magic
tech sky130A
magscale 1 2
timestamp 1643900835
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 252554 700380 252560 700392
rect 235224 700352 252560 700380
rect 235224 700340 235230 700352
rect 252554 700340 252560 700352
rect 252612 700340 252618 700392
rect 269758 700340 269764 700392
rect 269816 700380 269822 700392
rect 283834 700380 283840 700392
rect 269816 700352 283840 700380
rect 269816 700340 269822 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 395338 700340 395344 700392
rect 395396 700380 395402 700392
rect 494790 700380 494796 700392
rect 395396 700352 494796 700380
rect 395396 700340 395402 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 215938 700312 215944 700324
rect 24360 700284 215944 700312
rect 24360 700272 24366 700284
rect 215938 700272 215944 700284
rect 215996 700272 216002 700324
rect 238018 700272 238024 700324
rect 238076 700312 238082 700324
rect 413646 700312 413652 700324
rect 238076 700284 413652 700312
rect 238076 700272 238082 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 453298 700272 453304 700324
rect 453356 700312 453362 700324
rect 462314 700312 462320 700324
rect 453356 700284 462320 700312
rect 453356 700272 453362 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 497458 700272 497464 700324
rect 497516 700312 497522 700324
rect 559650 700312 559656 700324
rect 497516 700284 559656 700312
rect 497516 700272 497522 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 155218 700108 155224 700120
rect 154172 700080 155224 700108
rect 154172 700068 154178 700080
rect 155218 700068 155224 700080
rect 155276 700068 155282 700120
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 363598 699660 363604 699712
rect 363656 699700 363662 699712
rect 364978 699700 364984 699712
rect 363656 699672 364984 699700
rect 363656 699660 363662 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 475378 699660 475384 699712
rect 475436 699700 475442 699712
rect 478506 699700 478512 699712
rect 475436 699672 478512 699700
rect 475436 699660 475442 699672
rect 478506 699660 478512 699672
rect 478564 699660 478570 699712
rect 249058 698912 249064 698964
rect 249116 698952 249122 698964
rect 527174 698952 527180 698964
rect 249116 698924 527180 698952
rect 249116 698912 249122 698924
rect 527174 698912 527180 698924
rect 527232 698912 527238 698964
rect 266354 697620 266360 697672
rect 266412 697660 266418 697672
rect 267642 697660 267648 697672
rect 266412 697632 267648 697660
rect 266412 697620 266418 697632
rect 267642 697620 267648 697632
rect 267700 697620 267706 697672
rect 180702 697552 180708 697604
rect 180760 697592 180766 697604
rect 397454 697592 397460 697604
rect 180760 697564 397460 697592
rect 180760 697552 180766 697564
rect 397454 697552 397460 697564
rect 397512 697552 397518 697604
rect 222838 696192 222844 696244
rect 222896 696232 222902 696244
rect 348786 696232 348792 696244
rect 222896 696204 348792 696232
rect 222896 696192 222902 696204
rect 348786 696192 348792 696204
rect 348844 696192 348850 696244
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 196618 670732 196624 670744
rect 3568 670704 196624 670732
rect 3568 670692 3574 670704
rect 196618 670692 196624 670704
rect 196676 670692 196682 670744
rect 73062 665796 73068 665848
rect 73120 665836 73126 665848
rect 240502 665836 240508 665848
rect 73120 665808 240508 665836
rect 73120 665796 73126 665808
rect 240502 665796 240508 665808
rect 240560 665796 240566 665848
rect 202138 660288 202144 660340
rect 202196 660328 202202 660340
rect 331214 660328 331220 660340
rect 202196 660300 331220 660328
rect 202196 660288 202202 660300
rect 331214 660288 331220 660300
rect 331272 660288 331278 660340
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 112438 656928 112444 656940
rect 3568 656900 112444 656928
rect 3568 656888 3574 656900
rect 112438 656888 112444 656900
rect 112496 656888 112502 656940
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 166258 632108 166264 632120
rect 3568 632080 166264 632108
rect 3568 632068 3574 632080
rect 166258 632068 166264 632080
rect 166316 632068 166322 632120
rect 191742 623024 191748 623076
rect 191800 623064 191806 623076
rect 299474 623064 299480 623076
rect 191800 623036 299480 623064
rect 191800 623024 191806 623036
rect 299474 623024 299480 623036
rect 299532 623024 299538 623076
rect 2774 619080 2780 619132
rect 2832 619120 2838 619132
rect 4798 619120 4804 619132
rect 2832 619092 4804 619120
rect 2832 619080 2838 619092
rect 4798 619080 4804 619092
rect 4856 619080 4862 619132
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 220078 605860 220084 605872
rect 3568 605832 220084 605860
rect 3568 605820 3574 605832
rect 220078 605820 220084 605832
rect 220136 605820 220142 605872
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 226978 579680 226984 579692
rect 3384 579652 226984 579680
rect 3384 579640 3390 579652
rect 226978 579640 226984 579652
rect 227036 579640 227042 579692
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 68278 565876 68284 565888
rect 3292 565848 68284 565876
rect 3292 565836 3298 565848
rect 68278 565836 68284 565848
rect 68336 565836 68342 565888
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 35158 553432 35164 553444
rect 3384 553404 35164 553432
rect 3384 553392 3390 553404
rect 35158 553392 35164 553404
rect 35216 553392 35222 553444
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 71038 527184 71044 527196
rect 3016 527156 71044 527184
rect 3016 527144 3022 527156
rect 71038 527144 71044 527156
rect 71096 527144 71102 527196
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 162118 514808 162124 514820
rect 3568 514780 162124 514808
rect 3568 514768 3574 514780
rect 162118 514768 162124 514780
rect 162176 514768 162182 514820
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 233878 501004 233884 501016
rect 3108 500976 233884 501004
rect 3108 500964 3114 500976
rect 233878 500964 233884 500976
rect 233936 500964 233942 501016
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 244918 474756 244924 474768
rect 3108 474728 244924 474756
rect 3108 474716 3114 474728
rect 244918 474716 244924 474728
rect 244976 474716 244982 474768
rect 3418 462952 3424 463004
rect 3476 462992 3482 463004
rect 258074 462992 258080 463004
rect 3476 462964 258080 462992
rect 3476 462952 3482 462964
rect 258074 462952 258080 462964
rect 258132 462952 258138 463004
rect 188982 456764 188988 456816
rect 189040 456804 189046 456816
rect 580166 456804 580172 456816
rect 189040 456776 580172 456804
rect 189040 456764 189046 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 204898 448576 204904 448588
rect 3200 448548 204904 448576
rect 3200 448536 3206 448548
rect 204898 448536 204904 448548
rect 204956 448536 204962 448588
rect 309778 430584 309784 430636
rect 309836 430624 309842 430636
rect 580166 430624 580172 430636
rect 309836 430596 580172 430624
rect 309836 430584 309842 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 21358 422328 21364 422340
rect 3476 422300 21364 422328
rect 3476 422288 3482 422300
rect 21358 422288 21364 422300
rect 21416 422288 21422 422340
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 29638 409884 29644 409896
rect 2924 409856 29644 409884
rect 2924 409844 2930 409856
rect 29638 409844 29644 409856
rect 29696 409844 29702 409896
rect 206278 404336 206284 404388
rect 206336 404376 206342 404388
rect 580166 404376 580172 404388
rect 206336 404348 580172 404376
rect 206336 404336 206342 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 177298 397508 177304 397520
rect 3476 397480 177304 397508
rect 3476 397468 3482 397480
rect 177298 397468 177304 397480
rect 177356 397468 177362 397520
rect 21358 382916 21364 382968
rect 21416 382956 21422 382968
rect 209038 382956 209044 382968
rect 21416 382928 209044 382956
rect 21416 382916 21422 382928
rect 209038 382916 209044 382928
rect 209096 382916 209102 382968
rect 198642 380128 198648 380180
rect 198700 380168 198706 380180
rect 583570 380168 583576 380180
rect 198700 380140 583576 380168
rect 198700 380128 198706 380140
rect 583570 380128 583576 380140
rect 583628 380128 583634 380180
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 21358 371260 21364 371272
rect 3476 371232 21364 371260
rect 3476 371220 3482 371232
rect 21358 371220 21364 371232
rect 21416 371220 21422 371272
rect 305638 364352 305644 364404
rect 305696 364392 305702 364404
rect 579614 364392 579620 364404
rect 305696 364364 579620 364392
rect 305696 364352 305702 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 15838 357456 15844 357468
rect 3200 357428 15844 357456
rect 3200 357416 3206 357428
rect 15838 357416 15844 357428
rect 15896 357416 15902 357468
rect 246298 356668 246304 356720
rect 246356 356708 246362 356720
rect 583018 356708 583024 356720
rect 246356 356680 583024 356708
rect 246356 356668 246362 356680
rect 583018 356668 583024 356680
rect 583076 356668 583082 356720
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 232498 345080 232504 345092
rect 3384 345052 232504 345080
rect 3384 345040 3390 345052
rect 232498 345040 232504 345052
rect 232556 345040 232562 345092
rect 15838 338716 15844 338768
rect 15896 338756 15902 338768
rect 228358 338756 228364 338768
rect 15896 338728 228364 338756
rect 15896 338716 15902 338728
rect 228358 338716 228364 338728
rect 228416 338716 228422 338768
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 224218 318832 224224 318844
rect 3384 318804 224224 318832
rect 3384 318792 3390 318804
rect 224218 318792 224224 318804
rect 224276 318792 224282 318844
rect 566458 311856 566464 311908
rect 566516 311896 566522 311908
rect 579982 311896 579988 311908
rect 566516 311868 579988 311896
rect 566516 311856 566522 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3418 304988 3424 305040
rect 3476 305028 3482 305040
rect 249978 305028 249984 305040
rect 3476 305000 249984 305028
rect 3476 304988 3482 305000
rect 249978 304988 249984 305000
rect 250036 304988 250042 305040
rect 260190 302200 260196 302252
rect 260248 302240 260254 302252
rect 266354 302240 266360 302252
rect 260248 302212 266360 302240
rect 260248 302200 260254 302212
rect 266354 302200 266360 302212
rect 266412 302200 266418 302252
rect 226242 300092 226248 300144
rect 226300 300132 226306 300144
rect 583294 300132 583300 300144
rect 226300 300104 583300 300132
rect 226300 300092 226306 300104
rect 583294 300092 583300 300104
rect 583352 300092 583358 300144
rect 214558 298732 214564 298784
rect 214616 298772 214622 298784
rect 580258 298772 580264 298784
rect 214616 298744 580264 298772
rect 214616 298732 214622 298744
rect 580258 298732 580264 298744
rect 580316 298732 580322 298784
rect 209682 296692 209688 296744
rect 209740 296732 209746 296744
rect 264238 296732 264244 296744
rect 209740 296704 264244 296732
rect 209740 296692 209746 296704
rect 264238 296692 264244 296704
rect 264296 296692 264302 296744
rect 235718 295944 235724 295996
rect 235776 295984 235782 295996
rect 475378 295984 475384 295996
rect 235776 295956 475384 295984
rect 235776 295944 235782 295956
rect 475378 295944 475384 295956
rect 475436 295944 475442 295996
rect 202782 294652 202788 294704
rect 202840 294692 202846 294704
rect 244274 294692 244280 294704
rect 202840 294664 244280 294692
rect 202840 294652 202846 294664
rect 244274 294652 244280 294664
rect 244332 294652 244338 294704
rect 213822 294584 213828 294636
rect 213880 294624 213886 294636
rect 582374 294624 582380 294636
rect 213880 294596 582380 294624
rect 213880 294584 213886 294596
rect 582374 294584 582380 294596
rect 582432 294584 582438 294636
rect 227622 293972 227628 294024
rect 227680 294012 227686 294024
rect 273898 294012 273904 294024
rect 227680 293984 273904 294012
rect 227680 293972 227686 293984
rect 273898 293972 273904 293984
rect 273956 293972 273962 294024
rect 195790 293224 195796 293276
rect 195848 293264 195854 293276
rect 429194 293264 429200 293276
rect 195848 293236 429200 293264
rect 195848 293224 195854 293236
rect 429194 293224 429200 293236
rect 429252 293224 429258 293276
rect 219342 292680 219348 292732
rect 219400 292720 219406 292732
rect 251174 292720 251180 292732
rect 219400 292692 251180 292720
rect 219400 292680 219406 292692
rect 251174 292680 251180 292692
rect 251232 292680 251238 292732
rect 232590 292612 232596 292664
rect 232648 292652 232654 292664
rect 304994 292652 305000 292664
rect 232648 292624 305000 292652
rect 232648 292612 232654 292624
rect 304994 292612 305000 292624
rect 305052 292612 305058 292664
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 11698 292584 11704 292596
rect 3476 292556 11704 292584
rect 3476 292544 3482 292556
rect 11698 292544 11704 292556
rect 11756 292544 11762 292596
rect 236914 292544 236920 292596
rect 236972 292584 236978 292596
rect 583662 292584 583668 292596
rect 236972 292556 583668 292584
rect 236972 292544 236978 292556
rect 583662 292544 583668 292556
rect 583720 292544 583726 292596
rect 224218 291932 224224 291984
rect 224276 291972 224282 291984
rect 240134 291972 240140 291984
rect 224276 291944 240140 291972
rect 224276 291932 224282 291944
rect 240134 291932 240140 291944
rect 240192 291932 240198 291984
rect 112438 291864 112444 291916
rect 112496 291904 112502 291916
rect 245654 291904 245660 291916
rect 112496 291876 245660 291904
rect 112496 291864 112502 291876
rect 245654 291864 245660 291876
rect 245712 291864 245718 291916
rect 211062 291796 211068 291848
rect 211120 291836 211126 291848
rect 583018 291836 583024 291848
rect 211120 291808 583024 291836
rect 211120 291796 211126 291808
rect 583018 291796 583024 291808
rect 583076 291796 583082 291848
rect 224862 291252 224868 291304
rect 224920 291292 224926 291304
rect 247034 291292 247040 291304
rect 224920 291264 247040 291292
rect 224920 291252 224926 291264
rect 247034 291252 247040 291264
rect 247092 291252 247098 291304
rect 242710 291184 242716 291236
rect 242768 291224 242774 291236
rect 271138 291224 271144 291236
rect 242768 291196 271144 291224
rect 242768 291184 242774 291196
rect 271138 291184 271144 291196
rect 271196 291184 271202 291236
rect 89622 290504 89628 290556
rect 89680 290544 89686 290556
rect 232774 290544 232780 290556
rect 89680 290516 232780 290544
rect 89680 290504 89686 290516
rect 232774 290504 232780 290516
rect 232832 290504 232838 290556
rect 232498 290436 232504 290488
rect 232556 290476 232562 290488
rect 243814 290476 243820 290488
rect 232556 290448 243820 290476
rect 232556 290436 232562 290448
rect 243814 290436 243820 290448
rect 243872 290436 243878 290488
rect 14 290096 20 290148
rect 72 290136 78 290148
rect 242894 290136 242900 290148
rect 72 290108 242900 290136
rect 72 290096 78 290108
rect 242894 290096 242900 290108
rect 242952 290096 242958 290148
rect 216490 290028 216496 290080
rect 216548 290068 216554 290080
rect 253934 290068 253940 290080
rect 216548 290040 253940 290068
rect 216548 290028 216554 290040
rect 253934 290028 253940 290040
rect 253992 290028 253998 290080
rect 215202 289960 215208 290012
rect 215260 290000 215266 290012
rect 260834 290000 260840 290012
rect 215260 289972 260840 290000
rect 215260 289960 215266 289972
rect 260834 289960 260840 289972
rect 260892 289960 260898 290012
rect 235810 289892 235816 289944
rect 235868 289932 235874 289944
rect 260098 289932 260104 289944
rect 235868 289904 260104 289932
rect 235868 289892 235874 289904
rect 260098 289892 260104 289904
rect 260156 289892 260162 289944
rect 239950 289824 239956 289876
rect 240008 289864 240014 289876
rect 574738 289864 574744 289876
rect 240008 289836 574744 289864
rect 240008 289824 240014 289836
rect 574738 289824 574744 289836
rect 574796 289824 574802 289876
rect 215938 289756 215944 289808
rect 215996 289796 216002 289808
rect 218238 289796 218244 289808
rect 215996 289768 218244 289796
rect 215996 289756 216002 289768
rect 218238 289756 218244 289768
rect 218296 289756 218302 289808
rect 200390 289144 200396 289196
rect 200448 289184 200454 289196
rect 206278 289184 206284 289196
rect 200448 289156 206284 289184
rect 200448 289144 200454 289156
rect 206278 289144 206284 289156
rect 206336 289144 206342 289196
rect 155218 289076 155224 289128
rect 155276 289116 155282 289128
rect 204254 289116 204260 289128
rect 155276 289088 204260 289116
rect 155276 289076 155282 289088
rect 204254 289076 204260 289088
rect 204312 289076 204318 289128
rect 233878 289076 233884 289128
rect 233936 289116 233942 289128
rect 245838 289116 245844 289128
rect 233936 289088 245844 289116
rect 233936 289076 233942 289088
rect 245838 289076 245844 289088
rect 245896 289076 245902 289128
rect 236638 288600 236644 288652
rect 236696 288640 236702 288652
rect 249794 288640 249800 288652
rect 236696 288612 249800 288640
rect 236696 288600 236702 288612
rect 249794 288600 249800 288612
rect 249852 288600 249858 288652
rect 240870 288532 240876 288584
rect 240928 288572 240934 288584
rect 255958 288572 255964 288584
rect 240928 288544 255964 288572
rect 240928 288532 240934 288544
rect 255958 288532 255964 288544
rect 256016 288532 256022 288584
rect 237374 288464 237380 288516
rect 237432 288504 237438 288516
rect 265618 288504 265624 288516
rect 237432 288476 265624 288504
rect 237432 288464 237438 288476
rect 265618 288464 265624 288476
rect 265676 288464 265682 288516
rect 206646 288396 206652 288448
rect 206704 288436 206710 288448
rect 583018 288436 583024 288448
rect 206704 288408 583024 288436
rect 206704 288396 206710 288408
rect 583018 288396 583024 288408
rect 583076 288396 583082 288448
rect 220078 288328 220084 288380
rect 220136 288368 220142 288380
rect 225414 288368 225420 288380
rect 220136 288340 225420 288368
rect 220136 288328 220142 288340
rect 225414 288328 225420 288340
rect 225472 288328 225478 288380
rect 235902 288328 235908 288380
rect 235960 288368 235966 288380
rect 238018 288368 238024 288380
rect 235960 288340 238024 288368
rect 235960 288328 235966 288340
rect 238018 288328 238024 288340
rect 238076 288328 238082 288380
rect 229830 287376 229836 287428
rect 229888 287416 229894 287428
rect 255314 287416 255320 287428
rect 229888 287388 255320 287416
rect 229888 287376 229894 287388
rect 255314 287376 255320 287388
rect 255372 287376 255378 287428
rect 239582 287308 239588 287360
rect 239640 287348 239646 287360
rect 266998 287348 267004 287360
rect 239640 287320 267004 287348
rect 239640 287308 239646 287320
rect 266998 287308 267004 287320
rect 267056 287308 267062 287360
rect 57238 287240 57244 287292
rect 57296 287280 57302 287292
rect 230382 287280 230388 287292
rect 57296 287252 230388 287280
rect 57296 287240 57302 287252
rect 230382 287240 230388 287252
rect 230440 287240 230446 287292
rect 233142 287240 233148 287292
rect 233200 287280 233206 287292
rect 302878 287280 302884 287292
rect 233200 287252 302884 287280
rect 233200 287240 233206 287252
rect 302878 287240 302884 287252
rect 302936 287240 302942 287292
rect 201310 287172 201316 287224
rect 201368 287212 201374 287224
rect 309134 287212 309140 287224
rect 201368 287184 309140 287212
rect 201368 287172 201374 287184
rect 309134 287172 309140 287184
rect 309192 287172 309198 287224
rect 201678 287104 201684 287156
rect 201736 287144 201742 287156
rect 334618 287144 334624 287156
rect 201736 287116 334624 287144
rect 201736 287104 201742 287116
rect 334618 287104 334624 287116
rect 334676 287104 334682 287156
rect 196618 287036 196624 287088
rect 196676 287076 196682 287088
rect 202782 287076 202788 287088
rect 196676 287048 202788 287076
rect 196676 287036 196682 287048
rect 202782 287036 202788 287048
rect 202840 287036 202846 287088
rect 222102 287036 222108 287088
rect 222160 287076 222166 287088
rect 302234 287076 302240 287088
rect 222160 287048 302240 287076
rect 222160 287036 222166 287048
rect 302234 287036 302240 287048
rect 302292 287036 302298 287088
rect 218606 286424 218612 286476
rect 218664 286464 218670 286476
rect 222838 286464 222844 286476
rect 218664 286436 222844 286464
rect 218664 286424 218670 286436
rect 222838 286424 222844 286436
rect 222896 286424 222902 286476
rect 208486 286356 208492 286408
rect 208544 286396 208550 286408
rect 232590 286396 232596 286408
rect 208544 286368 232596 286396
rect 208544 286356 208550 286368
rect 232590 286356 232596 286368
rect 232648 286356 232654 286408
rect 210878 286288 210884 286340
rect 210936 286328 210942 286340
rect 236638 286328 236644 286340
rect 210936 286300 236644 286328
rect 210936 286288 210942 286300
rect 236638 286288 236644 286300
rect 236696 286288 236702 286340
rect 195882 286016 195888 286068
rect 195940 286056 195946 286068
rect 203150 286056 203156 286068
rect 195940 286028 203156 286056
rect 195940 286016 195946 286028
rect 203150 286016 203156 286028
rect 203208 286016 203214 286068
rect 231670 286016 231676 286068
rect 231728 286056 231734 286068
rect 243998 286056 244004 286068
rect 231728 286028 244004 286056
rect 231728 286016 231734 286028
rect 243998 286016 244004 286028
rect 244056 286016 244062 286068
rect 182082 285948 182088 286000
rect 182140 285988 182146 286000
rect 204622 285988 204628 286000
rect 182140 285960 204628 285988
rect 182140 285948 182146 285960
rect 204622 285948 204628 285960
rect 204680 285948 204686 286000
rect 236086 285948 236092 286000
rect 236144 285988 236150 286000
rect 253198 285988 253204 286000
rect 236144 285960 253204 285988
rect 236144 285948 236150 285960
rect 253198 285948 253204 285960
rect 253256 285948 253262 286000
rect 43438 285880 43444 285932
rect 43496 285920 43502 285932
rect 206094 285920 206100 285932
rect 43496 285892 206100 285920
rect 43496 285880 43502 285892
rect 206094 285880 206100 285892
rect 206152 285880 206158 285932
rect 232222 285880 232228 285932
rect 232280 285920 232286 285932
rect 262858 285920 262864 285932
rect 232280 285892 262864 285920
rect 232280 285880 232286 285892
rect 262858 285880 262864 285892
rect 262916 285880 262922 285932
rect 194502 285812 194508 285864
rect 194560 285852 194566 285864
rect 203702 285852 203708 285864
rect 194560 285824 203708 285852
rect 194560 285812 194566 285824
rect 203702 285812 203708 285824
rect 203760 285812 203766 285864
rect 207014 285852 207020 285864
rect 204732 285824 207020 285852
rect 200022 285744 200028 285796
rect 200080 285784 200086 285796
rect 204732 285784 204760 285824
rect 207014 285812 207020 285824
rect 207072 285812 207078 285864
rect 227806 285812 227812 285864
rect 227864 285852 227870 285864
rect 276658 285852 276664 285864
rect 227864 285824 276664 285852
rect 227864 285812 227870 285824
rect 276658 285812 276664 285824
rect 276716 285812 276722 285864
rect 205542 285784 205548 285796
rect 200080 285756 204760 285784
rect 204824 285756 205548 285784
rect 200080 285744 200086 285756
rect 199930 285676 199936 285728
rect 199988 285716 199994 285728
rect 204824 285716 204852 285756
rect 205542 285744 205548 285756
rect 205600 285744 205606 285796
rect 213454 285744 213460 285796
rect 213512 285784 213518 285796
rect 214558 285784 214564 285796
rect 213512 285756 214564 285784
rect 213512 285744 213518 285756
rect 214558 285744 214564 285756
rect 214616 285744 214622 285796
rect 214742 285744 214748 285796
rect 214800 285784 214806 285796
rect 221182 285784 221188 285796
rect 214800 285756 221188 285784
rect 214800 285744 214806 285756
rect 221182 285744 221188 285756
rect 221240 285744 221246 285796
rect 221550 285744 221556 285796
rect 221608 285784 221614 285796
rect 221608 285756 229094 285784
rect 221608 285744 221614 285756
rect 199988 285688 204852 285716
rect 199988 285676 199994 285688
rect 204898 285676 204904 285728
rect 204956 285716 204962 285728
rect 208118 285716 208124 285728
rect 204956 285688 208124 285716
rect 204956 285676 204962 285688
rect 208118 285676 208124 285688
rect 208176 285676 208182 285728
rect 209958 285676 209964 285728
rect 210016 285716 210022 285728
rect 211062 285716 211068 285728
rect 210016 285688 211068 285716
rect 210016 285676 210022 285688
rect 211062 285676 211068 285688
rect 211120 285676 211126 285728
rect 212902 285676 212908 285728
rect 212960 285716 212966 285728
rect 213822 285716 213828 285728
rect 212960 285688 213828 285716
rect 212960 285676 212966 285688
rect 213822 285676 213828 285688
rect 213880 285676 213886 285728
rect 214374 285676 214380 285728
rect 214432 285716 214438 285728
rect 215202 285716 215208 285728
rect 214432 285688 215208 285716
rect 214432 285676 214438 285688
rect 215202 285676 215208 285688
rect 215260 285676 215266 285728
rect 215294 285676 215300 285728
rect 215352 285716 215358 285728
rect 216582 285716 216588 285728
rect 215352 285688 216588 285716
rect 215352 285676 215358 285688
rect 216582 285676 216588 285688
rect 216640 285676 216646 285728
rect 223574 285676 223580 285728
rect 223632 285716 223638 285728
rect 224862 285716 224868 285728
rect 223632 285688 224868 285716
rect 223632 285676 223638 285688
rect 224862 285676 224868 285688
rect 224920 285676 224926 285728
rect 226518 285676 226524 285728
rect 226576 285716 226582 285728
rect 227622 285716 227628 285728
rect 226576 285688 227628 285716
rect 226576 285676 226582 285688
rect 227622 285676 227628 285688
rect 227680 285676 227686 285728
rect 229066 285716 229094 285756
rect 234614 285744 234620 285796
rect 234672 285784 234678 285796
rect 235718 285784 235724 285796
rect 234672 285756 235724 285784
rect 234672 285744 234678 285756
rect 235718 285744 235724 285756
rect 235776 285744 235782 285796
rect 239030 285744 239036 285796
rect 239088 285784 239094 285796
rect 239950 285784 239956 285796
rect 239088 285756 239956 285784
rect 239088 285744 239094 285756
rect 239950 285744 239956 285756
rect 240008 285744 240014 285796
rect 241974 285744 241980 285796
rect 242032 285784 242038 285796
rect 291194 285784 291200 285796
rect 242032 285756 291200 285784
rect 242032 285744 242038 285756
rect 291194 285744 291200 285756
rect 291252 285744 291258 285796
rect 303614 285716 303620 285728
rect 229066 285688 303620 285716
rect 303614 285676 303620 285688
rect 303672 285676 303678 285728
rect 240134 285268 240140 285320
rect 240192 285308 240198 285320
rect 241054 285308 241060 285320
rect 240192 285280 241060 285308
rect 240192 285268 240198 285280
rect 241054 285268 241060 285280
rect 241112 285268 241118 285320
rect 215846 284928 215852 284980
rect 215904 284968 215910 284980
rect 237374 284968 237380 284980
rect 215904 284940 237380 284968
rect 215904 284928 215910 284940
rect 237374 284928 237380 284940
rect 237432 284928 237438 284980
rect 221182 284656 221188 284708
rect 221240 284696 221246 284708
rect 264330 284696 264336 284708
rect 221240 284668 264336 284696
rect 221240 284656 221246 284668
rect 264330 284656 264336 284668
rect 264388 284656 264394 284708
rect 237006 284588 237012 284640
rect 237064 284628 237070 284640
rect 249886 284628 249892 284640
rect 237064 284600 249892 284628
rect 237064 284588 237070 284600
rect 249886 284588 249892 284600
rect 249944 284588 249950 284640
rect 212350 284520 212356 284572
rect 212408 284560 212414 284572
rect 249150 284560 249156 284572
rect 212408 284532 249156 284560
rect 212408 284520 212414 284532
rect 249150 284520 249156 284532
rect 249208 284520 249214 284572
rect 173158 284452 173164 284504
rect 173216 284492 173222 284504
rect 223942 284492 223948 284504
rect 173216 284464 223948 284492
rect 173216 284452 173222 284464
rect 223942 284452 223948 284464
rect 224000 284452 224006 284504
rect 238110 284452 238116 284504
rect 238168 284492 238174 284504
rect 261478 284492 261484 284504
rect 238168 284464 261484 284492
rect 238168 284452 238174 284464
rect 261478 284452 261484 284464
rect 261536 284452 261542 284504
rect 65518 284384 65524 284436
rect 65576 284424 65582 284436
rect 213822 284424 213828 284436
rect 65576 284396 213828 284424
rect 65576 284384 65582 284396
rect 213822 284384 213828 284396
rect 213880 284384 213886 284436
rect 237558 284384 237564 284436
rect 237616 284424 237622 284436
rect 244090 284424 244096 284436
rect 237616 284396 244096 284424
rect 237616 284384 237622 284396
rect 244090 284384 244096 284396
rect 244148 284384 244154 284436
rect 17218 284316 17224 284368
rect 17276 284356 17282 284368
rect 227438 284356 227444 284368
rect 17276 284328 227444 284356
rect 17276 284316 17282 284328
rect 227438 284316 227444 284328
rect 227496 284316 227502 284368
rect 239950 284316 239956 284368
rect 240008 284356 240014 284368
rect 299474 284356 299480 284368
rect 240008 284328 299480 284356
rect 240008 284316 240014 284328
rect 299474 284316 299480 284328
rect 299532 284316 299538 284368
rect 201494 284180 201500 284232
rect 201552 284220 201558 284232
rect 202138 284220 202144 284232
rect 201552 284192 202144 284220
rect 201552 284180 201558 284192
rect 202138 284180 202144 284192
rect 202196 284180 202202 284232
rect 234522 283908 234528 283960
rect 234580 283948 234586 283960
rect 234580 283920 238754 283948
rect 234580 283908 234586 283920
rect 238726 283880 238754 283920
rect 284294 283880 284300 283892
rect 238726 283852 284300 283880
rect 284294 283840 284300 283852
rect 284352 283840 284358 283892
rect 244090 283568 244096 283620
rect 244148 283608 244154 283620
rect 282914 283608 282920 283620
rect 244148 283580 282920 283608
rect 244148 283568 244154 283580
rect 282914 283568 282920 283580
rect 282972 283568 282978 283620
rect 246022 282820 246028 282872
rect 246080 282860 246086 282872
rect 583570 282860 583576 282872
rect 246080 282832 583576 282860
rect 246080 282820 246086 282832
rect 583570 282820 583576 282832
rect 583628 282820 583634 282872
rect 183462 281596 183468 281648
rect 183520 281636 183526 281648
rect 197446 281636 197452 281648
rect 183520 281608 197452 281636
rect 183520 281596 183526 281608
rect 197446 281596 197452 281608
rect 197504 281596 197510 281648
rect 51718 281528 51724 281580
rect 51776 281568 51782 281580
rect 197354 281568 197360 281580
rect 51776 281540 197360 281568
rect 51776 281528 51782 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 245930 281528 245936 281580
rect 245988 281568 245994 281580
rect 254026 281568 254032 281580
rect 245988 281540 254032 281568
rect 245988 281528 245994 281540
rect 254026 281528 254032 281540
rect 254084 281528 254090 281580
rect 246022 280236 246028 280288
rect 246080 280276 246086 280288
rect 268378 280276 268384 280288
rect 246080 280248 268384 280276
rect 246080 280236 246086 280248
rect 268378 280236 268384 280248
rect 268436 280236 268442 280288
rect 245930 280168 245936 280220
rect 245988 280208 245994 280220
rect 271230 280208 271236 280220
rect 245988 280180 271236 280208
rect 245988 280168 245994 280180
rect 271230 280168 271236 280180
rect 271288 280168 271294 280220
rect 188890 278740 188896 278792
rect 188948 278780 188954 278792
rect 197354 278780 197360 278792
rect 188948 278752 197360 278780
rect 188948 278740 188954 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 245930 278740 245936 278792
rect 245988 278780 245994 278792
rect 583570 278780 583576 278792
rect 245988 278752 583576 278780
rect 245988 278740 245994 278752
rect 583570 278740 583576 278752
rect 583628 278740 583634 278792
rect 245930 278128 245936 278180
rect 245988 278168 245994 278180
rect 249978 278168 249984 278180
rect 245988 278140 249984 278168
rect 245988 278128 245994 278140
rect 249978 278128 249984 278140
rect 250036 278128 250042 278180
rect 194410 277720 194416 277772
rect 194468 277760 194474 277772
rect 197354 277760 197360 277772
rect 194468 277732 197360 277760
rect 194468 277720 194474 277732
rect 197354 277720 197360 277732
rect 197412 277720 197418 277772
rect 245930 277380 245936 277432
rect 245988 277420 245994 277432
rect 583478 277420 583484 277432
rect 245988 277392 583484 277420
rect 245988 277380 245994 277392
rect 583478 277380 583484 277392
rect 583536 277380 583542 277432
rect 191650 276020 191656 276072
rect 191708 276060 191714 276072
rect 197446 276060 197452 276072
rect 191708 276032 197452 276060
rect 191708 276020 191714 276032
rect 197446 276020 197452 276032
rect 197504 276020 197510 276072
rect 246022 276020 246028 276072
rect 246080 276060 246086 276072
rect 280798 276060 280804 276072
rect 246080 276032 280804 276060
rect 246080 276020 246086 276032
rect 280798 276020 280804 276032
rect 280856 276020 280862 276072
rect 4798 275952 4804 276004
rect 4856 275992 4862 276004
rect 197354 275992 197360 276004
rect 4856 275964 197360 275992
rect 4856 275952 4862 275964
rect 197354 275952 197360 275964
rect 197412 275952 197418 276004
rect 245930 275952 245936 276004
rect 245988 275992 245994 276004
rect 583846 275992 583852 276004
rect 245988 275964 583852 275992
rect 245988 275952 245994 275964
rect 583846 275952 583852 275964
rect 583904 275952 583910 276004
rect 245930 275340 245936 275392
rect 245988 275380 245994 275392
rect 249058 275380 249064 275392
rect 245988 275352 249064 275380
rect 245988 275340 245994 275352
rect 249058 275340 249064 275352
rect 249116 275340 249122 275392
rect 187602 274660 187608 274712
rect 187660 274700 187666 274712
rect 197354 274700 197360 274712
rect 187660 274672 197360 274700
rect 187660 274660 187666 274672
rect 197354 274660 197360 274672
rect 197412 274660 197418 274712
rect 8202 273912 8208 273964
rect 8260 273952 8266 273964
rect 178034 273952 178040 273964
rect 8260 273924 178040 273952
rect 8260 273912 8266 273924
rect 178034 273912 178040 273924
rect 178092 273912 178098 273964
rect 190362 273300 190368 273352
rect 190420 273340 190426 273352
rect 197446 273340 197452 273352
rect 190420 273312 197452 273340
rect 190420 273300 190426 273312
rect 197446 273300 197452 273312
rect 197504 273300 197510 273352
rect 245930 273300 245936 273352
rect 245988 273340 245994 273352
rect 256694 273340 256700 273352
rect 245988 273312 256700 273340
rect 245988 273300 245994 273312
rect 256694 273300 256700 273312
rect 256752 273300 256758 273352
rect 184842 273232 184848 273284
rect 184900 273272 184906 273284
rect 197354 273272 197360 273284
rect 184900 273244 197360 273272
rect 184900 273232 184906 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 246022 273232 246028 273284
rect 246080 273272 246086 273284
rect 295334 273272 295340 273284
rect 246080 273244 295340 273272
rect 246080 273232 246086 273244
rect 295334 273232 295340 273244
rect 295392 273232 295398 273284
rect 171042 273164 171048 273216
rect 171100 273204 171106 273216
rect 197446 273204 197452 273216
rect 171100 273176 197452 273204
rect 171100 273164 171106 273176
rect 197446 273164 197452 273176
rect 197504 273164 197510 273216
rect 246022 271940 246028 271992
rect 246080 271980 246086 271992
rect 255406 271980 255412 271992
rect 246080 271952 255412 271980
rect 246080 271940 246086 271952
rect 255406 271940 255412 271952
rect 255464 271940 255470 271992
rect 245930 271872 245936 271924
rect 245988 271912 245994 271924
rect 267090 271912 267096 271924
rect 245988 271884 267096 271912
rect 245988 271872 245994 271884
rect 267090 271872 267096 271884
rect 267148 271872 267154 271924
rect 304258 271872 304264 271924
rect 304316 271912 304322 271924
rect 579798 271912 579804 271924
rect 304316 271884 579804 271912
rect 304316 271872 304322 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 300118 271124 300124 271176
rect 300176 271164 300182 271176
rect 580350 271164 580356 271176
rect 300176 271136 580356 271164
rect 300176 271124 300182 271136
rect 580350 271124 580356 271136
rect 580408 271124 580414 271176
rect 187510 270580 187516 270632
rect 187568 270620 187574 270632
rect 197354 270620 197360 270632
rect 187568 270592 197360 270620
rect 187568 270580 187574 270592
rect 197354 270580 197360 270592
rect 197412 270580 197418 270632
rect 246022 270580 246028 270632
rect 246080 270620 246086 270632
rect 258166 270620 258172 270632
rect 246080 270592 258172 270620
rect 246080 270580 246086 270592
rect 258166 270580 258172 270592
rect 258224 270580 258230 270632
rect 186222 270512 186228 270564
rect 186280 270552 186286 270564
rect 197446 270552 197452 270564
rect 186280 270524 197452 270552
rect 186280 270512 186286 270524
rect 197446 270512 197452 270524
rect 197504 270512 197510 270564
rect 245930 270512 245936 270564
rect 245988 270552 245994 270564
rect 276750 270552 276756 270564
rect 245988 270524 276756 270552
rect 245988 270512 245994 270524
rect 276750 270512 276756 270524
rect 276808 270512 276814 270564
rect 193122 269152 193128 269204
rect 193180 269192 193186 269204
rect 197446 269192 197452 269204
rect 193180 269164 197452 269192
rect 193180 269152 193186 269164
rect 197446 269152 197452 269164
rect 197504 269152 197510 269204
rect 54478 269084 54484 269136
rect 54536 269124 54542 269136
rect 197354 269124 197360 269136
rect 54536 269096 197360 269124
rect 54536 269084 54542 269096
rect 197354 269084 197360 269096
rect 197412 269084 197418 269136
rect 245930 269084 245936 269136
rect 245988 269124 245994 269136
rect 285674 269124 285680 269136
rect 245988 269096 285680 269124
rect 245988 269084 245994 269096
rect 285674 269084 285680 269096
rect 285732 269084 285738 269136
rect 68278 269016 68284 269068
rect 68336 269056 68342 269068
rect 197446 269056 197452 269068
rect 68336 269028 197452 269056
rect 68336 269016 68342 269028
rect 197446 269016 197452 269028
rect 197504 269016 197510 269068
rect 178034 268948 178040 269000
rect 178092 268988 178098 269000
rect 197354 268988 197360 269000
rect 178092 268960 197360 268988
rect 178092 268948 178098 268960
rect 197354 268948 197360 268960
rect 197412 268948 197418 269000
rect 246022 267792 246028 267844
rect 246080 267832 246086 267844
rect 268470 267832 268476 267844
rect 246080 267804 268476 267832
rect 246080 267792 246086 267804
rect 268470 267792 268476 267804
rect 268528 267792 268534 267844
rect 245930 267724 245936 267776
rect 245988 267764 245994 267776
rect 583846 267764 583852 267776
rect 245988 267736 583852 267764
rect 245988 267724 245994 267736
rect 583846 267724 583852 267736
rect 583904 267724 583910 267776
rect 166258 267656 166264 267708
rect 166316 267696 166322 267708
rect 197354 267696 197360 267708
rect 166316 267668 197360 267696
rect 166316 267656 166322 267668
rect 197354 267656 197360 267668
rect 197412 267656 197418 267708
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 170398 266404 170404 266416
rect 3108 266376 170404 266404
rect 3108 266364 3114 266376
rect 170398 266364 170404 266376
rect 170456 266364 170462 266416
rect 195606 266364 195612 266416
rect 195664 266404 195670 266416
rect 197906 266404 197912 266416
rect 195664 266376 197912 266404
rect 195664 266364 195670 266376
rect 197906 266364 197912 266376
rect 197964 266364 197970 266416
rect 246022 266364 246028 266416
rect 246080 266404 246086 266416
rect 269850 266404 269856 266416
rect 246080 266376 269856 266404
rect 246080 266364 246086 266376
rect 269850 266364 269856 266376
rect 269908 266364 269914 266416
rect 245930 266296 245936 266348
rect 245988 266336 245994 266348
rect 566458 266336 566464 266348
rect 245988 266308 566464 266336
rect 245988 266296 245994 266308
rect 566458 266296 566464 266308
rect 566516 266296 566522 266348
rect 15838 264936 15844 264988
rect 15896 264976 15902 264988
rect 197446 264976 197452 264988
rect 15896 264948 197452 264976
rect 15896 264936 15902 264948
rect 197446 264936 197452 264948
rect 197504 264936 197510 264988
rect 245838 264936 245844 264988
rect 245896 264976 245902 264988
rect 251266 264976 251272 264988
rect 245896 264948 251272 264976
rect 245896 264936 245902 264948
rect 251266 264936 251272 264948
rect 251324 264936 251330 264988
rect 35158 264868 35164 264920
rect 35216 264908 35222 264920
rect 197354 264908 197360 264920
rect 35216 264880 197360 264908
rect 35216 264868 35222 264880
rect 197354 264868 197360 264880
rect 197412 264868 197418 264920
rect 184750 263576 184756 263628
rect 184808 263616 184814 263628
rect 197354 263616 197360 263628
rect 184808 263588 197360 263616
rect 184808 263576 184814 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 245930 263576 245936 263628
rect 245988 263616 245994 263628
rect 248414 263616 248420 263628
rect 245988 263588 248420 263616
rect 245988 263576 245994 263588
rect 248414 263576 248420 263588
rect 248472 263576 248478 263628
rect 193030 262216 193036 262268
rect 193088 262256 193094 262268
rect 197446 262256 197452 262268
rect 193088 262228 197452 262256
rect 193088 262216 193094 262228
rect 197446 262216 197452 262228
rect 197504 262216 197510 262268
rect 245930 262216 245936 262268
rect 245988 262256 245994 262268
rect 259454 262256 259460 262268
rect 245988 262228 259460 262256
rect 245988 262216 245994 262228
rect 259454 262216 259460 262228
rect 259512 262216 259518 262268
rect 71038 262148 71044 262200
rect 71096 262188 71102 262200
rect 197354 262188 197360 262200
rect 71096 262160 197360 262188
rect 71096 262148 71102 262160
rect 197354 262148 197360 262160
rect 197412 262148 197418 262200
rect 245838 260856 245844 260908
rect 245896 260896 245902 260908
rect 258258 260896 258264 260908
rect 245896 260868 258264 260896
rect 245896 260856 245902 260868
rect 258258 260856 258264 260868
rect 258316 260856 258322 260908
rect 244918 260720 244924 260772
rect 244976 260760 244982 260772
rect 245838 260760 245844 260772
rect 244976 260732 245844 260760
rect 244976 260720 244982 260732
rect 245838 260720 245844 260732
rect 245896 260720 245902 260772
rect 187418 259428 187424 259480
rect 187476 259468 187482 259480
rect 197354 259468 197360 259480
rect 187476 259440 197360 259468
rect 187476 259428 187482 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 245930 259428 245936 259480
rect 245988 259468 245994 259480
rect 300854 259468 300860 259480
rect 245988 259440 300860 259468
rect 245988 259428 245994 259440
rect 300854 259428 300860 259440
rect 300912 259428 300918 259480
rect 249150 259360 249156 259412
rect 249208 259400 249214 259412
rect 580166 259400 580172 259412
rect 249208 259372 580172 259400
rect 249208 259360 249214 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 191558 258544 191564 258596
rect 191616 258584 191622 258596
rect 197446 258584 197452 258596
rect 191616 258556 197452 258584
rect 191616 258544 191622 258556
rect 197446 258544 197452 258556
rect 197504 258544 197510 258596
rect 246022 258136 246028 258188
rect 246080 258176 246086 258188
rect 287054 258176 287060 258188
rect 246080 258148 287060 258176
rect 246080 258136 246086 258148
rect 287054 258136 287060 258148
rect 287112 258136 287118 258188
rect 32398 258068 32404 258120
rect 32456 258108 32462 258120
rect 197354 258108 197360 258120
rect 32456 258080 197360 258108
rect 32456 258068 32462 258080
rect 197354 258068 197360 258080
rect 197412 258068 197418 258120
rect 245930 258068 245936 258120
rect 245988 258108 245994 258120
rect 294046 258108 294052 258120
rect 245988 258080 294052 258108
rect 245988 258068 245994 258080
rect 294046 258068 294052 258080
rect 294104 258068 294110 258120
rect 3510 257320 3516 257372
rect 3568 257360 3574 257372
rect 178678 257360 178684 257372
rect 3568 257332 178684 257360
rect 3568 257320 3574 257332
rect 178678 257320 178684 257332
rect 178736 257320 178742 257372
rect 246390 257320 246396 257372
rect 246448 257360 246454 257372
rect 583294 257360 583300 257372
rect 246448 257332 583300 257360
rect 246448 257320 246454 257332
rect 583294 257320 583300 257332
rect 583352 257320 583358 257372
rect 195698 256776 195704 256828
rect 195756 256816 195762 256828
rect 197538 256816 197544 256828
rect 195756 256788 197544 256816
rect 195756 256776 195762 256788
rect 197538 256776 197544 256788
rect 197596 256776 197602 256828
rect 188798 256708 188804 256760
rect 188856 256748 188862 256760
rect 197354 256748 197360 256760
rect 188856 256720 197360 256748
rect 188856 256708 188862 256720
rect 197354 256708 197360 256720
rect 197412 256708 197418 256760
rect 245930 256708 245936 256760
rect 245988 256748 245994 256760
rect 272518 256748 272524 256760
rect 245988 256720 272524 256748
rect 245988 256708 245994 256720
rect 272518 256708 272524 256720
rect 272576 256708 272582 256760
rect 195790 256640 195796 256692
rect 195848 256680 195854 256692
rect 197906 256680 197912 256692
rect 195848 256652 197912 256680
rect 195848 256640 195854 256652
rect 197906 256640 197912 256652
rect 197964 256640 197970 256692
rect 245746 256640 245752 256692
rect 245804 256680 245810 256692
rect 583386 256680 583392 256692
rect 245804 256652 583392 256680
rect 245804 256640 245810 256652
rect 583386 256640 583392 256652
rect 583444 256640 583450 256692
rect 192938 255280 192944 255332
rect 192996 255320 193002 255332
rect 197354 255320 197360 255332
rect 192996 255292 197360 255320
rect 192996 255280 193002 255292
rect 197354 255280 197360 255292
rect 197412 255280 197418 255332
rect 137922 254532 137928 254584
rect 137980 254572 137986 254584
rect 147674 254572 147680 254584
rect 137980 254544 147680 254572
rect 137980 254532 137986 254544
rect 147674 254532 147680 254544
rect 147732 254532 147738 254584
rect 246482 254532 246488 254584
rect 246540 254572 246546 254584
rect 582742 254572 582748 254584
rect 246540 254544 582748 254572
rect 246540 254532 246546 254544
rect 582742 254532 582748 254544
rect 582800 254532 582806 254584
rect 191466 253988 191472 254040
rect 191524 254028 191530 254040
rect 197446 254028 197452 254040
rect 191524 254000 197452 254028
rect 191524 253988 191530 254000
rect 197446 253988 197452 254000
rect 197504 253988 197510 254040
rect 18598 253920 18604 253972
rect 18656 253960 18662 253972
rect 197354 253960 197360 253972
rect 18656 253932 197360 253960
rect 18656 253920 18662 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 245930 253920 245936 253972
rect 245988 253960 245994 253972
rect 252646 253960 252652 253972
rect 245988 253932 252652 253960
rect 245988 253920 245994 253932
rect 252646 253920 252652 253932
rect 252704 253920 252710 253972
rect 186130 253172 186136 253224
rect 186188 253212 186194 253224
rect 197998 253212 198004 253224
rect 186188 253184 198004 253212
rect 186188 253172 186194 253184
rect 197998 253172 198004 253184
rect 198056 253172 198062 253224
rect 194318 252968 194324 253020
rect 194376 253008 194382 253020
rect 198090 253008 198096 253020
rect 194376 252980 198096 253008
rect 194376 252968 194382 252980
rect 198090 252968 198096 252980
rect 198148 252968 198154 253020
rect 245930 252628 245936 252680
rect 245988 252668 245994 252680
rect 306374 252668 306380 252680
rect 245988 252640 306380 252668
rect 245988 252628 245994 252640
rect 306374 252628 306380 252640
rect 306432 252628 306438 252680
rect 180610 252560 180616 252612
rect 180668 252600 180674 252612
rect 197354 252600 197360 252612
rect 180668 252572 197360 252600
rect 180668 252560 180674 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 245838 252560 245844 252612
rect 245896 252600 245902 252612
rect 306466 252600 306472 252612
rect 245896 252572 306472 252600
rect 245896 252560 245902 252572
rect 306466 252560 306472 252572
rect 306524 252560 306530 252612
rect 245930 252492 245936 252544
rect 245988 252532 245994 252544
rect 258074 252532 258080 252544
rect 245988 252504 258080 252532
rect 245988 252492 245994 252504
rect 258074 252492 258080 252504
rect 258132 252492 258138 252544
rect 245930 251200 245936 251252
rect 245988 251240 245994 251252
rect 583386 251240 583392 251252
rect 245988 251212 583392 251240
rect 245988 251200 245994 251212
rect 583386 251200 583392 251212
rect 583444 251200 583450 251252
rect 147674 251132 147680 251184
rect 147732 251172 147738 251184
rect 197354 251172 197360 251184
rect 147732 251144 197360 251172
rect 147732 251132 147738 251144
rect 197354 251132 197360 251144
rect 197412 251132 197418 251184
rect 255958 250452 255964 250504
rect 256016 250492 256022 250504
rect 582742 250492 582748 250504
rect 256016 250464 582748 250492
rect 256016 250452 256022 250464
rect 582742 250452 582748 250464
rect 582800 250452 582806 250504
rect 245838 249772 245844 249824
rect 245896 249812 245902 249824
rect 307754 249812 307760 249824
rect 245896 249784 307760 249812
rect 245896 249772 245902 249784
rect 307754 249772 307760 249784
rect 307812 249772 307818 249824
rect 245930 249704 245936 249756
rect 245988 249744 245994 249756
rect 252554 249744 252560 249756
rect 245988 249716 252560 249744
rect 245988 249704 245994 249716
rect 252554 249704 252560 249716
rect 252612 249704 252618 249756
rect 190270 248480 190276 248532
rect 190328 248520 190334 248532
rect 197354 248520 197360 248532
rect 190328 248492 197360 248520
rect 190328 248480 190334 248492
rect 197354 248480 197360 248492
rect 197412 248480 197418 248532
rect 188706 248412 188712 248464
rect 188764 248452 188770 248464
rect 197446 248452 197452 248464
rect 188764 248424 197452 248452
rect 188764 248412 188770 248424
rect 197446 248412 197452 248424
rect 197504 248412 197510 248464
rect 180702 248344 180708 248396
rect 180760 248384 180766 248396
rect 197354 248384 197360 248396
rect 180760 248356 197360 248384
rect 180760 248344 180766 248356
rect 197354 248344 197360 248356
rect 197412 248344 197418 248396
rect 245838 248344 245844 248396
rect 245896 248384 245902 248396
rect 583754 248384 583760 248396
rect 245896 248356 583760 248384
rect 245896 248344 245902 248356
rect 583754 248344 583760 248356
rect 583812 248344 583818 248396
rect 245930 248276 245936 248328
rect 245988 248316 245994 248328
rect 309778 248316 309784 248328
rect 245988 248288 309784 248316
rect 245988 248276 245994 248288
rect 309778 248276 309784 248288
rect 309836 248276 309842 248328
rect 195790 247052 195796 247104
rect 195848 247092 195854 247104
rect 197630 247092 197636 247104
rect 195848 247064 197636 247092
rect 195848 247052 195854 247064
rect 197630 247052 197636 247064
rect 197688 247052 197694 247104
rect 29638 246984 29644 247036
rect 29696 247024 29702 247036
rect 197354 247024 197360 247036
rect 29696 246996 197360 247024
rect 29696 246984 29702 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 245930 245624 245936 245676
rect 245988 245664 245994 245676
rect 305178 245664 305184 245676
rect 245988 245636 305184 245664
rect 245988 245624 245994 245636
rect 305178 245624 305184 245636
rect 305236 245624 305242 245676
rect 245930 244264 245936 244316
rect 245988 244304 245994 244316
rect 251358 244304 251364 244316
rect 245988 244276 251364 244304
rect 245988 244264 245994 244276
rect 251358 244264 251364 244276
rect 251416 244264 251422 244316
rect 11698 244196 11704 244248
rect 11756 244236 11762 244248
rect 197354 244236 197360 244248
rect 11756 244208 197360 244236
rect 11756 244196 11762 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 191742 244128 191748 244180
rect 191800 244168 191806 244180
rect 197446 244168 197452 244180
rect 191800 244140 197452 244168
rect 191800 244128 191806 244140
rect 197446 244128 197452 244140
rect 197504 244128 197510 244180
rect 583846 243584 583852 243636
rect 583904 243584 583910 243636
rect 582742 243516 582748 243568
rect 582800 243556 582806 243568
rect 583754 243556 583760 243568
rect 582800 243528 583760 243556
rect 582800 243516 582806 243528
rect 583754 243516 583760 243528
rect 583812 243516 583818 243568
rect 583864 243432 583892 243584
rect 583846 243380 583852 243432
rect 583904 243380 583910 243432
rect 245838 242904 245844 242956
rect 245896 242944 245902 242956
rect 273990 242944 273996 242956
rect 245896 242916 273996 242944
rect 245896 242904 245902 242916
rect 273990 242904 273996 242916
rect 274048 242904 274054 242956
rect 188982 242836 188988 242888
rect 189040 242876 189046 242888
rect 197354 242876 197360 242888
rect 189040 242848 197360 242876
rect 189040 242836 189046 242848
rect 197354 242836 197360 242848
rect 197412 242836 197418 242888
rect 3418 242156 3424 242208
rect 3476 242196 3482 242208
rect 180058 242196 180064 242208
rect 3476 242168 180064 242196
rect 3476 242156 3482 242168
rect 180058 242156 180064 242168
rect 180116 242156 180122 242208
rect 245838 241544 245844 241596
rect 245896 241584 245902 241596
rect 269942 241584 269948 241596
rect 245896 241556 269948 241584
rect 245896 241544 245902 241556
rect 269942 241544 269948 241556
rect 270000 241544 270006 241596
rect 191742 241476 191748 241528
rect 191800 241516 191806 241528
rect 197446 241516 197452 241528
rect 191800 241488 197452 241516
rect 191800 241476 191806 241488
rect 197446 241476 197452 241488
rect 197504 241476 197510 241528
rect 244090 241476 244096 241528
rect 244148 241516 244154 241528
rect 579614 241516 579620 241528
rect 244148 241488 579620 241516
rect 244148 241476 244154 241488
rect 579614 241476 579620 241488
rect 579672 241476 579678 241528
rect 240520 240468 244274 240496
rect 199102 240184 199108 240236
rect 199160 240224 199166 240236
rect 199160 240196 213224 240224
rect 199160 240184 199166 240196
rect 213196 240168 213224 240196
rect 240520 240168 240548 240468
rect 244246 240428 244274 240468
rect 246022 240428 246028 240440
rect 241486 240400 242020 240428
rect 244246 240400 246028 240428
rect 241486 240292 241514 240400
rect 240612 240264 241514 240292
rect 241992 240292 242020 240400
rect 246022 240388 246028 240400
rect 246080 240388 246086 240440
rect 245930 240320 245936 240372
rect 245988 240360 245994 240372
rect 255498 240360 255504 240372
rect 245988 240332 255504 240360
rect 245988 240320 245994 240332
rect 255498 240320 255504 240332
rect 255556 240320 255562 240372
rect 269758 240292 269764 240304
rect 241992 240264 269764 240292
rect 240612 240168 240640 240264
rect 269758 240252 269764 240264
rect 269816 240252 269822 240304
rect 453298 240224 453304 240236
rect 240980 240196 453304 240224
rect 240980 240168 241008 240196
rect 453298 240184 453304 240196
rect 453356 240184 453362 240236
rect 3418 240116 3424 240168
rect 3476 240156 3482 240168
rect 3476 240128 209774 240156
rect 3476 240116 3482 240128
rect 209746 240088 209774 240128
rect 213178 240116 213184 240168
rect 213236 240116 213242 240168
rect 240502 240116 240508 240168
rect 240560 240116 240566 240168
rect 240594 240116 240600 240168
rect 240652 240116 240658 240168
rect 240962 240116 240968 240168
rect 241020 240116 241026 240168
rect 582466 240156 582472 240168
rect 241072 240128 582472 240156
rect 225230 240088 225236 240100
rect 209746 240060 225236 240088
rect 225230 240048 225236 240060
rect 225288 240048 225294 240100
rect 235902 240048 235908 240100
rect 235960 240088 235966 240100
rect 241072 240088 241100 240128
rect 582466 240116 582472 240128
rect 582524 240116 582530 240168
rect 235960 240060 241100 240088
rect 235960 240048 235966 240060
rect 241146 240048 241152 240100
rect 241204 240088 241210 240100
rect 582558 240088 582564 240100
rect 241204 240060 582564 240088
rect 241204 240048 241210 240060
rect 582558 240048 582564 240060
rect 582616 240048 582622 240100
rect 170398 239980 170404 240032
rect 170456 240020 170462 240032
rect 212718 240020 212724 240032
rect 170456 239992 212724 240020
rect 170456 239980 170462 239992
rect 212718 239980 212724 239992
rect 212776 239980 212782 240032
rect 238846 239980 238852 240032
rect 238904 240020 238910 240032
rect 497458 240020 497464 240032
rect 238904 239992 241100 240020
rect 238904 239980 238910 239992
rect 234982 239912 234988 239964
rect 235040 239952 235046 239964
rect 240962 239952 240968 239964
rect 235040 239924 240968 239952
rect 235040 239912 235046 239924
rect 240962 239912 240968 239924
rect 241020 239912 241026 239964
rect 241072 239952 241100 239992
rect 244246 239992 497464 240020
rect 244246 239952 244274 239992
rect 497458 239980 497464 239992
rect 497516 239980 497522 240032
rect 395338 239952 395344 239964
rect 241072 239924 244274 239952
rect 248386 239924 395344 239952
rect 162118 239844 162124 239896
rect 162176 239884 162182 239896
rect 242710 239884 242716 239896
rect 162176 239856 242716 239884
rect 162176 239844 162182 239856
rect 242710 239844 242716 239856
rect 242768 239844 242774 239896
rect 232590 239776 232596 239828
rect 232648 239816 232654 239828
rect 248386 239816 248414 239924
rect 395338 239912 395344 239924
rect 395396 239912 395402 239964
rect 232648 239788 248414 239816
rect 232648 239776 232654 239788
rect 199838 239504 199844 239556
rect 199896 239544 199902 239556
rect 209130 239544 209136 239556
rect 199896 239516 209136 239544
rect 199896 239504 199902 239516
rect 209130 239504 209136 239516
rect 209188 239504 209194 239556
rect 207934 239436 207940 239488
rect 207992 239476 207998 239488
rect 288618 239476 288624 239488
rect 207992 239448 288624 239476
rect 207992 239436 207998 239448
rect 288618 239436 288624 239448
rect 288676 239436 288682 239488
rect 106182 239368 106188 239420
rect 106240 239408 106246 239420
rect 209774 239408 209780 239420
rect 106240 239380 209780 239408
rect 106240 239368 106246 239380
rect 209774 239368 209780 239380
rect 209832 239368 209838 239420
rect 209774 238688 209780 238740
rect 209832 238728 209838 238740
rect 214558 238728 214564 238740
rect 209832 238700 214564 238728
rect 209832 238688 209838 238700
rect 214558 238688 214564 238700
rect 214616 238688 214622 238740
rect 239214 238688 239220 238740
rect 239272 238728 239278 238740
rect 244090 238728 244096 238740
rect 239272 238700 244096 238728
rect 239272 238688 239278 238700
rect 244090 238688 244096 238700
rect 244148 238688 244154 238740
rect 180058 238620 180064 238672
rect 180116 238660 180122 238672
rect 231486 238660 231492 238672
rect 180116 238632 231492 238660
rect 180116 238620 180122 238632
rect 231486 238620 231492 238632
rect 231544 238620 231550 238672
rect 236454 238620 236460 238672
rect 236512 238660 236518 238672
rect 582926 238660 582932 238672
rect 236512 238632 582932 238660
rect 236512 238620 236518 238632
rect 582926 238620 582932 238632
rect 582984 238620 582990 238672
rect 177298 238552 177304 238604
rect 177356 238592 177362 238604
rect 209222 238592 209228 238604
rect 177356 238564 209228 238592
rect 177356 238552 177362 238564
rect 209222 238552 209228 238564
rect 209280 238552 209286 238604
rect 216030 238552 216036 238604
rect 216088 238592 216094 238604
rect 304258 238592 304264 238604
rect 216088 238564 304264 238592
rect 216088 238552 216094 238564
rect 304258 238552 304264 238564
rect 304316 238552 304322 238604
rect 216582 238484 216588 238536
rect 216640 238524 216646 238536
rect 300118 238524 300124 238536
rect 216640 238496 300124 238524
rect 216640 238484 216646 238496
rect 300118 238484 300124 238496
rect 300176 238484 300182 238536
rect 21358 238416 21364 238468
rect 21416 238456 21422 238468
rect 221918 238456 221924 238468
rect 21416 238428 221924 238456
rect 21416 238416 21422 238428
rect 221918 238416 221924 238428
rect 221976 238416 221982 238468
rect 227622 238416 227628 238468
rect 227680 238456 227686 238468
rect 260190 238456 260196 238468
rect 227680 238428 260196 238456
rect 227680 238416 227686 238428
rect 260190 238416 260196 238428
rect 260248 238416 260254 238468
rect 233510 238348 233516 238400
rect 233568 238388 233574 238400
rect 583110 238388 583116 238400
rect 233568 238360 583116 238388
rect 233568 238348 233574 238360
rect 583110 238348 583116 238360
rect 583168 238348 583174 238400
rect 223758 238280 223764 238332
rect 223816 238320 223822 238332
rect 224770 238320 224776 238332
rect 223816 238292 224776 238320
rect 223816 238280 223822 238292
rect 224770 238280 224776 238292
rect 224828 238280 224834 238332
rect 234062 238280 234068 238332
rect 234120 238320 234126 238332
rect 234522 238320 234528 238332
rect 234120 238292 234528 238320
rect 234120 238280 234126 238292
rect 234522 238280 234528 238292
rect 234580 238280 234586 238332
rect 206462 238212 206468 238264
rect 206520 238252 206526 238264
rect 206922 238252 206928 238264
rect 206520 238224 206928 238252
rect 206520 238212 206526 238224
rect 206922 238212 206928 238224
rect 206980 238212 206986 238264
rect 211246 238076 211252 238128
rect 211304 238116 211310 238128
rect 220078 238116 220084 238128
rect 211304 238088 220084 238116
rect 211304 238076 211310 238088
rect 220078 238076 220084 238088
rect 220136 238076 220142 238128
rect 214190 238008 214196 238060
rect 214248 238048 214254 238060
rect 215018 238048 215024 238060
rect 214248 238020 215024 238048
rect 214248 238008 214254 238020
rect 215018 238008 215024 238020
rect 215076 238008 215082 238060
rect 220446 238008 220452 238060
rect 220504 238048 220510 238060
rect 238754 238048 238760 238060
rect 220504 238020 238760 238048
rect 220504 238008 220510 238020
rect 238754 238008 238760 238020
rect 238812 238008 238818 238060
rect 222838 237940 222844 237992
rect 222896 237980 222902 237992
rect 223482 237980 223488 237992
rect 222896 237952 223488 237980
rect 222896 237940 222902 237952
rect 223482 237940 223488 237952
rect 223540 237940 223546 237992
rect 230566 237804 230572 237856
rect 230624 237844 230630 237856
rect 231762 237844 231768 237856
rect 230624 237816 231768 237844
rect 230624 237804 230630 237816
rect 231762 237804 231768 237816
rect 231820 237804 231826 237856
rect 201494 237736 201500 237788
rect 201552 237776 201558 237788
rect 202690 237776 202696 237788
rect 201552 237748 202696 237776
rect 201552 237736 201558 237748
rect 202690 237736 202696 237748
rect 202748 237736 202754 237788
rect 200206 237668 200212 237720
rect 200264 237708 200270 237720
rect 201310 237708 201316 237720
rect 200264 237680 201316 237708
rect 200264 237668 200270 237680
rect 201310 237668 201316 237680
rect 201368 237668 201374 237720
rect 205910 237668 205916 237720
rect 205968 237708 205974 237720
rect 206738 237708 206744 237720
rect 205968 237680 206744 237708
rect 205968 237668 205974 237680
rect 206738 237668 206744 237680
rect 206796 237668 206802 237720
rect 207382 237668 207388 237720
rect 207440 237708 207446 237720
rect 208210 237708 208216 237720
rect 207440 237680 208216 237708
rect 207440 237668 207446 237680
rect 208210 237668 208216 237680
rect 208268 237668 208274 237720
rect 201126 237532 201132 237584
rect 201184 237572 201190 237584
rect 209038 237572 209044 237584
rect 201184 237544 209044 237572
rect 201184 237532 201190 237544
rect 209038 237532 209044 237544
rect 209096 237532 209102 237584
rect 202966 237464 202972 237516
rect 203024 237504 203030 237516
rect 203886 237504 203892 237516
rect 203024 237476 203892 237504
rect 203024 237464 203030 237476
rect 203886 237464 203892 237476
rect 203944 237464 203950 237516
rect 218054 237464 218060 237516
rect 218112 237504 218118 237516
rect 220170 237504 220176 237516
rect 218112 237476 220176 237504
rect 218112 237464 218118 237476
rect 220170 237464 220176 237476
rect 220228 237464 220234 237516
rect 200574 237396 200580 237448
rect 200632 237436 200638 237448
rect 201402 237436 201408 237448
rect 200632 237408 201408 237436
rect 200632 237396 200638 237408
rect 201402 237396 201408 237408
rect 201460 237396 201466 237448
rect 203518 237396 203524 237448
rect 203576 237436 203582 237448
rect 203978 237436 203984 237448
rect 203576 237408 203984 237436
rect 203576 237396 203582 237408
rect 203978 237396 203984 237408
rect 204036 237396 204042 237448
rect 208394 237396 208400 237448
rect 208452 237436 208458 237448
rect 210326 237436 210332 237448
rect 208452 237408 210332 237436
rect 208452 237396 208458 237408
rect 210326 237396 210332 237408
rect 210384 237396 210390 237448
rect 211798 237396 211804 237448
rect 211856 237436 211862 237448
rect 212442 237436 212448 237448
rect 211856 237408 212448 237436
rect 211856 237396 211862 237408
rect 212442 237396 212448 237408
rect 212500 237396 212506 237448
rect 213086 237396 213092 237448
rect 213144 237436 213150 237448
rect 213730 237436 213736 237448
rect 213144 237408 213736 237436
rect 213144 237396 213150 237408
rect 213730 237396 213736 237408
rect 213788 237396 213794 237448
rect 215662 237396 215668 237448
rect 215720 237436 215726 237448
rect 216582 237436 216588 237448
rect 215720 237408 216588 237436
rect 215720 237396 215726 237408
rect 216582 237396 216588 237408
rect 216640 237396 216646 237448
rect 218422 237396 218428 237448
rect 218480 237436 218486 237448
rect 219250 237436 219256 237448
rect 218480 237408 219256 237436
rect 218480 237396 218486 237408
rect 219250 237396 219256 237408
rect 219308 237396 219314 237448
rect 219894 237396 219900 237448
rect 219952 237436 219958 237448
rect 220722 237436 220728 237448
rect 219952 237408 220728 237436
rect 219952 237396 219958 237408
rect 220722 237396 220728 237408
rect 220780 237396 220786 237448
rect 220998 237396 221004 237448
rect 221056 237436 221062 237448
rect 222010 237436 222016 237448
rect 221056 237408 222016 237436
rect 221056 237396 221062 237408
rect 222010 237396 222016 237408
rect 222068 237396 222074 237448
rect 225782 237396 225788 237448
rect 225840 237436 225846 237448
rect 226242 237436 226248 237448
rect 225840 237408 226248 237436
rect 225840 237396 225846 237408
rect 226242 237396 226248 237408
rect 226300 237396 226306 237448
rect 226702 237396 226708 237448
rect 226760 237436 226766 237448
rect 227622 237436 227628 237448
rect 226760 237408 227628 237436
rect 226760 237396 226766 237408
rect 227622 237396 227628 237408
rect 227680 237396 227686 237448
rect 232038 237396 232044 237448
rect 232096 237436 232102 237448
rect 233142 237436 233148 237448
rect 232096 237408 233148 237436
rect 232096 237396 232102 237408
rect 233142 237396 233148 237408
rect 233200 237396 233206 237448
rect 236822 237396 236828 237448
rect 236880 237436 236886 237448
rect 237282 237436 237288 237448
rect 236880 237408 237288 237436
rect 236880 237396 236886 237408
rect 237282 237396 237288 237408
rect 237340 237396 237346 237448
rect 237374 237396 237380 237448
rect 237432 237436 237438 237448
rect 238662 237436 238668 237448
rect 237432 237408 238668 237436
rect 237432 237396 237438 237408
rect 238662 237396 238668 237408
rect 238720 237396 238726 237448
rect 240318 237396 240324 237448
rect 240376 237436 240382 237448
rect 241422 237436 241428 237448
rect 240376 237408 241428 237436
rect 240376 237396 240382 237408
rect 241422 237396 241428 237408
rect 241480 237396 241486 237448
rect 41322 237328 41328 237380
rect 41380 237368 41386 237380
rect 219526 237368 219532 237380
rect 41380 237340 219532 237368
rect 41380 237328 41386 237340
rect 219526 237328 219532 237340
rect 219584 237328 219590 237380
rect 221366 237328 221372 237380
rect 221424 237368 221430 237380
rect 363598 237368 363604 237380
rect 221424 237340 363604 237368
rect 221424 237328 221430 237340
rect 363598 237328 363604 237340
rect 363656 237328 363662 237380
rect 235258 236784 235264 236836
rect 235316 236824 235322 236836
rect 243262 236824 243268 236836
rect 235316 236796 243268 236824
rect 235316 236784 235322 236796
rect 243262 236784 243268 236796
rect 243320 236784 243326 236836
rect 217134 236648 217140 236700
rect 217192 236688 217198 236700
rect 232130 236688 232136 236700
rect 217192 236660 232136 236688
rect 217192 236648 217198 236660
rect 232130 236648 232136 236660
rect 232188 236648 232194 236700
rect 235350 236648 235356 236700
rect 235408 236688 235414 236700
rect 582650 236688 582656 236700
rect 235408 236660 582656 236688
rect 235408 236648 235414 236660
rect 582650 236648 582656 236660
rect 582708 236648 582714 236700
rect 240502 236104 240508 236156
rect 240560 236144 240566 236156
rect 240962 236144 240968 236156
rect 240560 236116 240968 236144
rect 240560 236104 240566 236116
rect 240962 236104 240968 236116
rect 241020 236104 241026 236156
rect 202046 235900 202052 235952
rect 202104 235940 202110 235952
rect 305638 235940 305644 235952
rect 202104 235912 305644 235940
rect 202104 235900 202110 235912
rect 305638 235900 305644 235912
rect 305696 235900 305702 235952
rect 230198 235396 230204 235408
rect 219406 235368 230204 235396
rect 22738 235288 22744 235340
rect 22796 235328 22802 235340
rect 219406 235328 219434 235368
rect 230198 235356 230204 235368
rect 230256 235356 230262 235408
rect 22796 235300 219434 235328
rect 22796 235288 22802 235300
rect 229094 235288 229100 235340
rect 229152 235328 229158 235340
rect 295426 235328 295432 235340
rect 229152 235300 295432 235328
rect 229152 235288 229158 235300
rect 295426 235288 295432 235300
rect 295484 235288 295490 235340
rect 212166 235220 212172 235272
rect 212224 235260 212230 235272
rect 582466 235260 582472 235272
rect 212224 235232 582472 235260
rect 212224 235220 212230 235232
rect 582466 235220 582472 235232
rect 582524 235220 582530 235272
rect 243630 234064 243636 234116
rect 243688 234104 243694 234116
rect 293954 234104 293960 234116
rect 243688 234076 293960 234104
rect 243688 234064 243694 234076
rect 293954 234064 293960 234076
rect 294012 234064 294018 234116
rect 227254 233996 227260 234048
rect 227312 234036 227318 234048
rect 289814 234036 289820 234048
rect 227312 234008 289820 234036
rect 227312 233996 227318 234008
rect 289814 233996 289820 234008
rect 289872 233996 289878 234048
rect 170398 233928 170404 233980
rect 170456 233968 170462 233980
rect 245746 233968 245752 233980
rect 170456 233940 245752 233968
rect 170456 233928 170462 233940
rect 245746 233928 245752 233940
rect 245804 233928 245810 233980
rect 3418 233860 3424 233912
rect 3476 233900 3482 233912
rect 208394 233900 208400 233912
rect 3476 233872 208400 233900
rect 3476 233860 3482 233872
rect 208394 233860 208400 233872
rect 208452 233860 208458 233912
rect 209866 233860 209872 233912
rect 209924 233900 209930 233912
rect 582742 233900 582748 233912
rect 209924 233872 582748 233900
rect 209924 233860 209930 233872
rect 582742 233860 582748 233872
rect 582800 233860 582806 233912
rect 239398 233520 239404 233572
rect 239456 233560 239462 233572
rect 242158 233560 242164 233572
rect 239456 233532 242164 233560
rect 239456 233520 239462 233532
rect 242158 233520 242164 233532
rect 242216 233520 242222 233572
rect 231118 233180 231124 233232
rect 231176 233220 231182 233232
rect 233326 233220 233332 233232
rect 231176 233192 233332 233220
rect 231176 233180 231182 233192
rect 233326 233180 233332 233192
rect 233384 233180 233390 233232
rect 195606 232568 195612 232620
rect 195664 232608 195670 232620
rect 303706 232608 303712 232620
rect 195664 232580 303712 232608
rect 195664 232568 195670 232580
rect 303706 232568 303712 232580
rect 303764 232568 303770 232620
rect 4798 232500 4804 232552
rect 4856 232540 4862 232552
rect 229646 232540 229652 232552
rect 4856 232512 229652 232540
rect 4856 232500 4862 232512
rect 229646 232500 229652 232512
rect 229704 232500 229710 232552
rect 222286 231140 222292 231192
rect 222344 231180 222350 231192
rect 278038 231180 278044 231192
rect 222344 231152 278044 231180
rect 222344 231140 222350 231152
rect 278038 231140 278044 231152
rect 278096 231140 278102 231192
rect 204990 231072 204996 231124
rect 205048 231112 205054 231124
rect 582558 231112 582564 231124
rect 205048 231084 582564 231112
rect 205048 231072 205054 231084
rect 582558 231072 582564 231084
rect 582616 231072 582622 231124
rect 178678 229848 178684 229900
rect 178736 229888 178742 229900
rect 245654 229888 245660 229900
rect 178736 229860 245660 229888
rect 178736 229848 178742 229860
rect 245654 229848 245660 229860
rect 245712 229848 245718 229900
rect 218974 229780 218980 229832
rect 219032 229820 219038 229832
rect 288710 229820 288716 229832
rect 219032 229792 288716 229820
rect 219032 229780 219038 229792
rect 288710 229780 288716 229792
rect 288768 229780 288774 229832
rect 194318 229712 194324 229764
rect 194376 229752 194382 229764
rect 298278 229752 298284 229764
rect 194376 229724 298284 229752
rect 194376 229712 194382 229724
rect 298278 229712 298284 229724
rect 298336 229712 298342 229764
rect 241330 228420 241336 228472
rect 241388 228460 241394 228472
rect 291286 228460 291292 228472
rect 241388 228432 291292 228460
rect 241388 228420 241394 228432
rect 291286 228420 291292 228432
rect 291344 228420 291350 228472
rect 196986 228352 196992 228404
rect 197044 228392 197050 228404
rect 276842 228392 276848 228404
rect 197044 228364 276848 228392
rect 197044 228352 197050 228364
rect 276842 228352 276848 228364
rect 276900 228352 276906 228404
rect 222010 227060 222016 227112
rect 222068 227100 222074 227112
rect 302326 227100 302332 227112
rect 222068 227072 302332 227100
rect 222068 227060 222074 227072
rect 302326 227060 302332 227072
rect 302384 227060 302390 227112
rect 203978 226992 203984 227044
rect 204036 227032 204042 227044
rect 292574 227032 292580 227044
rect 204036 227004 292580 227032
rect 204036 226992 204042 227004
rect 292574 226992 292580 227004
rect 292632 226992 292638 227044
rect 226150 225564 226156 225616
rect 226208 225604 226214 225616
rect 305086 225604 305092 225616
rect 226208 225576 305092 225604
rect 226208 225564 226214 225576
rect 305086 225564 305092 225576
rect 305144 225564 305150 225616
rect 220722 224204 220728 224256
rect 220780 224244 220786 224256
rect 282178 224244 282184 224256
rect 220780 224216 282184 224244
rect 220780 224204 220786 224216
rect 282178 224204 282184 224216
rect 282236 224204 282242 224256
rect 352558 224204 352564 224256
rect 352616 224244 352622 224256
rect 580258 224244 580264 224256
rect 352616 224216 580264 224244
rect 352616 224204 352622 224216
rect 580258 224204 580264 224216
rect 580316 224204 580322 224256
rect 202690 221416 202696 221468
rect 202748 221456 202754 221468
rect 285766 221456 285772 221468
rect 202748 221428 285772 221456
rect 202748 221416 202754 221428
rect 285766 221416 285772 221428
rect 285824 221416 285830 221468
rect 224678 218696 224684 218748
rect 224736 218736 224742 218748
rect 299658 218736 299664 218748
rect 224736 218708 299664 218736
rect 224736 218696 224742 218708
rect 299658 218696 299664 218708
rect 299716 218696 299722 218748
rect 201310 215908 201316 215960
rect 201368 215948 201374 215960
rect 296806 215948 296812 215960
rect 201368 215920 296812 215948
rect 201368 215908 201374 215920
rect 296806 215908 296812 215920
rect 296864 215908 296870 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 15838 215268 15844 215280
rect 3384 215240 15844 215268
rect 3384 215228 3390 215240
rect 15838 215228 15844 215240
rect 15896 215228 15902 215280
rect 233142 213188 233148 213240
rect 233200 213228 233206 213240
rect 288526 213228 288532 213240
rect 233200 213200 288532 213228
rect 233200 213188 233206 213200
rect 288526 213188 288532 213200
rect 288584 213188 288590 213240
rect 188798 211760 188804 211812
rect 188856 211800 188862 211812
rect 296714 211800 296720 211812
rect 188856 211772 296720 211800
rect 188856 211760 188862 211772
rect 296714 211760 296720 211772
rect 296772 211760 296778 211812
rect 208210 210400 208216 210452
rect 208268 210440 208274 210452
rect 280154 210440 280160 210452
rect 208268 210412 280160 210440
rect 208268 210400 208274 210412
rect 280154 210400 280160 210412
rect 280212 210400 280218 210452
rect 191466 209040 191472 209092
rect 191524 209080 191530 209092
rect 582834 209080 582840 209092
rect 191524 209052 582840 209080
rect 191524 209040 191530 209052
rect 582834 209040 582840 209052
rect 582892 209040 582898 209092
rect 302878 206932 302884 206984
rect 302936 206972 302942 206984
rect 579798 206972 579804 206984
rect 302936 206944 579804 206972
rect 302936 206932 302942 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 219250 204892 219256 204944
rect 219308 204932 219314 204944
rect 284386 204932 284392 204944
rect 219308 204904 284392 204932
rect 219308 204892 219314 204904
rect 284386 204892 284392 204904
rect 284444 204892 284450 204944
rect 209130 203600 209136 203652
rect 209188 203640 209194 203652
rect 214558 203640 214564 203652
rect 209188 203612 214564 203640
rect 209188 203600 209194 203612
rect 214558 203600 214564 203612
rect 214616 203600 214622 203652
rect 205450 203532 205456 203584
rect 205508 203572 205514 203584
rect 289906 203572 289912 203584
rect 205508 203544 289912 203572
rect 205508 203532 205514 203544
rect 289906 203532 289912 203544
rect 289964 203532 289970 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 170398 202824 170404 202836
rect 3108 202796 170404 202824
rect 3108 202784 3114 202796
rect 170398 202784 170404 202796
rect 170456 202784 170462 202836
rect 215018 202104 215024 202156
rect 215076 202144 215082 202156
rect 307846 202144 307852 202156
rect 215076 202116 307852 202144
rect 215076 202104 215082 202116
rect 307846 202104 307852 202116
rect 307904 202104 307910 202156
rect 233878 201832 233884 201884
rect 233936 201872 233942 201884
rect 237926 201872 237932 201884
rect 233936 201844 237932 201872
rect 233936 201832 233942 201844
rect 237926 201832 237932 201844
rect 237984 201832 237990 201884
rect 204898 200744 204904 200796
rect 204956 200784 204962 200796
rect 299566 200784 299572 200796
rect 204956 200756 299572 200784
rect 204956 200744 204962 200756
rect 299566 200744 299572 200756
rect 299624 200744 299630 200796
rect 220170 199384 220176 199436
rect 220228 199424 220234 199436
rect 230750 199424 230756 199436
rect 220228 199396 230756 199424
rect 220228 199384 220234 199396
rect 230750 199384 230756 199396
rect 230808 199384 230814 199436
rect 227622 197956 227628 198008
rect 227680 197996 227686 198008
rect 291378 197996 291384 198008
rect 227680 197968 291384 197996
rect 227680 197956 227686 197968
rect 291378 197956 291384 197968
rect 291436 197956 291442 198008
rect 198458 196596 198464 196648
rect 198516 196636 198522 196648
rect 279050 196636 279056 196648
rect 198516 196608 279056 196636
rect 198516 196596 198522 196608
rect 279050 196596 279056 196608
rect 279108 196596 279114 196648
rect 199838 195304 199844 195356
rect 199896 195344 199902 195356
rect 245654 195344 245660 195356
rect 199896 195316 245660 195344
rect 199896 195304 199902 195316
rect 245654 195304 245660 195316
rect 245712 195304 245718 195356
rect 217870 195236 217876 195288
rect 217928 195276 217934 195288
rect 300946 195276 300952 195288
rect 217928 195248 300952 195276
rect 217928 195236 217934 195248
rect 300946 195236 300952 195248
rect 301004 195236 301010 195288
rect 180610 193808 180616 193860
rect 180668 193848 180674 193860
rect 271322 193848 271328 193860
rect 180668 193820 271328 193848
rect 180668 193808 180674 193820
rect 271322 193808 271328 193820
rect 271380 193808 271386 193860
rect 334618 193128 334624 193180
rect 334676 193168 334682 193180
rect 580166 193168 580172 193180
rect 334676 193140 580172 193168
rect 334676 193128 334682 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 187602 192516 187608 192568
rect 187660 192556 187666 192568
rect 242894 192556 242900 192568
rect 187660 192528 242900 192556
rect 187660 192516 187666 192528
rect 242894 192516 242900 192528
rect 242952 192516 242958 192568
rect 220078 192448 220084 192500
rect 220136 192488 220142 192500
rect 292758 192488 292764 192500
rect 220136 192460 292764 192488
rect 220136 192448 220142 192460
rect 292758 192448 292764 192460
rect 292816 192448 292822 192500
rect 214558 189932 214564 189984
rect 214616 189972 214622 189984
rect 240410 189972 240416 189984
rect 214616 189944 240416 189972
rect 214616 189932 214622 189944
rect 240410 189932 240416 189944
rect 240468 189932 240474 189984
rect 182082 189864 182088 189916
rect 182140 189904 182146 189916
rect 228358 189904 228364 189916
rect 182140 189876 228364 189904
rect 182140 189864 182146 189876
rect 228358 189864 228364 189876
rect 228416 189864 228422 189916
rect 197170 189796 197176 189848
rect 197228 189836 197234 189848
rect 278774 189836 278780 189848
rect 197228 189808 278780 189836
rect 197228 189796 197234 189808
rect 278774 189796 278780 189808
rect 278832 189796 278838 189848
rect 192938 189728 192944 189780
rect 192996 189768 193002 189780
rect 302418 189768 302424 189780
rect 192996 189740 302424 189768
rect 192996 189728 193002 189740
rect 302418 189728 302424 189740
rect 302476 189728 302482 189780
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 173158 189020 173164 189032
rect 3568 188992 173164 189020
rect 3568 188980 3574 188992
rect 173158 188980 173164 188992
rect 173216 188980 173222 189032
rect 195698 188368 195704 188420
rect 195756 188408 195762 188420
rect 230566 188408 230572 188420
rect 195756 188380 230572 188408
rect 195756 188368 195762 188380
rect 230566 188368 230572 188380
rect 230624 188368 230630 188420
rect 203886 188300 203892 188352
rect 203944 188340 203950 188352
rect 285858 188340 285864 188352
rect 203944 188312 285864 188340
rect 203944 188300 203950 188312
rect 285858 188300 285864 188312
rect 285916 188300 285922 188352
rect 204162 187076 204168 187128
rect 204220 187116 204226 187128
rect 244458 187116 244464 187128
rect 204220 187088 244464 187116
rect 204220 187076 204226 187088
rect 244458 187076 244464 187088
rect 244516 187076 244522 187128
rect 188706 187008 188712 187060
rect 188764 187048 188770 187060
rect 248506 187048 248512 187060
rect 188764 187020 248512 187048
rect 188764 187008 188770 187020
rect 248506 187008 248512 187020
rect 248564 187008 248570 187060
rect 193030 186940 193036 186992
rect 193088 186980 193094 186992
rect 287238 186980 287244 186992
rect 193088 186952 287244 186980
rect 193088 186940 193094 186952
rect 287238 186940 287244 186952
rect 287296 186940 287302 186992
rect 261478 185648 261484 185700
rect 261536 185688 261542 185700
rect 291470 185688 291476 185700
rect 261536 185660 291476 185688
rect 261536 185648 261542 185660
rect 291470 185648 291476 185660
rect 291528 185648 291534 185700
rect 226242 185580 226248 185632
rect 226300 185620 226306 185632
rect 226300 185592 277394 185620
rect 226300 185580 226306 185592
rect 277366 185552 277394 185592
rect 282178 185580 282184 185632
rect 282236 185620 282242 185632
rect 285950 185620 285956 185632
rect 282236 185592 285956 185620
rect 282236 185580 282242 185592
rect 285950 185580 285956 185592
rect 286008 185580 286014 185632
rect 284478 185552 284484 185564
rect 277366 185524 284484 185552
rect 284478 185512 284484 185524
rect 284536 185512 284542 185564
rect 213822 184492 213828 184544
rect 213880 184532 213886 184544
rect 242986 184532 242992 184544
rect 213880 184504 242992 184532
rect 213880 184492 213886 184504
rect 242986 184492 242992 184504
rect 243044 184492 243050 184544
rect 206830 184424 206836 184476
rect 206888 184464 206894 184476
rect 235994 184464 236000 184476
rect 206888 184436 236000 184464
rect 206888 184424 206894 184436
rect 235994 184424 236000 184436
rect 236052 184424 236058 184476
rect 197078 184356 197084 184408
rect 197136 184396 197142 184408
rect 240134 184396 240140 184408
rect 197136 184368 240140 184396
rect 197136 184356 197142 184368
rect 240134 184356 240140 184368
rect 240192 184356 240198 184408
rect 240410 184356 240416 184408
rect 240468 184396 240474 184408
rect 278130 184396 278136 184408
rect 240468 184368 278136 184396
rect 240468 184356 240474 184368
rect 278130 184356 278136 184368
rect 278188 184356 278194 184408
rect 199930 184288 199936 184340
rect 199988 184328 199994 184340
rect 245746 184328 245752 184340
rect 199988 184300 245752 184328
rect 199988 184288 199994 184300
rect 245746 184288 245752 184300
rect 245804 184288 245810 184340
rect 229002 184220 229008 184272
rect 229060 184260 229066 184272
rect 302510 184260 302516 184272
rect 229060 184232 302516 184260
rect 229060 184220 229066 184232
rect 302510 184220 302516 184232
rect 302568 184220 302574 184272
rect 191650 184152 191656 184204
rect 191708 184192 191714 184204
rect 290090 184192 290096 184204
rect 191708 184164 290096 184192
rect 191708 184152 191714 184164
rect 290090 184152 290096 184164
rect 290148 184152 290154 184204
rect 272518 182860 272524 182912
rect 272576 182900 272582 182912
rect 298370 182900 298376 182912
rect 272576 182872 298376 182900
rect 272576 182860 272582 182872
rect 298370 182860 298376 182872
rect 298428 182860 298434 182912
rect 246390 182792 246396 182844
rect 246448 182832 246454 182844
rect 287146 182832 287152 182844
rect 246448 182804 287152 182832
rect 246448 182792 246454 182804
rect 287146 182792 287152 182804
rect 287204 182792 287210 182844
rect 262858 181704 262864 181756
rect 262916 181744 262922 181756
rect 281534 181744 281540 181756
rect 262916 181716 281540 181744
rect 262916 181704 262922 181716
rect 281534 181704 281540 181716
rect 281592 181704 281598 181756
rect 183462 181636 183468 181688
rect 183520 181676 183526 181688
rect 241606 181676 241612 181688
rect 183520 181648 241612 181676
rect 183520 181636 183526 181648
rect 241606 181636 241612 181648
rect 241664 181636 241670 181688
rect 266998 181636 267004 181688
rect 267056 181676 267062 181688
rect 296898 181676 296904 181688
rect 267056 181648 296904 181676
rect 267056 181636 267062 181648
rect 296898 181636 296904 181648
rect 296956 181636 296962 181688
rect 187418 181568 187424 181620
rect 187476 181608 187482 181620
rect 247218 181608 247224 181620
rect 187476 181580 247224 181608
rect 187476 181568 187482 181580
rect 247218 181568 247224 181580
rect 247276 181568 247282 181620
rect 253198 181568 253204 181620
rect 253256 181608 253262 181620
rect 295610 181608 295616 181620
rect 253256 181580 295616 181608
rect 253256 181568 253262 181580
rect 295610 181568 295616 181580
rect 295668 181568 295674 181620
rect 234522 181500 234528 181552
rect 234580 181540 234586 181552
rect 303798 181540 303804 181552
rect 234580 181512 303804 181540
rect 234580 181500 234586 181512
rect 303798 181500 303804 181512
rect 303856 181500 303862 181552
rect 202598 181432 202604 181484
rect 202656 181472 202662 181484
rect 283466 181472 283472 181484
rect 202656 181444 283472 181472
rect 202656 181432 202662 181444
rect 283466 181432 283472 181444
rect 283524 181432 283530 181484
rect 130930 181024 130936 181076
rect 130988 181064 130994 181076
rect 173250 181064 173256 181076
rect 130988 181036 173256 181064
rect 130988 181024 130994 181036
rect 173250 181024 173256 181036
rect 173308 181024 173314 181076
rect 128170 180956 128176 181008
rect 128228 180996 128234 181008
rect 184382 180996 184388 181008
rect 128228 180968 184388 180996
rect 128228 180956 128234 180968
rect 184382 180956 184388 180968
rect 184440 180956 184446 181008
rect 102042 180888 102048 180940
rect 102100 180928 102106 180940
rect 169018 180928 169024 180940
rect 102100 180900 169024 180928
rect 102100 180888 102106 180900
rect 169018 180888 169024 180900
rect 169076 180888 169082 180940
rect 99466 180820 99472 180872
rect 99524 180860 99530 180872
rect 203518 180860 203524 180872
rect 99524 180832 203524 180860
rect 99524 180820 99530 180832
rect 203518 180820 203524 180832
rect 203576 180820 203582 180872
rect 273898 180276 273904 180328
rect 273956 180316 273962 180328
rect 294138 180316 294144 180328
rect 273956 180288 294144 180316
rect 273956 180276 273962 180288
rect 294138 180276 294144 180288
rect 294196 180276 294202 180328
rect 215202 180208 215208 180260
rect 215260 180248 215266 180260
rect 237558 180248 237564 180260
rect 215260 180220 237564 180248
rect 215260 180208 215266 180220
rect 237558 180208 237564 180220
rect 237616 180208 237622 180260
rect 260098 180208 260104 180260
rect 260156 180248 260162 180260
rect 292666 180248 292672 180260
rect 260156 180220 292672 180248
rect 260156 180208 260162 180220
rect 292666 180208 292672 180220
rect 292724 180208 292730 180260
rect 200022 180140 200028 180192
rect 200080 180180 200086 180192
rect 230658 180180 230664 180192
rect 200080 180152 230664 180180
rect 200080 180140 200086 180152
rect 230658 180140 230664 180152
rect 230716 180140 230722 180192
rect 237282 180140 237288 180192
rect 237340 180180 237346 180192
rect 283190 180180 283196 180192
rect 237340 180152 283196 180180
rect 237340 180140 237346 180152
rect 283190 180140 283196 180152
rect 283248 180140 283254 180192
rect 201402 180072 201408 180124
rect 201460 180112 201466 180124
rect 292850 180112 292856 180124
rect 201460 180084 292856 180112
rect 201460 180072 201466 180084
rect 292850 180072 292856 180084
rect 292908 180072 292914 180124
rect 129458 179732 129464 179784
rect 129516 179772 129522 179784
rect 168374 179772 168380 179784
rect 129516 179744 168380 179772
rect 129516 179732 129522 179744
rect 168374 179732 168380 179744
rect 168432 179732 168438 179784
rect 123294 179664 123300 179716
rect 123352 179704 123358 179716
rect 175918 179704 175924 179716
rect 123352 179676 175924 179704
rect 123352 179664 123358 179676
rect 175918 179664 175924 179676
rect 175976 179664 175982 179716
rect 121270 179596 121276 179648
rect 121328 179636 121334 179648
rect 177390 179636 177396 179648
rect 121328 179608 177396 179636
rect 121328 179596 121334 179608
rect 177390 179596 177396 179608
rect 177448 179596 177454 179648
rect 110690 179528 110696 179580
rect 110748 179568 110754 179580
rect 182818 179568 182824 179580
rect 110748 179540 182824 179568
rect 110748 179528 110754 179540
rect 182818 179528 182824 179540
rect 182876 179528 182882 179580
rect 108114 179460 108120 179512
rect 108172 179500 108178 179512
rect 181438 179500 181444 179512
rect 108172 179472 181444 179500
rect 108172 179460 108178 179472
rect 181438 179460 181444 179472
rect 181496 179460 181502 179512
rect 114554 179392 114560 179444
rect 114612 179432 114618 179444
rect 214558 179432 214564 179444
rect 114612 179404 214564 179432
rect 114612 179392 114618 179404
rect 214558 179392 214564 179404
rect 214616 179392 214622 179444
rect 224770 178984 224776 179036
rect 224828 179024 224834 179036
rect 231946 179024 231952 179036
rect 224828 178996 231952 179024
rect 224828 178984 224834 178996
rect 231946 178984 231952 178996
rect 232004 178984 232010 179036
rect 269942 178984 269948 179036
rect 270000 179024 270006 179036
rect 284570 179024 284576 179036
rect 270000 178996 284576 179024
rect 270000 178984 270006 178996
rect 284570 178984 284576 178996
rect 284628 178984 284634 179036
rect 212442 178916 212448 178968
rect 212500 178956 212506 178968
rect 229462 178956 229468 178968
rect 212500 178928 229468 178956
rect 212500 178916 212506 178928
rect 229462 178916 229468 178928
rect 229520 178916 229526 178968
rect 268378 178916 268384 178968
rect 268436 178956 268442 178968
rect 289998 178956 290004 178968
rect 268436 178928 290004 178956
rect 268436 178916 268442 178928
rect 289998 178916 290004 178928
rect 290056 178916 290062 178968
rect 206922 178848 206928 178900
rect 206980 178888 206986 178900
rect 237466 178888 237472 178900
rect 206980 178860 237472 178888
rect 206980 178848 206986 178860
rect 237466 178848 237472 178860
rect 237524 178848 237530 178900
rect 271230 178848 271236 178900
rect 271288 178888 271294 178900
rect 296990 178888 296996 178900
rect 271288 178860 296996 178888
rect 271288 178848 271294 178860
rect 296990 178848 296996 178860
rect 297048 178848 297054 178900
rect 195790 178780 195796 178832
rect 195848 178820 195854 178832
rect 236086 178820 236092 178832
rect 195848 178792 236092 178820
rect 195848 178780 195854 178792
rect 236086 178780 236092 178792
rect 236144 178780 236150 178832
rect 267090 178780 267096 178832
rect 267148 178820 267154 178832
rect 295518 178820 295524 178832
rect 267148 178792 295524 178820
rect 267148 178780 267154 178792
rect 295518 178780 295524 178792
rect 295576 178780 295582 178832
rect 186130 178712 186136 178764
rect 186188 178752 186194 178764
rect 229186 178752 229192 178764
rect 186188 178724 229192 178752
rect 186188 178712 186194 178724
rect 229186 178712 229192 178724
rect 229244 178712 229250 178764
rect 241422 178712 241428 178764
rect 241480 178752 241486 178764
rect 279234 178752 279240 178764
rect 241480 178724 279240 178752
rect 241480 178712 241486 178724
rect 279234 178712 279240 178724
rect 279292 178712 279298 178764
rect 184750 178644 184756 178696
rect 184808 178684 184814 178696
rect 236178 178684 236184 178696
rect 184808 178656 236184 178684
rect 184808 178644 184814 178656
rect 236178 178644 236184 178656
rect 236236 178644 236242 178696
rect 238662 178644 238668 178696
rect 238720 178684 238726 178696
rect 283374 178684 283380 178696
rect 238720 178656 283380 178684
rect 238720 178644 238726 178656
rect 283374 178644 283380 178656
rect 283432 178644 283438 178696
rect 132402 178372 132408 178424
rect 132460 178412 132466 178424
rect 165338 178412 165344 178424
rect 132460 178384 165344 178412
rect 132460 178372 132466 178384
rect 165338 178372 165344 178384
rect 165396 178372 165402 178424
rect 112254 178304 112260 178356
rect 112312 178344 112318 178356
rect 166350 178344 166356 178356
rect 112312 178316 166356 178344
rect 112312 178304 112318 178316
rect 166350 178304 166356 178316
rect 166408 178304 166414 178356
rect 116946 178236 116952 178288
rect 117004 178276 117010 178288
rect 174538 178276 174544 178288
rect 117004 178248 174544 178276
rect 117004 178236 117010 178248
rect 174538 178236 174544 178248
rect 174596 178236 174602 178288
rect 125962 178168 125968 178220
rect 126020 178208 126026 178220
rect 186958 178208 186964 178220
rect 126020 178180 186964 178208
rect 126020 178168 126026 178180
rect 186958 178168 186964 178180
rect 187016 178168 187022 178220
rect 109586 178100 109592 178152
rect 109644 178140 109650 178152
rect 180058 178140 180064 178152
rect 109644 178112 180064 178140
rect 109644 178100 109650 178112
rect 180058 178100 180064 178112
rect 180116 178100 180122 178152
rect 119522 178032 119528 178084
rect 119580 178072 119586 178084
rect 200758 178072 200764 178084
rect 119580 178044 200764 178072
rect 119580 178032 119586 178044
rect 200758 178032 200764 178044
rect 200816 178032 200822 178084
rect 223390 177964 223396 178016
rect 223448 178004 223454 178016
rect 229370 178004 229376 178016
rect 223448 177976 229376 178004
rect 223448 177964 223454 177976
rect 229370 177964 229376 177976
rect 229428 177964 229434 178016
rect 271322 177556 271328 177608
rect 271380 177596 271386 177608
rect 288434 177596 288440 177608
rect 271380 177568 288440 177596
rect 271380 177556 271386 177568
rect 288434 177556 288440 177568
rect 288492 177556 288498 177608
rect 278130 177488 278136 177540
rect 278188 177528 278194 177540
rect 301038 177528 301044 177540
rect 278188 177500 301044 177528
rect 278188 177488 278194 177500
rect 301038 177488 301044 177500
rect 301096 177488 301102 177540
rect 219342 177420 219348 177472
rect 219400 177460 219406 177472
rect 234798 177460 234804 177472
rect 219400 177432 234804 177460
rect 219400 177420 219406 177432
rect 234798 177420 234804 177432
rect 234856 177420 234862 177472
rect 269850 177420 269856 177472
rect 269908 177460 269914 177472
rect 294230 177460 294236 177472
rect 269908 177432 294236 177460
rect 269908 177420 269914 177432
rect 294230 177420 294236 177432
rect 294288 177420 294294 177472
rect 208302 177352 208308 177404
rect 208360 177392 208366 177404
rect 279142 177392 279148 177404
rect 208360 177364 279148 177392
rect 208360 177352 208366 177364
rect 279142 177352 279148 177364
rect 279200 177352 279206 177404
rect 198642 177284 198648 177336
rect 198700 177324 198706 177336
rect 280338 177324 280344 177336
rect 198700 177296 280344 177324
rect 198700 177284 198706 177296
rect 280338 177284 280344 177296
rect 280396 177284 280402 177336
rect 105722 177080 105728 177132
rect 105780 177120 105786 177132
rect 191098 177120 191104 177132
rect 105780 177092 191104 177120
rect 105780 177080 105786 177092
rect 191098 177080 191104 177092
rect 191156 177080 191162 177132
rect 134426 177012 134432 177064
rect 134484 177052 134490 177064
rect 165430 177052 165436 177064
rect 134484 177024 165436 177052
rect 134484 177012 134490 177024
rect 165430 177012 165436 177024
rect 165488 177012 165494 177064
rect 127158 176944 127164 176996
rect 127216 176984 127222 176996
rect 167730 176984 167736 176996
rect 127216 176956 167736 176984
rect 127216 176944 127222 176956
rect 167730 176944 167736 176956
rect 167788 176944 167794 176996
rect 158898 176876 158904 176928
rect 158956 176916 158962 176928
rect 207658 176916 207664 176928
rect 158956 176888 207664 176916
rect 158956 176876 158962 176888
rect 207658 176876 207664 176888
rect 207716 176876 207722 176928
rect 148226 176808 148232 176860
rect 148284 176848 148290 176860
rect 198090 176848 198096 176860
rect 148284 176820 198096 176848
rect 148284 176808 148290 176820
rect 198090 176808 198096 176820
rect 198148 176808 198154 176860
rect 107010 176740 107016 176792
rect 107068 176780 107074 176792
rect 170490 176780 170496 176792
rect 107068 176752 170496 176780
rect 107068 176740 107074 176752
rect 170490 176740 170496 176752
rect 170548 176740 170554 176792
rect 136082 176672 136088 176724
rect 136140 176712 136146 176724
rect 136140 176684 136772 176712
rect 136140 176672 136146 176684
rect 136744 176644 136772 176684
rect 213914 176644 213920 176656
rect 136744 176616 213920 176644
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 276842 176604 276848 176656
rect 276900 176644 276906 176656
rect 283006 176644 283012 176656
rect 276900 176616 283012 176644
rect 276900 176604 276906 176616
rect 283006 176604 283012 176616
rect 283064 176604 283070 176656
rect 191558 176536 191564 176588
rect 191616 176576 191622 176588
rect 241514 176576 241520 176588
rect 191616 176548 241520 176576
rect 191616 176536 191622 176548
rect 241514 176536 241520 176548
rect 241572 176536 241578 176588
rect 280798 176536 280804 176588
rect 280856 176576 280862 176588
rect 287330 176576 287336 176588
rect 280856 176548 287336 176576
rect 280856 176536 280862 176548
rect 287330 176536 287336 176548
rect 287388 176536 287394 176588
rect 278038 176468 278044 176520
rect 278096 176508 278102 176520
rect 280246 176508 280252 176520
rect 278096 176480 280252 176508
rect 278096 176468 278102 176480
rect 280246 176468 280252 176480
rect 280304 176468 280310 176520
rect 133138 176196 133144 176248
rect 133196 176236 133202 176248
rect 165522 176236 165528 176248
rect 133196 176208 165528 176236
rect 133196 176196 133202 176208
rect 165522 176196 165528 176208
rect 165580 176196 165586 176248
rect 124490 176128 124496 176180
rect 124548 176168 124554 176180
rect 166442 176168 166448 176180
rect 124548 176140 166448 176168
rect 124548 176128 124554 176140
rect 166442 176128 166448 176140
rect 166500 176128 166506 176180
rect 276750 176128 276756 176180
rect 276808 176168 276814 176180
rect 279326 176168 279332 176180
rect 276808 176140 279332 176168
rect 276808 176128 276814 176140
rect 279326 176128 279332 176140
rect 279384 176128 279390 176180
rect 121914 176060 121920 176112
rect 121972 176100 121978 176112
rect 169110 176100 169116 176112
rect 121972 176072 169116 176100
rect 121972 176060 121978 176072
rect 169110 176060 169116 176072
rect 169168 176060 169174 176112
rect 224862 176060 224868 176112
rect 224920 176100 224926 176112
rect 231854 176100 231860 176112
rect 224920 176072 231860 176100
rect 224920 176060 224926 176072
rect 231854 176060 231860 176072
rect 231912 176060 231918 176112
rect 276658 176060 276664 176112
rect 276716 176100 276722 176112
rect 280430 176100 280436 176112
rect 276716 176072 280436 176100
rect 276716 176060 276722 176072
rect 280430 176060 280436 176072
rect 280488 176060 280494 176112
rect 118418 175992 118424 176044
rect 118476 176032 118482 176044
rect 173158 176032 173164 176044
rect 118476 176004 173164 176032
rect 118476 175992 118482 176004
rect 173158 175992 173164 176004
rect 173216 175992 173222 176044
rect 223482 175992 223488 176044
rect 223540 176032 223546 176044
rect 232038 176032 232044 176044
rect 223540 176004 232044 176032
rect 223540 175992 223546 176004
rect 232038 175992 232044 176004
rect 232096 175992 232102 176044
rect 273990 175992 273996 176044
rect 274048 176032 274054 176044
rect 281626 176032 281632 176044
rect 274048 176004 281632 176032
rect 274048 175992 274054 176004
rect 281626 175992 281632 176004
rect 281684 175992 281690 176044
rect 115750 175924 115756 175976
rect 115808 175964 115814 175976
rect 184290 175964 184296 175976
rect 115808 175936 184296 175964
rect 115808 175924 115814 175936
rect 184290 175924 184296 175936
rect 184348 175924 184354 175976
rect 188890 175924 188896 175976
rect 188948 175964 188954 175976
rect 230934 175964 230940 175976
rect 188948 175936 230940 175964
rect 188948 175924 188954 175936
rect 230934 175924 230940 175936
rect 230992 175924 230998 175976
rect 268470 175924 268476 175976
rect 268528 175964 268534 175976
rect 281810 175964 281816 175976
rect 268528 175936 281816 175964
rect 268528 175924 268534 175936
rect 281810 175924 281816 175936
rect 281868 175924 281874 175976
rect 220906 175788 220912 175840
rect 220964 175788 220970 175840
rect 224218 175788 224224 175840
rect 224276 175788 224282 175840
rect 165430 175176 165436 175228
rect 165488 175216 165494 175228
rect 213914 175216 213920 175228
rect 165488 175188 213920 175216
rect 165488 175176 165494 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165522 175108 165528 175160
rect 165580 175148 165586 175160
rect 214006 175148 214012 175160
rect 165580 175120 214012 175148
rect 165580 175108 165586 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 220924 175148 220952 175788
rect 224236 175216 224264 175788
rect 246390 175244 246396 175296
rect 246448 175284 246454 175296
rect 264974 175284 264980 175296
rect 246448 175256 264980 175284
rect 246448 175244 246454 175256
rect 264974 175244 264980 175256
rect 265032 175244 265038 175296
rect 229278 175216 229284 175228
rect 224236 175188 229284 175216
rect 229278 175176 229284 175188
rect 229336 175176 229342 175228
rect 231118 175176 231124 175228
rect 231176 175216 231182 175228
rect 256694 175216 256700 175228
rect 231176 175188 256700 175216
rect 231176 175176 231182 175188
rect 256694 175176 256700 175188
rect 256752 175176 256758 175228
rect 229002 175148 229008 175160
rect 220924 175120 229008 175148
rect 229002 175108 229008 175120
rect 229060 175108 229066 175160
rect 231762 175108 231768 175160
rect 231820 175148 231826 175160
rect 255498 175148 255504 175160
rect 231820 175120 255504 175148
rect 231820 175108 231826 175120
rect 255498 175108 255504 175120
rect 255556 175108 255562 175160
rect 194502 175040 194508 175092
rect 194560 175080 194566 175092
rect 194560 175052 219434 175080
rect 194560 175040 194566 175052
rect 219406 175012 219434 175052
rect 230474 175012 230480 175024
rect 219406 174984 230480 175012
rect 230474 174972 230480 174984
rect 230532 174972 230538 175024
rect 209038 174496 209044 174548
rect 209096 174536 209102 174548
rect 237650 174536 237656 174548
rect 209096 174508 237656 174536
rect 209096 174496 209102 174508
rect 237650 174496 237656 174508
rect 237708 174496 237714 174548
rect 257430 174020 257436 174072
rect 257488 174060 257494 174072
rect 264974 174060 264980 174072
rect 257488 174032 264980 174060
rect 257488 174020 257494 174032
rect 264974 174020 264980 174032
rect 265032 174020 265038 174072
rect 229002 173952 229008 174004
rect 229060 173992 229066 174004
rect 229060 173952 229094 173992
rect 256142 173952 256148 174004
rect 256200 173992 256206 174004
rect 265066 173992 265072 174004
rect 256200 173964 265072 173992
rect 256200 173952 256206 173964
rect 265066 173952 265072 173964
rect 265124 173952 265130 174004
rect 229066 173924 229094 173952
rect 236270 173924 236276 173936
rect 229066 173896 236276 173924
rect 236270 173884 236276 173896
rect 236328 173884 236334 173936
rect 252094 173884 252100 173936
rect 252152 173924 252158 173936
rect 265250 173924 265256 173936
rect 252152 173896 265256 173924
rect 252152 173884 252158 173896
rect 265250 173884 265256 173896
rect 265308 173884 265314 173936
rect 165338 173816 165344 173868
rect 165396 173856 165402 173868
rect 213914 173856 213920 173868
rect 165396 173828 213920 173856
rect 165396 173816 165402 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231578 173816 231584 173868
rect 231636 173856 231642 173868
rect 247126 173856 247132 173868
rect 231636 173828 247132 173856
rect 231636 173816 231642 173828
rect 247126 173816 247132 173828
rect 247184 173816 247190 173868
rect 173250 173748 173256 173800
rect 173308 173788 173314 173800
rect 214006 173788 214012 173800
rect 173308 173760 214012 173788
rect 173308 173748 173314 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 229186 173612 229192 173664
rect 229244 173652 229250 173664
rect 229370 173652 229376 173664
rect 229244 173624 229376 173652
rect 229244 173612 229250 173624
rect 229370 173612 229376 173624
rect 229428 173612 229434 173664
rect 281718 173544 281724 173596
rect 281776 173584 281782 173596
rect 284294 173584 284300 173596
rect 281776 173556 284300 173584
rect 281776 173544 281782 173556
rect 284294 173544 284300 173556
rect 284352 173544 284358 173596
rect 229094 173204 229100 173256
rect 229152 173244 229158 173256
rect 229462 173244 229468 173256
rect 229152 173216 229468 173244
rect 229152 173204 229158 173216
rect 229462 173204 229468 173216
rect 229520 173204 229526 173256
rect 247954 173136 247960 173188
rect 248012 173176 248018 173188
rect 265158 173176 265164 173188
rect 248012 173148 265164 173176
rect 248012 173136 248018 173148
rect 265158 173136 265164 173148
rect 265216 173136 265222 173188
rect 240962 172660 240968 172712
rect 241020 172700 241026 172712
rect 264974 172700 264980 172712
rect 241020 172672 264980 172700
rect 241020 172660 241026 172672
rect 264974 172660 264980 172672
rect 265032 172660 265038 172712
rect 260374 172524 260380 172576
rect 260432 172564 260438 172576
rect 265066 172564 265072 172576
rect 260432 172536 265072 172564
rect 260432 172524 260438 172536
rect 265066 172524 265072 172536
rect 265124 172524 265130 172576
rect 168374 172456 168380 172508
rect 168432 172496 168438 172508
rect 213914 172496 213920 172508
rect 168432 172468 213920 172496
rect 168432 172456 168438 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 231670 172456 231676 172508
rect 231728 172496 231734 172508
rect 259454 172496 259460 172508
rect 231728 172468 259460 172496
rect 231728 172456 231734 172468
rect 259454 172456 259460 172468
rect 259512 172456 259518 172508
rect 184382 172388 184388 172440
rect 184440 172428 184446 172440
rect 214006 172428 214012 172440
rect 184440 172400 214012 172428
rect 184440 172388 184446 172400
rect 214006 172388 214012 172400
rect 214064 172388 214070 172440
rect 231762 172388 231768 172440
rect 231820 172428 231826 172440
rect 248414 172428 248420 172440
rect 231820 172400 248420 172428
rect 231820 172388 231826 172400
rect 248414 172388 248420 172400
rect 248472 172388 248478 172440
rect 282638 172388 282644 172440
rect 282696 172428 282702 172440
rect 285950 172428 285956 172440
rect 282696 172400 285956 172428
rect 282696 172388 282702 172400
rect 285950 172388 285956 172400
rect 286008 172388 286014 172440
rect 231486 172184 231492 172236
rect 231544 172224 231550 172236
rect 235258 172224 235264 172236
rect 231544 172196 235264 172224
rect 231544 172184 231550 172196
rect 235258 172184 235264 172196
rect 235316 172184 235322 172236
rect 262950 171504 262956 171556
rect 263008 171544 263014 171556
rect 264974 171544 264980 171556
rect 263008 171516 264980 171544
rect 263008 171504 263014 171516
rect 264974 171504 264980 171516
rect 265032 171504 265038 171556
rect 250438 171164 250444 171216
rect 250496 171204 250502 171216
rect 265066 171204 265072 171216
rect 250496 171176 265072 171204
rect 250496 171164 250502 171176
rect 265066 171164 265072 171176
rect 265124 171164 265130 171216
rect 167914 171096 167920 171148
rect 167972 171136 167978 171148
rect 184198 171136 184204 171148
rect 167972 171108 184204 171136
rect 167972 171096 167978 171108
rect 184198 171096 184204 171108
rect 184256 171096 184262 171148
rect 249150 171096 249156 171148
rect 249208 171136 249214 171148
rect 264974 171136 264980 171148
rect 249208 171108 264980 171136
rect 249208 171096 249214 171108
rect 264974 171096 264980 171108
rect 265032 171096 265038 171148
rect 167730 171028 167736 171080
rect 167788 171068 167794 171080
rect 213914 171068 213920 171080
rect 167788 171040 213920 171068
rect 167788 171028 167794 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 251174 171068 251180 171080
rect 231820 171040 251180 171068
rect 231820 171028 231826 171040
rect 251174 171028 251180 171040
rect 251232 171028 251238 171080
rect 186958 170960 186964 171012
rect 187016 171000 187022 171012
rect 214006 171000 214012 171012
rect 187016 170972 214012 171000
rect 187016 170960 187022 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 231486 170960 231492 171012
rect 231544 171000 231550 171012
rect 240226 171000 240232 171012
rect 231544 170972 240232 171000
rect 231544 170960 231550 170972
rect 240226 170960 240232 170972
rect 240284 170960 240290 171012
rect 231210 170756 231216 170808
rect 231268 170796 231274 170808
rect 236086 170796 236092 170808
rect 231268 170768 236092 170796
rect 231268 170756 231274 170768
rect 236086 170756 236092 170768
rect 236144 170756 236150 170808
rect 281718 170620 281724 170672
rect 281776 170660 281782 170672
rect 283466 170660 283472 170672
rect 281776 170632 283472 170660
rect 281776 170620 281782 170632
rect 283466 170620 283472 170632
rect 283524 170620 283530 170672
rect 258810 169872 258816 169924
rect 258868 169912 258874 169924
rect 265158 169912 265164 169924
rect 258868 169884 265164 169912
rect 258868 169872 258874 169884
rect 265158 169872 265164 169884
rect 265216 169872 265222 169924
rect 257338 169804 257344 169856
rect 257396 169844 257402 169856
rect 264974 169844 264980 169856
rect 257396 169816 264980 169844
rect 257396 169804 257402 169816
rect 264974 169804 264980 169816
rect 265032 169804 265038 169856
rect 239490 169736 239496 169788
rect 239548 169776 239554 169788
rect 265066 169776 265072 169788
rect 239548 169748 265072 169776
rect 239548 169736 239554 169748
rect 265066 169736 265072 169748
rect 265124 169736 265130 169788
rect 166442 169668 166448 169720
rect 166500 169708 166506 169720
rect 213914 169708 213920 169720
rect 166500 169680 213920 169708
rect 166500 169668 166506 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 231118 169668 231124 169720
rect 231176 169708 231182 169720
rect 233418 169708 233424 169720
rect 231176 169680 233424 169708
rect 231176 169668 231182 169680
rect 233418 169668 233424 169680
rect 233476 169668 233482 169720
rect 175918 169600 175924 169652
rect 175976 169640 175982 169652
rect 214006 169640 214012 169652
rect 175976 169612 214012 169640
rect 175976 169600 175982 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 231762 169532 231768 169584
rect 231820 169572 231826 169584
rect 238754 169572 238760 169584
rect 231820 169544 238760 169572
rect 231820 169532 231826 169544
rect 238754 169532 238760 169544
rect 238812 169532 238818 169584
rect 282730 168716 282736 168768
rect 282788 168756 282794 168768
rect 288618 168756 288624 168768
rect 282788 168728 288624 168756
rect 282788 168716 282794 168728
rect 288618 168716 288624 168728
rect 288676 168716 288682 168768
rect 282822 168648 282828 168700
rect 282880 168688 282886 168700
rect 287238 168688 287244 168700
rect 282880 168660 287244 168688
rect 282880 168648 282886 168660
rect 287238 168648 287244 168660
rect 287296 168648 287302 168700
rect 260282 168580 260288 168632
rect 260340 168620 260346 168632
rect 265250 168620 265256 168632
rect 260340 168592 265256 168620
rect 260340 168580 260346 168592
rect 265250 168580 265256 168592
rect 265308 168580 265314 168632
rect 254762 168512 254768 168564
rect 254820 168552 254826 168564
rect 265066 168552 265072 168564
rect 254820 168524 265072 168552
rect 254820 168512 254826 168524
rect 265066 168512 265072 168524
rect 265124 168512 265130 168564
rect 253474 168444 253480 168496
rect 253532 168484 253538 168496
rect 264974 168484 264980 168496
rect 253532 168456 264980 168484
rect 253532 168444 253538 168456
rect 264974 168444 264980 168456
rect 265032 168444 265038 168496
rect 244918 168376 244924 168428
rect 244976 168416 244982 168428
rect 265158 168416 265164 168428
rect 244976 168388 265164 168416
rect 244976 168376 244982 168388
rect 265158 168376 265164 168388
rect 265216 168376 265222 168428
rect 169110 168308 169116 168360
rect 169168 168348 169174 168360
rect 213914 168348 213920 168360
rect 169168 168320 213920 168348
rect 169168 168308 169174 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 251358 168348 251364 168360
rect 231820 168320 251364 168348
rect 231820 168308 231826 168320
rect 251358 168308 251364 168320
rect 251416 168308 251422 168360
rect 282730 168308 282736 168360
rect 282788 168348 282794 168360
rect 301038 168348 301044 168360
rect 282788 168320 301044 168348
rect 282788 168308 282794 168320
rect 301038 168308 301044 168320
rect 301096 168308 301102 168360
rect 177390 168240 177396 168292
rect 177448 168280 177454 168292
rect 214006 168280 214012 168292
rect 177448 168252 214012 168280
rect 177448 168240 177454 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 231394 168240 231400 168292
rect 231452 168280 231458 168292
rect 247034 168280 247040 168292
rect 231452 168252 247040 168280
rect 231452 168240 231458 168252
rect 247034 168240 247040 168252
rect 247092 168240 247098 168292
rect 282822 168240 282828 168292
rect 282880 168280 282886 168292
rect 288434 168280 288440 168292
rect 282880 168252 288440 168280
rect 282880 168240 282886 168252
rect 288434 168240 288440 168252
rect 288492 168240 288498 168292
rect 231670 168036 231676 168088
rect 231728 168076 231734 168088
rect 234798 168076 234804 168088
rect 231728 168048 234804 168076
rect 231728 168036 231734 168048
rect 234798 168036 234804 168048
rect 234856 168036 234862 168088
rect 261754 167084 261760 167136
rect 261812 167124 261818 167136
rect 265158 167124 265164 167136
rect 261812 167096 265164 167124
rect 261812 167084 261818 167096
rect 265158 167084 265164 167096
rect 265216 167084 265222 167136
rect 241146 167016 241152 167068
rect 241204 167056 241210 167068
rect 264974 167056 264980 167068
rect 241204 167028 264980 167056
rect 241204 167016 241210 167028
rect 264974 167016 264980 167028
rect 265032 167016 265038 167068
rect 173158 166948 173164 167000
rect 173216 166988 173222 167000
rect 214098 166988 214104 167000
rect 173216 166960 214104 166988
rect 173216 166948 173222 166960
rect 214098 166948 214104 166960
rect 214156 166948 214162 167000
rect 174538 166880 174544 166932
rect 174596 166920 174602 166932
rect 214006 166920 214012 166932
rect 174596 166892 214012 166920
rect 174596 166880 174602 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 200758 166812 200764 166864
rect 200816 166852 200822 166864
rect 213914 166852 213920 166864
rect 200816 166824 213920 166852
rect 200816 166812 200822 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 231026 166676 231032 166728
rect 231084 166716 231090 166728
rect 233878 166716 233884 166728
rect 231084 166688 233884 166716
rect 231084 166676 231090 166688
rect 233878 166676 233884 166688
rect 233936 166676 233942 166728
rect 231302 166540 231308 166592
rect 231360 166580 231366 166592
rect 236178 166580 236184 166592
rect 231360 166552 236184 166580
rect 231360 166540 231366 166552
rect 236178 166540 236184 166552
rect 236236 166540 236242 166592
rect 251818 166336 251824 166388
rect 251876 166376 251882 166388
rect 265066 166376 265072 166388
rect 251876 166348 265072 166376
rect 251876 166336 251882 166348
rect 265066 166336 265072 166348
rect 265124 166336 265130 166388
rect 231118 166268 231124 166320
rect 231176 166308 231182 166320
rect 252646 166308 252652 166320
rect 231176 166280 252652 166308
rect 231176 166268 231182 166280
rect 252646 166268 252652 166280
rect 252704 166268 252710 166320
rect 230474 165860 230480 165912
rect 230532 165900 230538 165912
rect 232130 165900 232136 165912
rect 230532 165872 232136 165900
rect 230532 165860 230538 165872
rect 232130 165860 232136 165872
rect 232188 165860 232194 165912
rect 253290 165656 253296 165708
rect 253348 165696 253354 165708
rect 264974 165696 264980 165708
rect 253348 165668 264980 165696
rect 253348 165656 253354 165668
rect 264974 165656 264980 165668
rect 265032 165656 265038 165708
rect 242434 165588 242440 165640
rect 242492 165628 242498 165640
rect 265066 165628 265072 165640
rect 242492 165600 265072 165628
rect 242492 165588 242498 165600
rect 265066 165588 265072 165600
rect 265124 165588 265130 165640
rect 171778 165520 171784 165572
rect 171836 165560 171842 165572
rect 214006 165560 214012 165572
rect 171836 165532 214012 165560
rect 171836 165520 171842 165532
rect 214006 165520 214012 165532
rect 214064 165520 214070 165572
rect 231394 165520 231400 165572
rect 231452 165560 231458 165572
rect 249886 165560 249892 165572
rect 231452 165532 249892 165560
rect 231452 165520 231458 165532
rect 249886 165520 249892 165532
rect 249944 165520 249950 165572
rect 281994 165520 282000 165572
rect 282052 165560 282058 165572
rect 299658 165560 299664 165572
rect 282052 165532 299664 165560
rect 282052 165520 282058 165532
rect 299658 165520 299664 165532
rect 299716 165520 299722 165572
rect 184290 165452 184296 165504
rect 184348 165492 184354 165504
rect 213914 165492 213920 165504
rect 184348 165464 213920 165492
rect 184348 165452 184354 165464
rect 213914 165452 213920 165464
rect 213972 165452 213978 165504
rect 282822 165452 282828 165504
rect 282880 165492 282886 165504
rect 296806 165492 296812 165504
rect 282880 165464 296812 165492
rect 282880 165452 282886 165464
rect 296806 165452 296812 165464
rect 296864 165452 296870 165504
rect 231302 165112 231308 165164
rect 231360 165152 231366 165164
rect 237558 165152 237564 165164
rect 231360 165124 237564 165152
rect 231360 165112 231366 165124
rect 237558 165112 237564 165124
rect 237616 165112 237622 165164
rect 250714 164840 250720 164892
rect 250772 164880 250778 164892
rect 265158 164880 265164 164892
rect 250772 164852 265164 164880
rect 250772 164840 250778 164852
rect 265158 164840 265164 164852
rect 265216 164840 265222 164892
rect 261478 164296 261484 164348
rect 261536 164336 261542 164348
rect 265066 164336 265072 164348
rect 261536 164308 265072 164336
rect 261536 164296 261542 164308
rect 265066 164296 265072 164308
rect 265124 164296 265130 164348
rect 236822 164228 236828 164280
rect 236880 164268 236886 164280
rect 264974 164268 264980 164280
rect 236880 164240 264980 164268
rect 236880 164228 236886 164240
rect 264974 164228 264980 164240
rect 265032 164228 265038 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 65518 164200 65524 164212
rect 3292 164172 65524 164200
rect 3292 164160 3298 164172
rect 65518 164160 65524 164172
rect 65576 164160 65582 164212
rect 166350 164160 166356 164212
rect 166408 164200 166414 164212
rect 213914 164200 213920 164212
rect 166408 164172 213920 164200
rect 166408 164160 166414 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 231394 164160 231400 164212
rect 231452 164200 231458 164212
rect 238846 164200 238852 164212
rect 231452 164172 238852 164200
rect 231452 164160 231458 164172
rect 238846 164160 238852 164172
rect 238904 164160 238910 164212
rect 178770 163480 178776 163532
rect 178828 163520 178834 163532
rect 214926 163520 214932 163532
rect 178828 163492 214932 163520
rect 178828 163480 178834 163492
rect 214926 163480 214932 163492
rect 214984 163480 214990 163532
rect 235534 163072 235540 163124
rect 235592 163112 235598 163124
rect 265158 163112 265164 163124
rect 235592 163084 265164 163112
rect 235592 163072 235598 163084
rect 265158 163072 265164 163084
rect 265216 163072 265222 163124
rect 246298 163004 246304 163056
rect 246356 163044 246362 163056
rect 265066 163044 265072 163056
rect 246356 163016 265072 163044
rect 246356 163004 246362 163016
rect 265066 163004 265072 163016
rect 265124 163004 265130 163056
rect 242342 162936 242348 162988
rect 242400 162976 242406 162988
rect 264974 162976 264980 162988
rect 242400 162948 264980 162976
rect 242400 162936 242406 162948
rect 264974 162936 264980 162948
rect 265032 162936 265038 162988
rect 180058 162800 180064 162852
rect 180116 162840 180122 162852
rect 214006 162840 214012 162852
rect 180116 162812 214012 162840
rect 180116 162800 180122 162812
rect 214006 162800 214012 162812
rect 214064 162800 214070 162852
rect 231394 162800 231400 162852
rect 231452 162840 231458 162852
rect 258258 162840 258264 162852
rect 231452 162812 258264 162840
rect 231452 162800 231458 162812
rect 258258 162800 258264 162812
rect 258316 162800 258322 162852
rect 282086 162800 282092 162852
rect 282144 162840 282150 162852
rect 295610 162840 295616 162852
rect 282144 162812 295616 162840
rect 282144 162800 282150 162812
rect 295610 162800 295616 162812
rect 295668 162800 295674 162852
rect 182818 162732 182824 162784
rect 182876 162772 182882 162784
rect 213914 162772 213920 162784
rect 182876 162744 213920 162772
rect 182876 162732 182882 162744
rect 213914 162732 213920 162744
rect 213972 162732 213978 162784
rect 230934 162732 230940 162784
rect 230992 162772 230998 162784
rect 241606 162772 241612 162784
rect 230992 162744 241612 162772
rect 230992 162732 230998 162744
rect 241606 162732 241612 162744
rect 241664 162732 241670 162784
rect 231394 161848 231400 161900
rect 231452 161888 231458 161900
rect 237466 161888 237472 161900
rect 231452 161860 237472 161888
rect 231452 161848 231458 161860
rect 237466 161848 237472 161860
rect 237524 161848 237530 161900
rect 247862 161508 247868 161560
rect 247920 161548 247926 161560
rect 264974 161548 264980 161560
rect 247920 161520 264980 161548
rect 247920 161508 247926 161520
rect 264974 161508 264980 161520
rect 265032 161508 265038 161560
rect 238018 161440 238024 161492
rect 238076 161480 238082 161492
rect 265158 161480 265164 161492
rect 238076 161452 265164 161480
rect 238076 161440 238082 161452
rect 265158 161440 265164 161452
rect 265216 161440 265222 161492
rect 170490 161372 170496 161424
rect 170548 161412 170554 161424
rect 214006 161412 214012 161424
rect 170548 161384 214012 161412
rect 170548 161372 170554 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 230934 161372 230940 161424
rect 230992 161412 230998 161424
rect 234430 161412 234436 161424
rect 230992 161384 234436 161412
rect 230992 161372 230998 161384
rect 234430 161372 234436 161384
rect 234488 161372 234494 161424
rect 181438 161304 181444 161356
rect 181496 161344 181502 161356
rect 213914 161344 213920 161356
rect 181496 161316 213920 161344
rect 181496 161304 181502 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 231394 161168 231400 161220
rect 231452 161208 231458 161220
rect 236270 161208 236276 161220
rect 231452 161180 236276 161208
rect 231452 161168 231458 161180
rect 236270 161168 236276 161180
rect 236328 161168 236334 161220
rect 282454 161168 282460 161220
rect 282512 161208 282518 161220
rect 287330 161208 287336 161220
rect 282512 161180 287336 161208
rect 282512 161168 282518 161180
rect 287330 161168 287336 161180
rect 287388 161168 287394 161220
rect 229830 160760 229836 160812
rect 229888 160800 229894 160812
rect 240134 160800 240140 160812
rect 229888 160772 240140 160800
rect 229888 160760 229894 160772
rect 240134 160760 240140 160772
rect 240192 160760 240198 160812
rect 234154 160692 234160 160744
rect 234212 160732 234218 160744
rect 264974 160732 264980 160744
rect 234212 160704 264980 160732
rect 234212 160692 234218 160704
rect 264974 160692 264980 160704
rect 265032 160692 265038 160744
rect 260098 160216 260104 160268
rect 260156 160256 260162 160268
rect 265158 160256 265164 160268
rect 260156 160228 265164 160256
rect 260156 160216 260162 160228
rect 265158 160216 265164 160228
rect 265216 160216 265222 160268
rect 243722 160148 243728 160200
rect 243780 160188 243786 160200
rect 265066 160188 265072 160200
rect 243780 160160 265072 160188
rect 243780 160148 243786 160160
rect 265066 160148 265072 160160
rect 265124 160148 265130 160200
rect 240870 160080 240876 160132
rect 240928 160120 240934 160132
rect 264974 160120 264980 160132
rect 240928 160092 264980 160120
rect 240928 160080 240934 160092
rect 264974 160080 264980 160092
rect 265032 160080 265038 160132
rect 170398 160012 170404 160064
rect 170456 160052 170462 160064
rect 214006 160052 214012 160064
rect 170456 160024 214012 160052
rect 170456 160012 170462 160024
rect 214006 160012 214012 160024
rect 214064 160012 214070 160064
rect 231394 160012 231400 160064
rect 231452 160052 231458 160064
rect 255406 160052 255412 160064
rect 231452 160024 255412 160052
rect 231452 160012 231458 160024
rect 255406 160012 255412 160024
rect 255464 160012 255470 160064
rect 282086 160012 282092 160064
rect 282144 160052 282150 160064
rect 292850 160052 292856 160064
rect 282144 160024 292856 160052
rect 282144 160012 282150 160024
rect 292850 160012 292856 160024
rect 292908 160012 292914 160064
rect 191098 159944 191104 159996
rect 191156 159984 191162 159996
rect 213914 159984 213920 159996
rect 191156 159956 213920 159984
rect 191156 159944 191162 159956
rect 213914 159944 213920 159956
rect 213972 159944 213978 159996
rect 230934 159944 230940 159996
rect 230992 159984 230998 159996
rect 254026 159984 254032 159996
rect 230992 159956 254032 159984
rect 230992 159944 230998 159956
rect 254026 159944 254032 159956
rect 254084 159944 254090 159996
rect 258718 158856 258724 158908
rect 258776 158896 258782 158908
rect 265158 158896 265164 158908
rect 258776 158868 265164 158896
rect 258776 158856 258782 158868
rect 265158 158856 265164 158868
rect 265216 158856 265222 158908
rect 257614 158788 257620 158840
rect 257672 158828 257678 158840
rect 265066 158828 265072 158840
rect 257672 158800 265072 158828
rect 257672 158788 257678 158800
rect 265066 158788 265072 158800
rect 265124 158788 265130 158840
rect 236730 158720 236736 158772
rect 236788 158760 236794 158772
rect 264974 158760 264980 158772
rect 236788 158732 264980 158760
rect 236788 158720 236794 158732
rect 264974 158720 264980 158732
rect 265032 158720 265038 158772
rect 167638 158652 167644 158704
rect 167696 158692 167702 158704
rect 213914 158692 213920 158704
rect 167696 158664 213920 158692
rect 167696 158652 167702 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 282822 158652 282828 158704
rect 282880 158692 282886 158704
rect 294046 158692 294052 158704
rect 282880 158664 294052 158692
rect 282880 158652 282886 158664
rect 294046 158652 294052 158664
rect 294104 158652 294110 158704
rect 169018 158584 169024 158636
rect 169076 158624 169082 158636
rect 214006 158624 214012 158636
rect 169076 158596 214012 158624
rect 169076 158584 169082 158596
rect 214006 158584 214012 158596
rect 214064 158584 214070 158636
rect 231210 157972 231216 158024
rect 231268 158012 231274 158024
rect 240962 158012 240968 158024
rect 231268 157984 240968 158012
rect 231268 157972 231274 157984
rect 240962 157972 240968 157984
rect 241020 157972 241026 158024
rect 258902 157496 258908 157548
rect 258960 157536 258966 157548
rect 265158 157536 265164 157548
rect 258960 157508 265164 157536
rect 258960 157496 258966 157508
rect 265158 157496 265164 157508
rect 265216 157496 265222 157548
rect 254854 157428 254860 157480
rect 254912 157468 254918 157480
rect 265066 157468 265072 157480
rect 254912 157440 265072 157468
rect 254912 157428 254918 157440
rect 265066 157428 265072 157440
rect 265124 157428 265130 157480
rect 238294 157360 238300 157412
rect 238352 157400 238358 157412
rect 264974 157400 264980 157412
rect 238352 157372 264980 157400
rect 238352 157360 238358 157372
rect 264974 157360 264980 157372
rect 265032 157360 265038 157412
rect 203518 157292 203524 157344
rect 203576 157332 203582 157344
rect 213914 157332 213920 157344
rect 203576 157304 213920 157332
rect 203576 157292 203582 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 255314 157332 255320 157344
rect 231820 157304 255320 157332
rect 231820 157292 231826 157304
rect 255314 157292 255320 157304
rect 255372 157292 255378 157344
rect 231118 157224 231124 157276
rect 231176 157264 231182 157276
rect 244366 157264 244372 157276
rect 231176 157236 244372 157264
rect 231176 157224 231182 157236
rect 244366 157224 244372 157236
rect 244424 157224 244430 157276
rect 255958 156068 255964 156120
rect 256016 156108 256022 156120
rect 265066 156108 265072 156120
rect 256016 156080 265072 156108
rect 256016 156068 256022 156080
rect 265066 156068 265072 156080
rect 265124 156068 265130 156120
rect 241238 156000 241244 156052
rect 241296 156040 241302 156052
rect 264974 156040 264980 156052
rect 241296 156012 264980 156040
rect 241296 156000 241302 156012
rect 264974 156000 264980 156012
rect 265032 156000 265038 156052
rect 234062 155932 234068 155984
rect 234120 155972 234126 155984
rect 265158 155972 265164 155984
rect 234120 155944 265164 155972
rect 234120 155932 234126 155944
rect 265158 155932 265164 155944
rect 265216 155932 265222 155984
rect 166258 155864 166264 155916
rect 166316 155904 166322 155916
rect 213914 155904 213920 155916
rect 166316 155876 213920 155904
rect 166316 155864 166322 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 230934 155864 230940 155916
rect 230992 155904 230998 155916
rect 234706 155904 234712 155916
rect 230992 155876 234712 155904
rect 230992 155864 230998 155876
rect 234706 155864 234712 155876
rect 234764 155864 234770 155916
rect 177298 155796 177304 155848
rect 177356 155836 177362 155848
rect 214006 155836 214012 155848
rect 177356 155808 214012 155836
rect 177356 155796 177362 155808
rect 214006 155796 214012 155808
rect 214064 155796 214070 155848
rect 232498 155184 232504 155236
rect 232556 155224 232562 155236
rect 265618 155224 265624 155236
rect 232556 155196 265624 155224
rect 232556 155184 232562 155196
rect 265618 155184 265624 155196
rect 265676 155184 265682 155236
rect 249334 154640 249340 154692
rect 249392 154680 249398 154692
rect 265066 154680 265072 154692
rect 249392 154652 265072 154680
rect 249392 154640 249398 154652
rect 265066 154640 265072 154652
rect 265124 154640 265130 154692
rect 239674 154572 239680 154624
rect 239732 154612 239738 154624
rect 264974 154612 264980 154624
rect 239732 154584 264980 154612
rect 239732 154572 239738 154584
rect 264974 154572 264980 154584
rect 265032 154572 265038 154624
rect 231762 154504 231768 154556
rect 231820 154544 231826 154556
rect 242986 154544 242992 154556
rect 231820 154516 242992 154544
rect 231820 154504 231826 154516
rect 242986 154504 242992 154516
rect 243044 154504 243050 154556
rect 281718 154504 281724 154556
rect 281776 154544 281782 154556
rect 307846 154544 307852 154556
rect 281776 154516 307852 154544
rect 281776 154504 281782 154516
rect 307846 154504 307852 154516
rect 307904 154504 307910 154556
rect 231486 153960 231492 154012
rect 231544 154000 231550 154012
rect 237650 154000 237656 154012
rect 231544 153972 237656 154000
rect 231544 153960 231550 153972
rect 237650 153960 237656 153972
rect 237708 153960 237714 154012
rect 253382 153824 253388 153876
rect 253440 153864 253446 153876
rect 265158 153864 265164 153876
rect 253440 153836 265164 153864
rect 253440 153824 253446 153836
rect 265158 153824 265164 153836
rect 265216 153824 265222 153876
rect 180058 153280 180064 153332
rect 180116 153320 180122 153332
rect 214006 153320 214012 153332
rect 180116 153292 214012 153320
rect 180116 153280 180122 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 252002 153280 252008 153332
rect 252060 153320 252066 153332
rect 265066 153320 265072 153332
rect 252060 153292 265072 153320
rect 252060 153280 252066 153292
rect 265066 153280 265072 153292
rect 265124 153280 265130 153332
rect 166258 153212 166264 153264
rect 166316 153252 166322 153264
rect 213914 153252 213920 153264
rect 166316 153224 213920 153252
rect 166316 153212 166322 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 232774 153212 232780 153264
rect 232832 153252 232838 153264
rect 264974 153252 264980 153264
rect 232832 153224 264980 153252
rect 232832 153212 232838 153224
rect 264974 153212 264980 153224
rect 265032 153212 265038 153264
rect 231394 153144 231400 153196
rect 231452 153184 231458 153196
rect 251266 153184 251272 153196
rect 231452 153156 251272 153184
rect 231452 153144 231458 153156
rect 251266 153144 251272 153156
rect 251324 153144 251330 153196
rect 231762 153076 231768 153128
rect 231820 153116 231826 153128
rect 245746 153116 245752 153128
rect 231820 153088 245752 153116
rect 231820 153076 231826 153088
rect 245746 153076 245752 153088
rect 245804 153076 245810 153128
rect 229738 152532 229744 152584
rect 229796 152572 229802 152584
rect 248506 152572 248512 152584
rect 229796 152544 248512 152572
rect 229796 152532 229802 152544
rect 248506 152532 248512 152544
rect 248564 152532 248570 152584
rect 229922 152464 229928 152516
rect 229980 152504 229986 152516
rect 265342 152504 265348 152516
rect 229980 152476 265348 152504
rect 229980 152464 229986 152476
rect 265342 152464 265348 152476
rect 265400 152464 265406 152516
rect 184290 151852 184296 151904
rect 184348 151892 184354 151904
rect 213914 151892 213920 151904
rect 184348 151864 213920 151892
rect 184348 151852 184354 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 251910 151852 251916 151904
rect 251968 151892 251974 151904
rect 265066 151892 265072 151904
rect 251968 151864 265072 151892
rect 251968 151852 251974 151864
rect 265066 151852 265072 151864
rect 265124 151852 265130 151904
rect 170398 151784 170404 151836
rect 170456 151824 170462 151836
rect 214006 151824 214012 151836
rect 170456 151796 214012 151824
rect 170456 151784 170462 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 245102 151784 245108 151836
rect 245160 151824 245166 151836
rect 264974 151824 264980 151836
rect 245160 151796 264980 151824
rect 245160 151784 245166 151796
rect 264974 151784 264980 151796
rect 265032 151784 265038 151836
rect 282822 151716 282828 151768
rect 282880 151756 282886 151768
rect 302510 151756 302516 151768
rect 282880 151728 302516 151756
rect 282880 151716 282886 151728
rect 302510 151716 302516 151728
rect 302568 151716 302574 151768
rect 231210 151580 231216 151632
rect 231268 151620 231274 151632
rect 233326 151620 233332 151632
rect 231268 151592 233332 151620
rect 231268 151580 231274 151592
rect 233326 151580 233332 151592
rect 233384 151580 233390 151632
rect 282638 151240 282644 151292
rect 282696 151280 282702 151292
rect 285858 151280 285864 151292
rect 282696 151252 285864 151280
rect 282696 151240 282702 151252
rect 285858 151240 285864 151252
rect 285916 151240 285922 151292
rect 250622 151104 250628 151156
rect 250680 151144 250686 151156
rect 265158 151144 265164 151156
rect 250680 151116 265164 151144
rect 250680 151104 250686 151116
rect 265158 151104 265164 151116
rect 265216 151104 265222 151156
rect 200758 151036 200764 151088
rect 200816 151076 200822 151088
rect 214466 151076 214472 151088
rect 200816 151048 214472 151076
rect 200816 151036 200822 151048
rect 214466 151036 214472 151048
rect 214524 151036 214530 151088
rect 231210 151036 231216 151088
rect 231268 151076 231274 151088
rect 252094 151076 252100 151088
rect 231268 151048 252100 151076
rect 231268 151036 231274 151048
rect 252094 151036 252100 151048
rect 252152 151036 252158 151088
rect 197998 150424 198004 150476
rect 198056 150464 198062 150476
rect 213914 150464 213920 150476
rect 198056 150436 213920 150464
rect 198056 150424 198062 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 249058 150424 249064 150476
rect 249116 150464 249122 150476
rect 264974 150464 264980 150476
rect 249116 150436 264980 150464
rect 249116 150424 249122 150436
rect 264974 150424 264980 150436
rect 265032 150424 265038 150476
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 43438 150396 43444 150408
rect 3568 150368 43444 150396
rect 3568 150356 3574 150368
rect 43438 150356 43444 150368
rect 43496 150356 43502 150408
rect 184198 150356 184204 150408
rect 184256 150396 184262 150408
rect 214006 150396 214012 150408
rect 184256 150368 214012 150396
rect 184256 150356 184262 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 230934 150356 230940 150408
rect 230992 150396 230998 150408
rect 253934 150396 253940 150408
rect 230992 150368 253940 150396
rect 230992 150356 230998 150368
rect 253934 150356 253940 150368
rect 253992 150356 253998 150408
rect 282822 150356 282828 150408
rect 282880 150396 282886 150408
rect 290090 150396 290096 150408
rect 282880 150368 290096 150396
rect 282880 150356 282886 150368
rect 290090 150356 290096 150368
rect 290148 150356 290154 150408
rect 198090 150288 198096 150340
rect 198148 150328 198154 150340
rect 213914 150328 213920 150340
rect 198148 150300 213920 150328
rect 198148 150288 198154 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 230842 150288 230848 150340
rect 230900 150328 230906 150340
rect 240778 150328 240784 150340
rect 230900 150300 240784 150328
rect 230900 150288 230906 150300
rect 240778 150288 240784 150300
rect 240836 150288 240842 150340
rect 234246 149744 234252 149796
rect 234304 149784 234310 149796
rect 249794 149784 249800 149796
rect 234304 149756 249800 149784
rect 234304 149744 234310 149756
rect 249794 149744 249800 149756
rect 249852 149744 249858 149796
rect 246574 149676 246580 149728
rect 246632 149716 246638 149728
rect 265250 149716 265256 149728
rect 246632 149688 265256 149716
rect 246632 149676 246638 149688
rect 265250 149676 265256 149688
rect 265308 149676 265314 149728
rect 281718 149608 281724 149660
rect 281776 149648 281782 149660
rect 284570 149648 284576 149660
rect 281776 149620 284576 149648
rect 281776 149608 281782 149620
rect 284570 149608 284576 149620
rect 284628 149608 284634 149660
rect 263042 149200 263048 149252
rect 263100 149240 263106 149252
rect 265434 149240 265440 149252
rect 263100 149212 265440 149240
rect 263100 149200 263106 149212
rect 265434 149200 265440 149212
rect 265492 149200 265498 149252
rect 253198 149132 253204 149184
rect 253256 149172 253262 149184
rect 264974 149172 264980 149184
rect 253256 149144 264980 149172
rect 253256 149132 253262 149144
rect 264974 149132 264980 149144
rect 265032 149132 265038 149184
rect 235442 149064 235448 149116
rect 235500 149104 235506 149116
rect 265066 149104 265072 149116
rect 235500 149076 265072 149104
rect 235500 149064 235506 149076
rect 265066 149064 265072 149076
rect 265124 149064 265130 149116
rect 207658 148996 207664 149048
rect 207716 149036 207722 149048
rect 213914 149036 213920 149048
rect 207716 149008 213920 149036
rect 207716 148996 207722 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 244458 149036 244464 149048
rect 231820 149008 244464 149036
rect 231820 148996 231826 149008
rect 244458 148996 244464 149008
rect 244516 148996 244522 149048
rect 282730 148996 282736 149048
rect 282788 149036 282794 149048
rect 292758 149036 292764 149048
rect 282788 149008 292764 149036
rect 282788 148996 282794 149008
rect 292758 148996 292764 149008
rect 292816 148996 292822 149048
rect 282822 148928 282828 148980
rect 282880 148968 282886 148980
rect 287054 148968 287060 148980
rect 282880 148940 287060 148968
rect 282880 148928 282886 148940
rect 287054 148928 287060 148940
rect 287112 148928 287118 148980
rect 231118 148316 231124 148368
rect 231176 148356 231182 148368
rect 234614 148356 234620 148368
rect 231176 148328 234620 148356
rect 231176 148316 231182 148328
rect 234614 148316 234620 148328
rect 234672 148316 234678 148368
rect 257430 148356 257436 148368
rect 238726 148328 257436 148356
rect 231394 148248 231400 148300
rect 231452 148288 231458 148300
rect 238726 148288 238754 148328
rect 257430 148316 257436 148328
rect 257488 148316 257494 148368
rect 231452 148260 238754 148288
rect 231452 148248 231458 148260
rect 262858 147840 262864 147892
rect 262916 147880 262922 147892
rect 265342 147880 265348 147892
rect 262916 147852 265348 147880
rect 262916 147840 262922 147852
rect 265342 147840 265348 147852
rect 265400 147840 265406 147892
rect 260466 147772 260472 147824
rect 260524 147812 260530 147824
rect 265066 147812 265072 147824
rect 260524 147784 265072 147812
rect 260524 147772 260530 147784
rect 265066 147772 265072 147784
rect 265124 147772 265130 147824
rect 264422 147704 264428 147756
rect 264480 147744 264486 147756
rect 266078 147744 266084 147756
rect 264480 147716 266084 147744
rect 264480 147704 264486 147716
rect 266078 147704 266084 147716
rect 266136 147704 266142 147756
rect 166350 147636 166356 147688
rect 166408 147676 166414 147688
rect 213914 147676 213920 147688
rect 166408 147648 213920 147676
rect 166408 147636 166414 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 250530 147636 250536 147688
rect 250588 147676 250594 147688
rect 264974 147676 264980 147688
rect 250588 147648 264980 147676
rect 250588 147636 250594 147648
rect 264974 147636 264980 147648
rect 265032 147636 265038 147688
rect 256050 146888 256056 146940
rect 256108 146928 256114 146940
rect 265158 146928 265164 146940
rect 256108 146900 265164 146928
rect 256108 146888 256114 146900
rect 265158 146888 265164 146900
rect 265216 146888 265222 146940
rect 202138 146344 202144 146396
rect 202196 146384 202202 146396
rect 214006 146384 214012 146396
rect 202196 146356 214012 146384
rect 202196 146344 202202 146356
rect 214006 146344 214012 146356
rect 214064 146344 214070 146396
rect 245194 146344 245200 146396
rect 245252 146384 245258 146396
rect 265066 146384 265072 146396
rect 245252 146356 265072 146384
rect 245252 146344 245258 146356
rect 265066 146344 265072 146356
rect 265124 146344 265130 146396
rect 195238 146276 195244 146328
rect 195296 146316 195302 146328
rect 213914 146316 213920 146328
rect 195296 146288 213920 146316
rect 195296 146276 195302 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 232590 146276 232596 146328
rect 232648 146316 232654 146328
rect 264974 146316 264980 146328
rect 232648 146288 264980 146316
rect 232648 146276 232654 146288
rect 264974 146276 264980 146288
rect 265032 146276 265038 146328
rect 231762 146208 231768 146260
rect 231820 146248 231826 146260
rect 247218 146248 247224 146260
rect 231820 146220 247224 146248
rect 231820 146208 231826 146220
rect 247218 146208 247224 146220
rect 247276 146208 247282 146260
rect 281994 146208 282000 146260
rect 282052 146248 282058 146260
rect 302418 146248 302424 146260
rect 282052 146220 302424 146248
rect 282052 146208 282058 146220
rect 302418 146208 302424 146220
rect 302476 146208 302482 146260
rect 282822 146140 282828 146192
rect 282880 146180 282886 146192
rect 291194 146180 291200 146192
rect 282880 146152 291200 146180
rect 282880 146140 282886 146152
rect 291194 146140 291200 146152
rect 291252 146140 291258 146192
rect 231670 145392 231676 145444
rect 231728 145432 231734 145444
rect 235994 145432 236000 145444
rect 231728 145404 236000 145432
rect 231728 145392 231734 145404
rect 235994 145392 236000 145404
rect 236052 145392 236058 145444
rect 247770 145052 247776 145104
rect 247828 145092 247834 145104
rect 265066 145092 265072 145104
rect 247828 145064 265072 145092
rect 247828 145052 247834 145064
rect 265066 145052 265072 145064
rect 265124 145052 265130 145104
rect 191098 144984 191104 145036
rect 191156 145024 191162 145036
rect 213914 145024 213920 145036
rect 191156 144996 213920 145024
rect 191156 144984 191162 144996
rect 213914 144984 213920 144996
rect 213972 144984 213978 145036
rect 242158 144984 242164 145036
rect 242216 145024 242222 145036
rect 264974 145024 264980 145036
rect 242216 144996 264980 145024
rect 242216 144984 242222 144996
rect 264974 144984 264980 144996
rect 265032 144984 265038 145036
rect 184198 144916 184204 144968
rect 184256 144956 184262 144968
rect 214006 144956 214012 144968
rect 184256 144928 214012 144956
rect 184256 144916 184262 144928
rect 214006 144916 214012 144928
rect 214064 144916 214070 144968
rect 235350 144916 235356 144968
rect 235408 144956 235414 144968
rect 265158 144956 265164 144968
rect 235408 144928 265164 144956
rect 235408 144916 235414 144928
rect 265158 144916 265164 144928
rect 265216 144916 265222 144968
rect 231302 144848 231308 144900
rect 231360 144888 231366 144900
rect 244274 144888 244280 144900
rect 231360 144860 244280 144888
rect 231360 144848 231366 144860
rect 244274 144848 244280 144860
rect 244332 144848 244338 144900
rect 282822 144848 282828 144900
rect 282880 144888 282886 144900
rect 294230 144888 294236 144900
rect 282880 144860 294236 144888
rect 282880 144848 282886 144860
rect 294230 144848 294236 144860
rect 294288 144848 294294 144900
rect 231486 144780 231492 144832
rect 231544 144820 231550 144832
rect 239398 144820 239404 144832
rect 231544 144792 239404 144820
rect 231544 144780 231550 144792
rect 239398 144780 239404 144792
rect 239456 144780 239462 144832
rect 237374 144168 237380 144220
rect 237432 144208 237438 144220
rect 241790 144208 241796 144220
rect 237432 144180 241796 144208
rect 237432 144168 237438 144180
rect 241790 144168 241796 144180
rect 241848 144168 241854 144220
rect 249242 144168 249248 144220
rect 249300 144208 249306 144220
rect 265250 144208 265256 144220
rect 249300 144180 265256 144208
rect 249300 144168 249306 144180
rect 265250 144168 265256 144180
rect 265308 144168 265314 144220
rect 198090 143624 198096 143676
rect 198148 143664 198154 143676
rect 214006 143664 214012 143676
rect 198148 143636 214012 143664
rect 198148 143624 198154 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 242250 143624 242256 143676
rect 242308 143664 242314 143676
rect 265066 143664 265072 143676
rect 242308 143636 265072 143664
rect 242308 143624 242314 143636
rect 265066 143624 265072 143636
rect 265124 143624 265130 143676
rect 188338 143556 188344 143608
rect 188396 143596 188402 143608
rect 213914 143596 213920 143608
rect 188396 143568 213920 143596
rect 188396 143556 188402 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 239582 143556 239588 143608
rect 239640 143596 239646 143608
rect 264974 143596 264980 143608
rect 239640 143568 264980 143596
rect 239640 143556 239646 143568
rect 264974 143556 264980 143568
rect 265032 143556 265038 143608
rect 281626 143488 281632 143540
rect 281684 143528 281690 143540
rect 296990 143528 296996 143540
rect 281684 143500 296996 143528
rect 281684 143488 281690 143500
rect 296990 143488 296996 143500
rect 297048 143488 297054 143540
rect 231302 143352 231308 143404
rect 231360 143392 231366 143404
rect 237374 143392 237380 143404
rect 231360 143364 237380 143392
rect 231360 143352 231366 143364
rect 237374 143352 237380 143364
rect 237432 143352 237438 143404
rect 256234 142264 256240 142316
rect 256292 142304 256298 142316
rect 264974 142304 264980 142316
rect 256292 142276 264980 142304
rect 256292 142264 256298 142276
rect 264974 142264 264980 142276
rect 265032 142264 265038 142316
rect 241054 142196 241060 142248
rect 241112 142236 241118 142248
rect 265158 142236 265164 142248
rect 241112 142208 265164 142236
rect 241112 142196 241118 142208
rect 265158 142196 265164 142208
rect 265216 142196 265222 142248
rect 186958 142128 186964 142180
rect 187016 142168 187022 142180
rect 213914 142168 213920 142180
rect 187016 142140 213920 142168
rect 187016 142128 187022 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 238202 142128 238208 142180
rect 238260 142168 238266 142180
rect 265066 142168 265072 142180
rect 238260 142140 265072 142168
rect 238260 142128 238266 142140
rect 265066 142128 265072 142140
rect 265124 142128 265130 142180
rect 231762 142060 231768 142112
rect 231820 142100 231826 142112
rect 258166 142100 258172 142112
rect 231820 142072 258172 142100
rect 231820 142060 231826 142072
rect 258166 142060 258172 142072
rect 258224 142060 258230 142112
rect 282730 142060 282736 142112
rect 282788 142100 282794 142112
rect 299750 142100 299756 142112
rect 282788 142072 299756 142100
rect 282788 142060 282794 142072
rect 299750 142060 299756 142072
rect 299808 142060 299814 142112
rect 282822 141992 282828 142044
rect 282880 142032 282886 142044
rect 298370 142032 298376 142044
rect 282880 142004 298376 142032
rect 282880 141992 282886 142004
rect 298370 141992 298376 142004
rect 298428 141992 298434 142044
rect 282822 141380 282828 141432
rect 282880 141420 282886 141432
rect 291470 141420 291476 141432
rect 282880 141392 291476 141420
rect 282880 141380 282886 141392
rect 291470 141380 291476 141392
rect 291528 141380 291534 141432
rect 252094 140904 252100 140956
rect 252152 140944 252158 140956
rect 264974 140944 264980 140956
rect 252152 140916 264980 140944
rect 252152 140904 252158 140916
rect 264974 140904 264980 140916
rect 265032 140904 265038 140956
rect 189718 140836 189724 140888
rect 189776 140876 189782 140888
rect 213914 140876 213920 140888
rect 189776 140848 213920 140876
rect 189776 140836 189782 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 240962 140836 240968 140888
rect 241020 140876 241026 140888
rect 265066 140876 265072 140888
rect 241020 140848 265072 140876
rect 241020 140836 241026 140848
rect 265066 140836 265072 140848
rect 265124 140836 265130 140888
rect 177390 140768 177396 140820
rect 177448 140808 177454 140820
rect 214006 140808 214012 140820
rect 177448 140780 214012 140808
rect 177448 140768 177454 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 233878 140768 233884 140820
rect 233936 140808 233942 140820
rect 265158 140808 265164 140820
rect 233936 140780 265164 140808
rect 233936 140768 233942 140780
rect 265158 140768 265164 140780
rect 265216 140768 265222 140820
rect 231670 140700 231676 140752
rect 231728 140740 231734 140752
rect 260834 140740 260840 140752
rect 231728 140712 260840 140740
rect 231728 140700 231734 140712
rect 260834 140700 260840 140712
rect 260892 140700 260898 140752
rect 281902 140700 281908 140752
rect 281960 140740 281966 140752
rect 289998 140740 290004 140752
rect 281960 140712 290004 140740
rect 281960 140700 281966 140712
rect 289998 140700 290004 140712
rect 290056 140700 290062 140752
rect 231762 140632 231768 140684
rect 231820 140672 231826 140684
rect 242894 140672 242900 140684
rect 231820 140644 242900 140672
rect 231820 140632 231826 140644
rect 242894 140632 242900 140644
rect 242952 140632 242958 140684
rect 206370 139476 206376 139528
rect 206428 139516 206434 139528
rect 214006 139516 214012 139528
rect 206428 139488 214012 139516
rect 206428 139476 206434 139488
rect 214006 139476 214012 139488
rect 214064 139476 214070 139528
rect 187142 139408 187148 139460
rect 187200 139448 187206 139460
rect 213914 139448 213920 139460
rect 187200 139420 213920 139448
rect 187200 139408 187206 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 243538 139408 243544 139460
rect 243596 139448 243602 139460
rect 264974 139448 264980 139460
rect 243596 139420 264980 139448
rect 243596 139408 243602 139420
rect 264974 139408 264980 139420
rect 265032 139408 265038 139460
rect 231762 139340 231768 139392
rect 231820 139380 231826 139392
rect 245654 139380 245660 139392
rect 231820 139352 245660 139380
rect 231820 139340 231826 139352
rect 245654 139340 245660 139352
rect 245712 139340 245718 139392
rect 583386 139340 583392 139392
rect 583444 139380 583450 139392
rect 583846 139380 583852 139392
rect 583444 139352 583852 139380
rect 583444 139340 583450 139352
rect 583846 139340 583852 139352
rect 583904 139340 583910 139392
rect 177298 138660 177304 138712
rect 177356 138700 177362 138712
rect 214926 138700 214932 138712
rect 177356 138672 214932 138700
rect 177356 138660 177362 138672
rect 214926 138660 214932 138672
rect 214984 138660 214990 138712
rect 231302 138660 231308 138712
rect 231360 138700 231366 138712
rect 239490 138700 239496 138712
rect 231360 138672 239496 138700
rect 231360 138660 231366 138672
rect 239490 138660 239496 138672
rect 239548 138660 239554 138712
rect 254670 138048 254676 138100
rect 254728 138088 254734 138100
rect 265066 138088 265072 138100
rect 254728 138060 265072 138088
rect 254728 138048 254734 138060
rect 265066 138048 265072 138060
rect 265124 138048 265130 138100
rect 185578 137980 185584 138032
rect 185636 138020 185642 138032
rect 214006 138020 214012 138032
rect 185636 137992 214012 138020
rect 185636 137980 185642 137992
rect 214006 137980 214012 137992
rect 214064 137980 214070 138032
rect 239398 137980 239404 138032
rect 239456 138020 239462 138032
rect 264974 138020 264980 138032
rect 239456 137992 264980 138020
rect 239456 137980 239462 137992
rect 264974 137980 264980 137992
rect 265032 137980 265038 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 32398 137952 32404 137964
rect 3568 137924 32404 137952
rect 3568 137912 3574 137924
rect 32398 137912 32404 137924
rect 32456 137912 32462 137964
rect 282822 137912 282828 137964
rect 282880 137952 282886 137964
rect 306466 137952 306472 137964
rect 282880 137924 306472 137952
rect 282880 137912 282886 137924
rect 306466 137912 306472 137924
rect 306524 137912 306530 137964
rect 231670 137844 231676 137896
rect 231728 137884 231734 137896
rect 234246 137884 234252 137896
rect 231728 137856 234252 137884
rect 231728 137844 231734 137856
rect 234246 137844 234252 137856
rect 234304 137844 234310 137896
rect 240778 136756 240784 136808
rect 240836 136796 240842 136808
rect 265066 136796 265072 136808
rect 240836 136768 265072 136796
rect 240836 136756 240842 136768
rect 265066 136756 265072 136768
rect 265124 136756 265130 136808
rect 236638 136688 236644 136740
rect 236696 136728 236702 136740
rect 264974 136728 264980 136740
rect 236696 136700 264980 136728
rect 236696 136688 236702 136700
rect 264974 136688 264980 136700
rect 265032 136688 265038 136740
rect 169018 136620 169024 136672
rect 169076 136660 169082 136672
rect 213914 136660 213920 136672
rect 169076 136632 213920 136660
rect 169076 136620 169082 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 233970 136620 233976 136672
rect 234028 136660 234034 136672
rect 265250 136660 265256 136672
rect 234028 136632 265256 136660
rect 234028 136620 234034 136632
rect 265250 136620 265256 136632
rect 265308 136620 265314 136672
rect 282362 136552 282368 136604
rect 282420 136592 282426 136604
rect 304994 136592 305000 136604
rect 282420 136564 305000 136592
rect 282420 136552 282426 136564
rect 304994 136552 305000 136564
rect 305052 136552 305058 136604
rect 282546 136348 282552 136400
rect 282604 136388 282610 136400
rect 285766 136388 285772 136400
rect 282604 136360 285772 136388
rect 282604 136348 282610 136360
rect 285766 136348 285772 136360
rect 285824 136348 285830 136400
rect 182818 135872 182824 135924
rect 182876 135912 182882 135924
rect 214098 135912 214104 135924
rect 182876 135884 214104 135912
rect 182876 135872 182882 135884
rect 214098 135872 214104 135884
rect 214156 135872 214162 135924
rect 231118 135872 231124 135924
rect 231176 135912 231182 135924
rect 264514 135912 264520 135924
rect 231176 135884 264520 135912
rect 231176 135872 231182 135884
rect 264514 135872 264520 135884
rect 264572 135872 264578 135924
rect 229738 135464 229744 135516
rect 229796 135504 229802 135516
rect 265066 135504 265072 135516
rect 229796 135476 265072 135504
rect 229796 135464 229802 135476
rect 265066 135464 265072 135476
rect 265124 135464 265130 135516
rect 257430 135396 257436 135448
rect 257488 135436 257494 135448
rect 265158 135436 265164 135448
rect 257488 135408 265164 135436
rect 257488 135396 257494 135408
rect 265158 135396 265164 135408
rect 265216 135396 265222 135448
rect 209130 135328 209136 135380
rect 209188 135368 209194 135380
rect 214006 135368 214012 135380
rect 209188 135340 214012 135368
rect 209188 135328 209194 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 245010 135328 245016 135380
rect 245068 135368 245074 135380
rect 264974 135368 264980 135380
rect 245068 135340 264980 135368
rect 245068 135328 245074 135340
rect 264974 135328 264980 135340
rect 265032 135328 265038 135380
rect 181438 135260 181444 135312
rect 181496 135300 181502 135312
rect 213914 135300 213920 135312
rect 181496 135272 213920 135300
rect 181496 135260 181502 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 231762 135192 231768 135244
rect 231820 135232 231826 135244
rect 256142 135232 256148 135244
rect 231820 135204 256148 135232
rect 231820 135192 231826 135204
rect 256142 135192 256148 135204
rect 256200 135192 256206 135244
rect 231670 135124 231676 135176
rect 231728 135164 231734 135176
rect 247954 135164 247960 135176
rect 231728 135136 247960 135164
rect 231728 135124 231734 135136
rect 247954 135124 247960 135136
rect 248012 135124 248018 135176
rect 247678 134036 247684 134088
rect 247736 134076 247742 134088
rect 265066 134076 265072 134088
rect 247736 134048 265072 134076
rect 247736 134036 247742 134048
rect 265066 134036 265072 134048
rect 265124 134036 265130 134088
rect 239490 133968 239496 134020
rect 239548 134008 239554 134020
rect 264974 134008 264980 134020
rect 239548 133980 264980 134008
rect 239548 133968 239554 133980
rect 264974 133968 264980 133980
rect 265032 133968 265038 134020
rect 173342 133900 173348 133952
rect 173400 133940 173406 133952
rect 213914 133940 213920 133952
rect 173400 133912 213920 133940
rect 173400 133900 173406 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 238110 133900 238116 133952
rect 238168 133940 238174 133952
rect 265158 133940 265164 133952
rect 238168 133912 265164 133940
rect 238168 133900 238174 133912
rect 265158 133900 265164 133912
rect 265216 133900 265222 133952
rect 231670 133832 231676 133884
rect 231728 133872 231734 133884
rect 262950 133872 262956 133884
rect 231728 133844 262956 133872
rect 231728 133832 231734 133844
rect 262950 133832 262956 133844
rect 263008 133832 263014 133884
rect 231762 133764 231768 133816
rect 231820 133804 231826 133816
rect 260374 133804 260380 133816
rect 231820 133776 260380 133804
rect 231820 133764 231826 133776
rect 260374 133764 260380 133776
rect 260432 133764 260438 133816
rect 231210 133560 231216 133612
rect 231268 133600 231274 133612
rect 238294 133600 238300 133612
rect 231268 133572 238300 133600
rect 231268 133560 231274 133572
rect 238294 133560 238300 133572
rect 238352 133560 238358 133612
rect 260190 132812 260196 132864
rect 260248 132852 260254 132864
rect 265066 132852 265072 132864
rect 260248 132824 265072 132852
rect 260248 132812 260254 132824
rect 265066 132812 265072 132824
rect 265124 132812 265130 132864
rect 261846 132744 261852 132796
rect 261904 132784 261910 132796
rect 264974 132784 264980 132796
rect 261904 132756 264980 132784
rect 261904 132744 261910 132756
rect 264974 132744 264980 132756
rect 265032 132744 265038 132796
rect 263134 132608 263140 132660
rect 263192 132648 263198 132660
rect 265894 132648 265900 132660
rect 263192 132620 265900 132648
rect 263192 132608 263198 132620
rect 265894 132608 265900 132620
rect 265952 132608 265958 132660
rect 175918 132540 175924 132592
rect 175976 132580 175982 132592
rect 214006 132580 214012 132592
rect 175976 132552 214012 132580
rect 175976 132540 175982 132552
rect 214006 132540 214012 132552
rect 214064 132540 214070 132592
rect 173250 132472 173256 132524
rect 173308 132512 173314 132524
rect 213914 132512 213920 132524
rect 173308 132484 213920 132512
rect 173308 132472 173314 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 250438 132444 250444 132456
rect 231820 132416 250444 132444
rect 231820 132404 231826 132416
rect 250438 132404 250444 132416
rect 250496 132404 250502 132456
rect 282730 132404 282736 132456
rect 282788 132444 282794 132456
rect 296898 132444 296904 132456
rect 282788 132416 296904 132444
rect 282788 132404 282794 132416
rect 296898 132404 296904 132416
rect 296956 132404 296962 132456
rect 231670 132336 231676 132388
rect 231728 132376 231734 132388
rect 249150 132376 249156 132388
rect 231728 132348 249156 132376
rect 231728 132336 231734 132348
rect 249150 132336 249156 132348
rect 249208 132336 249214 132388
rect 282822 132336 282828 132388
rect 282880 132376 282886 132388
rect 295334 132376 295340 132388
rect 282880 132348 295340 132376
rect 282880 132336 282886 132348
rect 295334 132336 295340 132348
rect 295392 132336 295398 132388
rect 250806 131724 250812 131776
rect 250864 131764 250870 131776
rect 265802 131764 265808 131776
rect 250864 131736 265808 131764
rect 250864 131724 250870 131736
rect 265802 131724 265808 131736
rect 265860 131724 265866 131776
rect 167730 131112 167736 131164
rect 167788 131152 167794 131164
rect 213914 131152 213920 131164
rect 167788 131124 213920 131152
rect 167788 131112 167794 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 258810 131084 258816 131096
rect 231820 131056 258816 131084
rect 231820 131044 231826 131056
rect 258810 131044 258816 131056
rect 258868 131044 258874 131096
rect 282822 131044 282828 131096
rect 282880 131084 282886 131096
rect 307754 131084 307760 131096
rect 282880 131056 307760 131084
rect 282880 131044 282886 131056
rect 307754 131044 307760 131056
rect 307812 131044 307818 131096
rect 231670 130976 231676 131028
rect 231728 131016 231734 131028
rect 257338 131016 257344 131028
rect 231728 130988 257344 131016
rect 231728 130976 231734 130988
rect 257338 130976 257344 130988
rect 257396 130976 257402 131028
rect 282178 130976 282184 131028
rect 282236 131016 282242 131028
rect 300946 131016 300952 131028
rect 282236 130988 300952 131016
rect 282236 130976 282242 130988
rect 300946 130976 300952 130988
rect 301004 130976 301010 131028
rect 231578 130908 231584 130960
rect 231636 130948 231642 130960
rect 254762 130948 254768 130960
rect 231636 130920 254768 130948
rect 231636 130908 231642 130920
rect 254762 130908 254768 130920
rect 254820 130908 254826 130960
rect 210418 129820 210424 129872
rect 210476 129860 210482 129872
rect 214006 129860 214012 129872
rect 210476 129832 214012 129860
rect 210476 129820 210482 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 261662 129820 261668 129872
rect 261720 129860 261726 129872
rect 265066 129860 265072 129872
rect 261720 129832 265072 129860
rect 261720 129820 261726 129832
rect 265066 129820 265072 129832
rect 265124 129820 265130 129872
rect 174630 129752 174636 129804
rect 174688 129792 174694 129804
rect 213914 129792 213920 129804
rect 174688 129764 213920 129792
rect 174688 129752 174694 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 254578 129752 254584 129804
rect 254636 129792 254642 129804
rect 264974 129792 264980 129804
rect 254636 129764 264980 129792
rect 254636 129752 254642 129764
rect 264974 129752 264980 129764
rect 265032 129752 265038 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 253474 129724 253480 129736
rect 231820 129696 253480 129724
rect 231820 129684 231826 129696
rect 253474 129684 253480 129696
rect 253532 129684 253538 129736
rect 231670 129616 231676 129668
rect 231728 129656 231734 129668
rect 244918 129656 244924 129668
rect 231728 129628 244924 129656
rect 231728 129616 231734 129628
rect 244918 129616 244924 129628
rect 244976 129616 244982 129668
rect 231118 129072 231124 129124
rect 231176 129112 231182 129124
rect 242434 129112 242440 129124
rect 231176 129084 242440 129112
rect 231176 129072 231182 129084
rect 242434 129072 242440 129084
rect 242492 129072 242498 129124
rect 231578 129004 231584 129056
rect 231636 129044 231642 129056
rect 246298 129044 246304 129056
rect 231636 129016 246304 129044
rect 231636 129004 231642 129016
rect 246298 129004 246304 129016
rect 246356 129004 246362 129056
rect 204990 128392 204996 128444
rect 205048 128432 205054 128444
rect 213914 128432 213920 128444
rect 205048 128404 213920 128432
rect 205048 128392 205054 128404
rect 213914 128392 213920 128404
rect 213972 128392 213978 128444
rect 257338 128392 257344 128444
rect 257396 128432 257402 128444
rect 265066 128432 265072 128444
rect 257396 128404 265072 128432
rect 257396 128392 257402 128404
rect 265066 128392 265072 128404
rect 265124 128392 265130 128444
rect 59262 128324 59268 128376
rect 59320 128364 59326 128376
rect 66162 128364 66168 128376
rect 59320 128336 66168 128364
rect 59320 128324 59326 128336
rect 66162 128324 66168 128336
rect 66220 128324 66226 128376
rect 170490 128324 170496 128376
rect 170548 128364 170554 128376
rect 214006 128364 214012 128376
rect 170548 128336 214012 128364
rect 170548 128324 170554 128336
rect 214006 128324 214012 128336
rect 214064 128324 214070 128376
rect 246482 128324 246488 128376
rect 246540 128364 246546 128376
rect 264974 128364 264980 128376
rect 246540 128336 264980 128364
rect 246540 128324 246546 128336
rect 264974 128324 264980 128336
rect 265032 128324 265038 128376
rect 230842 128256 230848 128308
rect 230900 128296 230906 128308
rect 261754 128296 261760 128308
rect 230900 128268 261760 128296
rect 230900 128256 230906 128268
rect 261754 128256 261760 128268
rect 261812 128256 261818 128308
rect 281718 128256 281724 128308
rect 281776 128296 281782 128308
rect 295426 128296 295432 128308
rect 281776 128268 295432 128296
rect 281776 128256 281782 128268
rect 295426 128256 295432 128268
rect 295484 128256 295490 128308
rect 231762 128188 231768 128240
rect 231820 128228 231826 128240
rect 260282 128228 260288 128240
rect 231820 128200 260288 128228
rect 231820 128188 231826 128200
rect 260282 128188 260288 128200
rect 260340 128188 260346 128240
rect 282822 128188 282828 128240
rect 282880 128228 282886 128240
rect 289906 128228 289912 128240
rect 282880 128200 289912 128228
rect 282880 128188 282886 128200
rect 289906 128188 289912 128200
rect 289964 128188 289970 128240
rect 231026 127576 231032 127628
rect 231084 127616 231090 127628
rect 239582 127616 239588 127628
rect 231084 127588 239588 127616
rect 231084 127576 231090 127588
rect 239582 127576 239588 127588
rect 239640 127576 239646 127628
rect 253566 127576 253572 127628
rect 253624 127616 253630 127628
rect 265710 127616 265716 127628
rect 253624 127588 265716 127616
rect 253624 127576 253630 127588
rect 265710 127576 265716 127588
rect 265768 127576 265774 127628
rect 202322 127032 202328 127084
rect 202380 127072 202386 127084
rect 213914 127072 213920 127084
rect 202380 127044 213920 127072
rect 202380 127032 202386 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 174538 126964 174544 127016
rect 174596 127004 174602 127016
rect 214006 127004 214012 127016
rect 174596 126976 214012 127004
rect 174596 126964 174602 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 261570 126964 261576 127016
rect 261628 127004 261634 127016
rect 264974 127004 264980 127016
rect 261628 126976 264980 127004
rect 261628 126964 261634 126976
rect 264974 126964 264980 126976
rect 265032 126964 265038 127016
rect 231762 126896 231768 126948
rect 231820 126936 231826 126948
rect 251818 126936 251824 126948
rect 231820 126908 251824 126936
rect 231820 126896 231826 126908
rect 251818 126896 251824 126908
rect 251876 126896 251882 126948
rect 281902 126896 281908 126948
rect 281960 126936 281966 126948
rect 285674 126936 285680 126948
rect 281960 126908 285680 126936
rect 281960 126896 281966 126908
rect 285674 126896 285680 126908
rect 285732 126896 285738 126948
rect 231670 126828 231676 126880
rect 231728 126868 231734 126880
rect 250714 126868 250720 126880
rect 231728 126840 250720 126868
rect 231728 126828 231734 126840
rect 250714 126828 250720 126840
rect 250772 126828 250778 126880
rect 257522 125740 257528 125792
rect 257580 125780 257586 125792
rect 264974 125780 264980 125792
rect 257580 125752 264980 125780
rect 257580 125740 257586 125752
rect 264974 125740 264980 125752
rect 265032 125740 265038 125792
rect 193950 125672 193956 125724
rect 194008 125712 194014 125724
rect 213914 125712 213920 125724
rect 194008 125684 213920 125712
rect 194008 125672 194014 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 254762 125672 254768 125724
rect 254820 125712 254826 125724
rect 265066 125712 265072 125724
rect 254820 125684 265072 125712
rect 254820 125672 254826 125684
rect 265066 125672 265072 125684
rect 265124 125672 265130 125724
rect 167638 125604 167644 125656
rect 167696 125644 167702 125656
rect 214006 125644 214012 125656
rect 167696 125616 214012 125644
rect 167696 125604 167702 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 236914 125604 236920 125656
rect 236972 125644 236978 125656
rect 265158 125644 265164 125656
rect 236972 125616 265164 125644
rect 236972 125604 236978 125616
rect 265158 125604 265164 125616
rect 265216 125604 265222 125656
rect 231486 125536 231492 125588
rect 231544 125576 231550 125588
rect 261478 125576 261484 125588
rect 231544 125548 261484 125576
rect 231544 125536 231550 125548
rect 261478 125536 261484 125548
rect 261536 125536 261542 125588
rect 282822 125536 282828 125588
rect 282880 125576 282886 125588
rect 305178 125576 305184 125588
rect 282880 125548 305184 125576
rect 282880 125536 282886 125548
rect 305178 125536 305184 125548
rect 305236 125536 305242 125588
rect 231762 125468 231768 125520
rect 231820 125508 231826 125520
rect 253290 125508 253296 125520
rect 231820 125480 253296 125508
rect 231820 125468 231826 125480
rect 253290 125468 253296 125480
rect 253348 125468 253354 125520
rect 282730 125468 282736 125520
rect 282788 125508 282794 125520
rect 298186 125508 298192 125520
rect 282788 125480 298192 125508
rect 282788 125468 282794 125480
rect 298186 125468 298192 125480
rect 298244 125468 298250 125520
rect 231762 125060 231768 125112
rect 231820 125100 231826 125112
rect 236822 125100 236828 125112
rect 231820 125072 236828 125100
rect 231820 125060 231826 125072
rect 236822 125060 236828 125072
rect 236880 125060 236886 125112
rect 230934 124584 230940 124636
rect 230992 124624 230998 124636
rect 235534 124624 235540 124636
rect 230992 124596 235540 124624
rect 230992 124584 230998 124596
rect 235534 124584 235540 124596
rect 235592 124584 235598 124636
rect 252186 124312 252192 124364
rect 252244 124352 252250 124364
rect 264974 124352 264980 124364
rect 252244 124324 264980 124352
rect 252244 124312 252250 124324
rect 264974 124312 264980 124324
rect 265032 124312 265038 124364
rect 195422 124244 195428 124296
rect 195480 124284 195486 124296
rect 213914 124284 213920 124296
rect 195480 124256 213920 124284
rect 195480 124244 195486 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 239582 124244 239588 124296
rect 239640 124284 239646 124296
rect 265066 124284 265072 124296
rect 239640 124256 265072 124284
rect 239640 124244 239646 124256
rect 265066 124244 265072 124256
rect 265124 124244 265130 124296
rect 178770 124176 178776 124228
rect 178828 124216 178834 124228
rect 214006 124216 214012 124228
rect 178828 124188 214012 124216
rect 178828 124176 178834 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 235258 124176 235264 124228
rect 235316 124216 235322 124228
rect 265158 124216 265164 124228
rect 235316 124188 265164 124216
rect 235316 124176 235322 124188
rect 265158 124176 265164 124188
rect 265216 124176 265222 124228
rect 230750 124108 230756 124160
rect 230808 124148 230814 124160
rect 232498 124148 232504 124160
rect 230808 124120 232504 124148
rect 230808 124108 230814 124120
rect 232498 124108 232504 124120
rect 232556 124108 232562 124160
rect 282638 124108 282644 124160
rect 282696 124148 282702 124160
rect 306374 124148 306380 124160
rect 282696 124120 306380 124148
rect 282696 124108 282702 124120
rect 306374 124108 306380 124120
rect 306432 124108 306438 124160
rect 282822 124040 282828 124092
rect 282880 124080 282886 124092
rect 295518 124080 295524 124092
rect 282880 124052 295524 124080
rect 282880 124040 282886 124052
rect 295518 124040 295524 124052
rect 295576 124040 295582 124092
rect 230750 123564 230756 123616
rect 230808 123604 230814 123616
rect 238018 123604 238024 123616
rect 230808 123576 238024 123604
rect 230808 123564 230814 123576
rect 238018 123564 238024 123576
rect 238076 123564 238082 123616
rect 282730 123428 282736 123480
rect 282788 123468 282794 123480
rect 303614 123468 303620 123480
rect 282788 123440 303620 123468
rect 282788 123428 282794 123440
rect 303614 123428 303620 123440
rect 303672 123428 303678 123480
rect 250714 122952 250720 123004
rect 250772 122992 250778 123004
rect 264974 122992 264980 123004
rect 250772 122964 264980 122992
rect 250772 122952 250778 122964
rect 264974 122952 264980 122964
rect 265032 122952 265038 123004
rect 173434 122884 173440 122936
rect 173492 122924 173498 122936
rect 214006 122924 214012 122936
rect 173492 122896 214012 122924
rect 173492 122884 173498 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 232682 122884 232688 122936
rect 232740 122924 232746 122936
rect 265066 122924 265072 122936
rect 232740 122896 265072 122924
rect 232740 122884 232746 122896
rect 265066 122884 265072 122896
rect 265124 122884 265130 122936
rect 171778 122816 171784 122868
rect 171836 122856 171842 122868
rect 213914 122856 213920 122868
rect 171836 122828 213920 122856
rect 171836 122816 171842 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 229830 122816 229836 122868
rect 229888 122856 229894 122868
rect 265158 122856 265164 122868
rect 229888 122828 265164 122856
rect 229888 122816 229894 122828
rect 265158 122816 265164 122828
rect 265216 122816 265222 122868
rect 231670 122748 231676 122800
rect 231728 122788 231734 122800
rect 264238 122788 264244 122800
rect 231728 122760 264244 122788
rect 231728 122748 231734 122760
rect 264238 122748 264244 122760
rect 264296 122748 264302 122800
rect 282822 122748 282828 122800
rect 282880 122788 282886 122800
rect 292574 122788 292580 122800
rect 282880 122760 292580 122788
rect 282880 122748 282886 122760
rect 292574 122748 292580 122760
rect 292632 122748 292638 122800
rect 231762 122680 231768 122732
rect 231820 122720 231826 122732
rect 242342 122720 242348 122732
rect 231820 122692 242348 122720
rect 231820 122680 231826 122692
rect 242342 122680 242348 122692
rect 242400 122680 242406 122732
rect 231670 122068 231676 122120
rect 231728 122108 231734 122120
rect 243722 122108 243728 122120
rect 231728 122080 243728 122108
rect 231728 122068 231734 122080
rect 243722 122068 243728 122080
rect 243780 122068 243786 122120
rect 256326 121592 256332 121644
rect 256384 121632 256390 121644
rect 265066 121632 265072 121644
rect 256384 121604 265072 121632
rect 256384 121592 256390 121604
rect 265066 121592 265072 121604
rect 265124 121592 265130 121644
rect 206462 121524 206468 121576
rect 206520 121564 206526 121576
rect 213914 121564 213920 121576
rect 206520 121536 213920 121564
rect 206520 121524 206526 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 246298 121524 246304 121576
rect 246356 121564 246362 121576
rect 264974 121564 264980 121576
rect 246356 121536 264980 121564
rect 246356 121524 246362 121536
rect 264974 121524 264980 121536
rect 265032 121524 265038 121576
rect 63402 121456 63408 121508
rect 63460 121496 63466 121508
rect 65978 121496 65984 121508
rect 63460 121468 65984 121496
rect 63460 121456 63466 121468
rect 65978 121456 65984 121468
rect 66036 121456 66042 121508
rect 203518 121456 203524 121508
rect 203576 121496 203582 121508
rect 214006 121496 214012 121508
rect 203576 121468 214012 121496
rect 203576 121456 203582 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 243630 121456 243636 121508
rect 243688 121496 243694 121508
rect 265158 121496 265164 121508
rect 243688 121468 265164 121496
rect 243688 121456 243694 121468
rect 265158 121456 265164 121468
rect 265216 121456 265222 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 247862 121428 247868 121440
rect 231820 121400 247868 121428
rect 231820 121388 231826 121400
rect 247862 121388 247868 121400
rect 247920 121388 247926 121440
rect 281534 121320 281540 121372
rect 281592 121360 281598 121372
rect 284386 121360 284392 121372
rect 281592 121332 284392 121360
rect 281592 121320 281598 121332
rect 284386 121320 284392 121332
rect 284444 121320 284450 121372
rect 231578 121252 231584 121304
rect 231636 121292 231642 121304
rect 234154 121292 234160 121304
rect 231636 121264 234160 121292
rect 231636 121252 231642 121264
rect 234154 121252 234160 121264
rect 234212 121252 234218 121304
rect 230750 120708 230756 120760
rect 230808 120748 230814 120760
rect 257614 120748 257620 120760
rect 230808 120720 257620 120748
rect 230808 120708 230814 120720
rect 257614 120708 257620 120720
rect 257672 120708 257678 120760
rect 242526 120232 242532 120284
rect 242584 120272 242590 120284
rect 264974 120272 264980 120284
rect 242584 120244 264980 120272
rect 242584 120232 242590 120244
rect 264974 120232 264980 120244
rect 265032 120232 265038 120284
rect 207658 120164 207664 120216
rect 207716 120204 207722 120216
rect 214006 120204 214012 120216
rect 207716 120176 214012 120204
rect 207716 120164 207722 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 238294 120164 238300 120216
rect 238352 120204 238358 120216
rect 265158 120204 265164 120216
rect 238352 120176 265164 120204
rect 238352 120164 238358 120176
rect 265158 120164 265164 120176
rect 265216 120164 265222 120216
rect 62022 120096 62028 120148
rect 62080 120136 62086 120148
rect 65886 120136 65892 120148
rect 62080 120108 65892 120136
rect 62080 120096 62086 120108
rect 65886 120096 65892 120108
rect 65944 120096 65950 120148
rect 196802 120096 196808 120148
rect 196860 120136 196866 120148
rect 213914 120136 213920 120148
rect 196860 120108 213920 120136
rect 196860 120096 196866 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 232498 120096 232504 120148
rect 232556 120136 232562 120148
rect 265066 120136 265072 120148
rect 232556 120108 265072 120136
rect 232556 120096 232562 120108
rect 265066 120096 265072 120108
rect 265124 120096 265130 120148
rect 230934 120028 230940 120080
rect 230992 120068 230998 120080
rect 260098 120068 260104 120080
rect 230992 120040 260104 120068
rect 230992 120028 230998 120040
rect 260098 120028 260104 120040
rect 260156 120028 260162 120080
rect 282086 120028 282092 120080
rect 282144 120068 282150 120080
rect 291286 120068 291292 120080
rect 282144 120040 291292 120068
rect 282144 120028 282150 120040
rect 291286 120028 291292 120040
rect 291344 120028 291350 120080
rect 231394 119960 231400 120012
rect 231452 120000 231458 120012
rect 240870 120000 240876 120012
rect 231452 119972 240876 120000
rect 231452 119960 231458 119972
rect 240870 119960 240876 119972
rect 240928 119960 240934 120012
rect 209222 118804 209228 118856
rect 209280 118844 209286 118856
rect 213914 118844 213920 118856
rect 209280 118816 213920 118844
rect 209280 118804 209286 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 193858 118736 193864 118788
rect 193916 118776 193922 118788
rect 214098 118776 214104 118788
rect 193916 118748 214104 118776
rect 193916 118736 193922 118748
rect 214098 118736 214104 118748
rect 214156 118736 214162 118788
rect 192478 118668 192484 118720
rect 192536 118708 192542 118720
rect 214006 118708 214012 118720
rect 192536 118680 214012 118708
rect 192536 118668 192542 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 231302 118668 231308 118720
rect 231360 118708 231366 118720
rect 232774 118708 232780 118720
rect 231360 118680 232780 118708
rect 231360 118668 231366 118680
rect 232774 118668 232780 118680
rect 232832 118668 232838 118720
rect 258810 118668 258816 118720
rect 258868 118708 258874 118720
rect 264974 118708 264980 118720
rect 258868 118680 264980 118708
rect 258868 118668 258874 118680
rect 264974 118668 264980 118680
rect 265032 118668 265038 118720
rect 231486 118600 231492 118652
rect 231544 118640 231550 118652
rect 258902 118640 258908 118652
rect 231544 118612 258908 118640
rect 231544 118600 231550 118612
rect 258902 118600 258908 118612
rect 258960 118600 258966 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 289814 118640 289820 118652
rect 282880 118612 289820 118640
rect 282880 118600 282886 118612
rect 289814 118600 289820 118612
rect 289872 118600 289878 118652
rect 231762 118532 231768 118584
rect 231820 118572 231826 118584
rect 258718 118572 258724 118584
rect 231820 118544 258724 118572
rect 231820 118532 231826 118544
rect 258718 118532 258724 118544
rect 258776 118532 258782 118584
rect 282730 118532 282736 118584
rect 282788 118572 282794 118584
rect 288710 118572 288716 118584
rect 282788 118544 288716 118572
rect 282788 118532 282794 118544
rect 288710 118532 288716 118544
rect 288768 118532 288774 118584
rect 231670 118396 231676 118448
rect 231728 118436 231734 118448
rect 236730 118436 236736 118448
rect 231728 118408 236736 118436
rect 231728 118396 231734 118408
rect 236730 118396 236736 118408
rect 236788 118396 236794 118448
rect 189810 117376 189816 117428
rect 189868 117416 189874 117428
rect 214006 117416 214012 117428
rect 189868 117388 214012 117416
rect 189868 117376 189874 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 261478 117376 261484 117428
rect 261536 117416 261542 117428
rect 265066 117416 265072 117428
rect 261536 117388 265072 117416
rect 261536 117376 261542 117388
rect 265066 117376 265072 117388
rect 265124 117376 265130 117428
rect 171870 117308 171876 117360
rect 171928 117348 171934 117360
rect 213914 117348 213920 117360
rect 171928 117320 213920 117348
rect 171928 117308 171934 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 247862 117308 247868 117360
rect 247920 117348 247926 117360
rect 264974 117348 264980 117360
rect 247920 117320 264980 117348
rect 247920 117308 247926 117320
rect 264974 117308 264980 117320
rect 265032 117308 265038 117360
rect 231762 117240 231768 117292
rect 231820 117280 231826 117292
rect 254854 117280 254860 117292
rect 231820 117252 254860 117280
rect 231820 117240 231826 117252
rect 254854 117240 254860 117252
rect 254912 117240 254918 117292
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 298278 117280 298284 117292
rect 282880 117252 298284 117280
rect 282880 117240 282886 117252
rect 298278 117240 298284 117252
rect 298336 117240 298342 117292
rect 282730 117172 282736 117224
rect 282788 117212 282794 117224
rect 288526 117212 288532 117224
rect 282788 117184 288532 117212
rect 282788 117172 282794 117184
rect 288526 117172 288532 117184
rect 288584 117172 288590 117224
rect 230658 116968 230664 117020
rect 230716 117008 230722 117020
rect 234062 117008 234068 117020
rect 230716 116980 234068 117008
rect 230716 116968 230722 116980
rect 234062 116968 234068 116980
rect 234120 116968 234126 117020
rect 234154 116560 234160 116612
rect 234212 116600 234218 116612
rect 261846 116600 261852 116612
rect 234212 116572 261852 116600
rect 234212 116560 234218 116572
rect 261846 116560 261852 116572
rect 261904 116560 261910 116612
rect 253474 116152 253480 116204
rect 253532 116192 253538 116204
rect 264974 116192 264980 116204
rect 253532 116164 264980 116192
rect 253532 116152 253538 116164
rect 264974 116152 264980 116164
rect 265032 116152 265038 116204
rect 260098 116084 260104 116136
rect 260156 116124 260162 116136
rect 265158 116124 265164 116136
rect 260156 116096 265164 116124
rect 260156 116084 260162 116096
rect 265158 116084 265164 116096
rect 265216 116084 265222 116136
rect 258718 116016 258724 116068
rect 258776 116056 258782 116068
rect 264974 116056 264980 116068
rect 258776 116028 264980 116056
rect 258776 116016 258782 116028
rect 264974 116016 264980 116028
rect 265032 116016 265038 116068
rect 181530 115948 181536 116000
rect 181588 115988 181594 116000
rect 213914 115988 213920 116000
rect 181588 115960 213920 115988
rect 181588 115948 181594 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 262950 115948 262956 116000
rect 263008 115988 263014 116000
rect 265066 115988 265072 116000
rect 263008 115960 265072 115988
rect 263008 115948 263014 115960
rect 265066 115948 265072 115960
rect 265124 115948 265130 116000
rect 231762 115880 231768 115932
rect 231820 115920 231826 115932
rect 255958 115920 255964 115932
rect 231820 115892 255964 115920
rect 231820 115880 231826 115892
rect 255958 115880 255964 115892
rect 256016 115880 256022 115932
rect 281718 115880 281724 115932
rect 281776 115920 281782 115932
rect 309134 115920 309140 115932
rect 281776 115892 309140 115920
rect 281776 115880 281782 115892
rect 309134 115880 309140 115892
rect 309192 115880 309198 115932
rect 231670 115812 231676 115864
rect 231728 115852 231734 115864
rect 249334 115852 249340 115864
rect 231728 115824 249340 115852
rect 231728 115812 231734 115824
rect 249334 115812 249340 115824
rect 249392 115812 249398 115864
rect 282086 115812 282092 115864
rect 282144 115852 282150 115864
rect 296714 115852 296720 115864
rect 282144 115824 296720 115852
rect 282144 115812 282150 115824
rect 296714 115812 296720 115824
rect 296772 115812 296778 115864
rect 231762 115268 231768 115320
rect 231820 115308 231826 115320
rect 239674 115308 239680 115320
rect 231820 115280 239680 115308
rect 231820 115268 231826 115280
rect 239674 115268 239680 115280
rect 239732 115268 239738 115320
rect 230014 115200 230020 115252
rect 230072 115240 230078 115252
rect 267274 115240 267280 115252
rect 230072 115212 267280 115240
rect 230072 115200 230078 115212
rect 267274 115200 267280 115212
rect 267332 115200 267338 115252
rect 185670 114588 185676 114640
rect 185728 114628 185734 114640
rect 214006 114628 214012 114640
rect 185728 114600 214012 114628
rect 185728 114588 185734 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 177574 114520 177580 114572
rect 177632 114560 177638 114572
rect 213914 114560 213920 114572
rect 177632 114532 213920 114560
rect 177632 114520 177638 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 249150 114520 249156 114572
rect 249208 114560 249214 114572
rect 264974 114560 264980 114572
rect 249208 114532 264980 114560
rect 249208 114520 249214 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 231486 114452 231492 114504
rect 231544 114492 231550 114504
rect 253382 114492 253388 114504
rect 231544 114464 253388 114492
rect 231544 114452 231550 114464
rect 253382 114452 253388 114464
rect 253440 114452 253446 114504
rect 282822 114452 282828 114504
rect 282880 114492 282886 114504
rect 302326 114492 302332 114504
rect 282880 114464 302332 114492
rect 282880 114452 282886 114464
rect 302326 114452 302332 114464
rect 302384 114452 302390 114504
rect 282730 114384 282736 114436
rect 282788 114424 282794 114436
rect 299566 114424 299572 114436
rect 282788 114396 299572 114424
rect 282788 114384 282794 114396
rect 299566 114384 299572 114396
rect 299624 114384 299630 114436
rect 230842 113772 230848 113824
rect 230900 113812 230906 113824
rect 263042 113812 263048 113824
rect 230900 113784 263048 113812
rect 230900 113772 230906 113784
rect 263042 113772 263048 113784
rect 263100 113772 263106 113824
rect 200850 113228 200856 113280
rect 200908 113268 200914 113280
rect 214006 113268 214012 113280
rect 200908 113240 214012 113268
rect 200908 113228 200914 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 196710 113160 196716 113212
rect 196768 113200 196774 113212
rect 213914 113200 213920 113212
rect 196768 113172 213920 113200
rect 196768 113160 196774 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 252002 113132 252008 113144
rect 231820 113104 252008 113132
rect 231820 113092 231826 113104
rect 252002 113092 252008 113104
rect 252060 113092 252066 113144
rect 282086 113092 282092 113144
rect 282144 113132 282150 113144
rect 300854 113132 300860 113144
rect 282144 113104 300860 113132
rect 282144 113092 282150 113104
rect 300854 113092 300860 113104
rect 300912 113092 300918 113144
rect 231670 113024 231676 113076
rect 231728 113064 231734 113076
rect 250622 113064 250628 113076
rect 231728 113036 250628 113064
rect 231728 113024 231734 113036
rect 250622 113024 250628 113036
rect 250680 113024 250686 113076
rect 258902 111936 258908 111988
rect 258960 111976 258966 111988
rect 265158 111976 265164 111988
rect 258960 111948 265164 111976
rect 258960 111936 258966 111948
rect 265158 111936 265164 111948
rect 265216 111936 265222 111988
rect 211798 111868 211804 111920
rect 211856 111908 211862 111920
rect 214006 111908 214012 111920
rect 211856 111880 214012 111908
rect 211856 111868 211862 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 251818 111868 251824 111920
rect 251876 111908 251882 111920
rect 264974 111908 264980 111920
rect 251876 111880 264980 111908
rect 251876 111868 251882 111880
rect 264974 111868 264980 111880
rect 265032 111868 265038 111920
rect 169110 111800 169116 111852
rect 169168 111840 169174 111852
rect 213914 111840 213920 111852
rect 169168 111812 213920 111840
rect 169168 111800 169174 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 244918 111800 244924 111852
rect 244976 111840 244982 111852
rect 265066 111840 265072 111852
rect 244976 111812 265072 111840
rect 244976 111800 244982 111812
rect 265066 111800 265072 111812
rect 265124 111800 265130 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 22738 111772 22744 111784
rect 3200 111744 22744 111772
rect 3200 111732 3206 111744
rect 22738 111732 22744 111744
rect 22796 111732 22802 111784
rect 167822 111732 167828 111784
rect 167880 111772 167886 111784
rect 197998 111772 198004 111784
rect 167880 111744 198004 111772
rect 167880 111732 167886 111744
rect 197998 111732 198004 111744
rect 198056 111732 198062 111784
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 251910 111772 251916 111784
rect 231820 111744 251916 111772
rect 231820 111732 231826 111744
rect 251910 111732 251916 111744
rect 251968 111732 251974 111784
rect 282730 111732 282736 111784
rect 282788 111772 282794 111784
rect 303706 111772 303712 111784
rect 282788 111744 303712 111772
rect 282788 111732 282794 111744
rect 303706 111732 303712 111744
rect 303764 111732 303770 111784
rect 230566 111664 230572 111716
rect 230624 111704 230630 111716
rect 246574 111704 246580 111716
rect 230624 111676 246580 111704
rect 230624 111664 230630 111676
rect 246574 111664 246580 111676
rect 246632 111664 246638 111716
rect 282822 111664 282828 111716
rect 282880 111704 282886 111716
rect 298094 111704 298100 111716
rect 282880 111676 298100 111704
rect 282880 111664 282886 111676
rect 298094 111664 298100 111676
rect 298152 111664 298158 111716
rect 231302 111052 231308 111104
rect 231360 111092 231366 111104
rect 260466 111092 260472 111104
rect 231360 111064 260472 111092
rect 231360 111052 231366 111064
rect 260466 111052 260472 111064
rect 260524 111052 260530 111104
rect 260374 110576 260380 110628
rect 260432 110616 260438 110628
rect 265158 110616 265164 110628
rect 260432 110588 265164 110616
rect 260432 110576 260438 110588
rect 265158 110576 265164 110588
rect 265216 110576 265222 110628
rect 178862 110508 178868 110560
rect 178920 110548 178926 110560
rect 213914 110548 213920 110560
rect 178920 110520 213920 110548
rect 178920 110508 178926 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 256142 110508 256148 110560
rect 256200 110548 256206 110560
rect 264974 110548 264980 110560
rect 256200 110520 264980 110548
rect 256200 110508 256206 110520
rect 264974 110508 264980 110520
rect 265032 110508 265038 110560
rect 177482 110440 177488 110492
rect 177540 110480 177546 110492
rect 214006 110480 214012 110492
rect 177540 110452 214012 110480
rect 177540 110440 177546 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 236730 110440 236736 110492
rect 236788 110480 236794 110492
rect 265066 110480 265072 110492
rect 236788 110452 265072 110480
rect 236788 110440 236794 110452
rect 265066 110440 265072 110452
rect 265124 110440 265130 110492
rect 167822 110372 167828 110424
rect 167880 110412 167886 110424
rect 215294 110412 215300 110424
rect 167880 110384 215300 110412
rect 167880 110372 167886 110384
rect 215294 110372 215300 110384
rect 215352 110372 215358 110424
rect 231670 110372 231676 110424
rect 231728 110412 231734 110424
rect 264422 110412 264428 110424
rect 231728 110384 264428 110412
rect 231728 110372 231734 110384
rect 264422 110372 264428 110384
rect 264480 110372 264486 110424
rect 282086 110372 282092 110424
rect 282144 110412 282150 110424
rect 302234 110412 302240 110424
rect 282144 110384 302240 110412
rect 282144 110372 282150 110384
rect 302234 110372 302240 110384
rect 302292 110372 302298 110424
rect 230566 110304 230572 110356
rect 230624 110344 230630 110356
rect 262858 110344 262864 110356
rect 230624 110316 262864 110344
rect 230624 110304 230630 110316
rect 262858 110304 262864 110316
rect 262916 110304 262922 110356
rect 282270 110304 282276 110356
rect 282328 110344 282334 110356
rect 292666 110344 292672 110356
rect 282328 110316 292672 110344
rect 282328 110304 282334 110316
rect 292666 110304 292672 110316
rect 292724 110304 292730 110356
rect 231762 110236 231768 110288
rect 231820 110276 231826 110288
rect 245102 110276 245108 110288
rect 231820 110248 245108 110276
rect 231820 110236 231826 110248
rect 245102 110236 245108 110248
rect 245160 110236 245166 110288
rect 260282 109148 260288 109200
rect 260340 109188 260346 109200
rect 265158 109188 265164 109200
rect 260340 109160 265164 109188
rect 260340 109148 260346 109160
rect 265158 109148 265164 109160
rect 265216 109148 265222 109200
rect 198182 109080 198188 109132
rect 198240 109120 198246 109132
rect 214006 109120 214012 109132
rect 198240 109092 214012 109120
rect 198240 109080 198246 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 253290 109080 253296 109132
rect 253348 109120 253354 109132
rect 264974 109120 264980 109132
rect 253348 109092 264980 109120
rect 253348 109080 253354 109092
rect 264974 109080 264980 109092
rect 265032 109080 265038 109132
rect 166442 109012 166448 109064
rect 166500 109052 166506 109064
rect 213914 109052 213920 109064
rect 166500 109024 213920 109052
rect 166500 109012 166506 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 238018 109012 238024 109064
rect 238076 109052 238082 109064
rect 265066 109052 265072 109064
rect 238076 109024 265072 109052
rect 238076 109012 238082 109024
rect 265066 109012 265072 109024
rect 265124 109012 265130 109064
rect 167822 108944 167828 108996
rect 167880 108984 167886 108996
rect 200758 108984 200764 108996
rect 167880 108956 200764 108984
rect 167880 108944 167886 108956
rect 200758 108944 200764 108956
rect 200816 108944 200822 108996
rect 231762 108944 231768 108996
rect 231820 108984 231826 108996
rect 249058 108984 249064 108996
rect 231820 108956 249064 108984
rect 231820 108944 231826 108956
rect 249058 108944 249064 108956
rect 249116 108944 249122 108996
rect 281718 108944 281724 108996
rect 281776 108984 281782 108996
rect 303798 108984 303804 108996
rect 281776 108956 303804 108984
rect 281776 108944 281782 108956
rect 303798 108944 303804 108956
rect 303856 108944 303862 108996
rect 282086 108876 282092 108928
rect 282144 108916 282150 108928
rect 293954 108916 293960 108928
rect 282144 108888 293960 108916
rect 282144 108876 282150 108888
rect 293954 108876 293960 108888
rect 294012 108876 294018 108928
rect 231486 108604 231492 108656
rect 231544 108644 231550 108656
rect 235442 108644 235448 108656
rect 231544 108616 235448 108644
rect 231544 108604 231550 108616
rect 235442 108604 235448 108616
rect 235500 108604 235506 108656
rect 231394 108264 231400 108316
rect 231452 108304 231458 108316
rect 241054 108304 241060 108316
rect 231452 108276 241060 108304
rect 231452 108264 231458 108276
rect 241054 108264 241060 108276
rect 241112 108264 241118 108316
rect 241146 107856 241152 107908
rect 241204 107896 241210 107908
rect 265066 107896 265072 107908
rect 241204 107868 265072 107896
rect 241204 107856 241210 107868
rect 265066 107856 265072 107868
rect 265124 107856 265130 107908
rect 246574 107788 246580 107840
rect 246632 107828 246638 107840
rect 264974 107828 264980 107840
rect 246632 107800 264980 107828
rect 246632 107788 246638 107800
rect 264974 107788 264980 107800
rect 265032 107788 265038 107840
rect 191282 107720 191288 107772
rect 191340 107760 191346 107772
rect 214006 107760 214012 107772
rect 191340 107732 214012 107760
rect 191340 107720 191346 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 243722 107720 243728 107772
rect 243780 107760 243786 107772
rect 265158 107760 265164 107772
rect 243780 107732 265164 107760
rect 243780 107720 243786 107732
rect 265158 107720 265164 107732
rect 265216 107720 265222 107772
rect 167822 107652 167828 107704
rect 167880 107692 167886 107704
rect 213914 107692 213920 107704
rect 167880 107664 213920 107692
rect 167880 107652 167886 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 231486 107584 231492 107636
rect 231544 107624 231550 107636
rect 256050 107624 256056 107636
rect 231544 107596 256056 107624
rect 231544 107584 231550 107596
rect 256050 107584 256056 107596
rect 256108 107584 256114 107636
rect 231762 107516 231768 107568
rect 231820 107556 231826 107568
rect 253198 107556 253204 107568
rect 231820 107528 253204 107556
rect 231820 107516 231826 107528
rect 253198 107516 253204 107528
rect 253256 107516 253262 107568
rect 169202 106904 169208 106956
rect 169260 106944 169266 106956
rect 214650 106944 214656 106956
rect 169260 106916 214656 106944
rect 169260 106904 169266 106916
rect 214650 106904 214656 106916
rect 214708 106904 214714 106956
rect 231210 106904 231216 106956
rect 231268 106944 231274 106956
rect 246390 106944 246396 106956
rect 231268 106916 246396 106944
rect 231268 106904 231274 106916
rect 246390 106904 246396 106916
rect 246448 106904 246454 106956
rect 242342 106428 242348 106480
rect 242400 106468 242406 106480
rect 264974 106468 264980 106480
rect 242400 106440 264980 106468
rect 242400 106428 242406 106440
rect 264974 106428 264980 106440
rect 265032 106428 265038 106480
rect 199378 106360 199384 106412
rect 199436 106400 199442 106412
rect 214006 106400 214012 106412
rect 199436 106372 214012 106400
rect 199436 106360 199442 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 249058 106360 249064 106412
rect 249116 106400 249122 106412
rect 265066 106400 265072 106412
rect 249116 106372 265072 106400
rect 249116 106360 249122 106372
rect 265066 106360 265072 106372
rect 265124 106360 265130 106412
rect 182910 106292 182916 106344
rect 182968 106332 182974 106344
rect 213914 106332 213920 106344
rect 182968 106304 213920 106332
rect 182968 106292 182974 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 231670 106224 231676 106276
rect 231728 106264 231734 106276
rect 250806 106264 250812 106276
rect 231728 106236 250812 106264
rect 231728 106224 231734 106236
rect 250806 106224 250812 106236
rect 250864 106224 250870 106276
rect 281534 106224 281540 106276
rect 281592 106264 281598 106276
rect 284478 106264 284484 106276
rect 281592 106236 284484 106264
rect 281592 106224 281598 106236
rect 284478 106224 284484 106236
rect 284536 106224 284542 106276
rect 231762 106156 231768 106208
rect 231820 106196 231826 106208
rect 250530 106196 250536 106208
rect 231820 106168 250536 106196
rect 231820 106156 231826 106168
rect 250530 106156 250536 106168
rect 250588 106156 250594 106208
rect 230566 106088 230572 106140
rect 230624 106128 230630 106140
rect 245194 106128 245200 106140
rect 230624 106100 245200 106128
rect 230624 106088 230630 106100
rect 245194 106088 245200 106100
rect 245252 106088 245258 106140
rect 258994 105000 259000 105052
rect 259052 105040 259058 105052
rect 265066 105040 265072 105052
rect 259052 105012 265072 105040
rect 259052 105000 259058 105012
rect 265066 105000 265072 105012
rect 265124 105000 265130 105052
rect 184382 104932 184388 104984
rect 184440 104972 184446 104984
rect 214006 104972 214012 104984
rect 184440 104944 214012 104972
rect 184440 104932 184446 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 263042 104932 263048 104984
rect 263100 104972 263106 104984
rect 265434 104972 265440 104984
rect 263100 104944 265440 104972
rect 263100 104932 263106 104944
rect 265434 104932 265440 104944
rect 265492 104932 265498 104984
rect 180150 104864 180156 104916
rect 180208 104904 180214 104916
rect 213914 104904 213920 104916
rect 180208 104876 213920 104904
rect 180208 104864 180214 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 250438 104864 250444 104916
rect 250496 104904 250502 104916
rect 264974 104904 264980 104916
rect 250496 104876 264980 104904
rect 250496 104864 250502 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 282822 104796 282828 104848
rect 282880 104836 282886 104848
rect 305086 104836 305092 104848
rect 282880 104808 305092 104836
rect 282880 104796 282886 104808
rect 305086 104796 305092 104808
rect 305144 104796 305150 104848
rect 230842 104728 230848 104780
rect 230900 104768 230906 104780
rect 232590 104768 232596 104780
rect 230900 104740 232596 104768
rect 230900 104728 230906 104740
rect 232590 104728 232596 104740
rect 232648 104728 232654 104780
rect 231762 104660 231768 104712
rect 231820 104700 231826 104712
rect 249242 104700 249248 104712
rect 231820 104672 249248 104700
rect 231820 104660 231826 104672
rect 249242 104660 249248 104672
rect 249300 104660 249306 104712
rect 230750 104184 230756 104236
rect 230808 104224 230814 104236
rect 256234 104224 256240 104236
rect 230808 104196 256240 104224
rect 230808 104184 230814 104196
rect 256234 104184 256240 104196
rect 256292 104184 256298 104236
rect 235442 104116 235448 104168
rect 235500 104156 235506 104168
rect 262950 104156 262956 104168
rect 235500 104128 262956 104156
rect 235500 104116 235506 104128
rect 262950 104116 262956 104128
rect 263008 104116 263014 104168
rect 231486 103844 231492 103896
rect 231544 103884 231550 103896
rect 235350 103884 235356 103896
rect 231544 103856 235356 103884
rect 231544 103844 231550 103856
rect 235350 103844 235356 103856
rect 235408 103844 235414 103896
rect 256050 103640 256056 103692
rect 256108 103680 256114 103692
rect 265066 103680 265072 103692
rect 256108 103652 265072 103680
rect 256108 103640 256114 103652
rect 265066 103640 265072 103652
rect 265124 103640 265130 103692
rect 253198 103572 253204 103624
rect 253256 103612 253262 103624
rect 265158 103612 265164 103624
rect 253256 103584 265164 103612
rect 253256 103572 253262 103584
rect 265158 103572 265164 103584
rect 265216 103572 265222 103624
rect 170582 103504 170588 103556
rect 170640 103544 170646 103556
rect 213914 103544 213920 103556
rect 170640 103516 213920 103544
rect 170640 103504 170646 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 249334 103504 249340 103556
rect 249392 103544 249398 103556
rect 264974 103544 264980 103556
rect 249392 103516 264980 103544
rect 249392 103504 249398 103516
rect 264974 103504 264980 103516
rect 265032 103504 265038 103556
rect 231762 103436 231768 103488
rect 231820 103476 231826 103488
rect 247770 103476 247776 103488
rect 231820 103448 247776 103476
rect 231820 103436 231826 103448
rect 247770 103436 247776 103448
rect 247828 103436 247834 103488
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 299474 103476 299480 103488
rect 282880 103448 299480 103476
rect 282880 103436 282886 103448
rect 299474 103436 299480 103448
rect 299532 103436 299538 103488
rect 231670 103368 231676 103420
rect 231728 103408 231734 103420
rect 242158 103408 242164 103420
rect 231728 103380 242164 103408
rect 231728 103368 231734 103380
rect 242158 103368 242164 103380
rect 242216 103368 242222 103420
rect 231578 103300 231584 103352
rect 231636 103340 231642 103352
rect 242250 103340 242256 103352
rect 231636 103312 242256 103340
rect 231636 103300 231642 103312
rect 242250 103300 242256 103312
rect 242308 103300 242314 103352
rect 240870 102348 240876 102400
rect 240928 102388 240934 102400
rect 265066 102388 265072 102400
rect 240928 102360 265072 102388
rect 240928 102348 240934 102360
rect 265066 102348 265072 102360
rect 265124 102348 265130 102400
rect 255958 102280 255964 102332
rect 256016 102320 256022 102332
rect 264974 102320 264980 102332
rect 256016 102292 264980 102320
rect 256016 102280 256022 102292
rect 264974 102280 264980 102292
rect 265032 102280 265038 102332
rect 242434 102212 242440 102264
rect 242492 102252 242498 102264
rect 265158 102252 265164 102264
rect 242492 102224 265164 102252
rect 242492 102212 242498 102224
rect 265158 102212 265164 102224
rect 265216 102212 265222 102264
rect 195514 102144 195520 102196
rect 195572 102184 195578 102196
rect 213914 102184 213920 102196
rect 195572 102156 213920 102184
rect 195572 102144 195578 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 262858 102144 262864 102196
rect 262916 102184 262922 102196
rect 265250 102184 265256 102196
rect 262916 102156 265256 102184
rect 262916 102144 262922 102156
rect 265250 102144 265256 102156
rect 265308 102144 265314 102196
rect 231762 102076 231768 102128
rect 231820 102116 231826 102128
rect 253566 102116 253572 102128
rect 231820 102088 253572 102116
rect 231820 102076 231826 102088
rect 253566 102076 253572 102088
rect 253624 102076 253630 102128
rect 231670 101396 231676 101448
rect 231728 101436 231734 101448
rect 252094 101436 252100 101448
rect 231728 101408 252100 101436
rect 231728 101396 231734 101408
rect 252094 101396 252100 101408
rect 252152 101396 252158 101448
rect 261294 100852 261300 100904
rect 261352 100892 261358 100904
rect 265066 100892 265072 100904
rect 261352 100864 265072 100892
rect 261352 100852 261358 100864
rect 265066 100852 265072 100864
rect 265124 100852 265130 100904
rect 262950 100784 262956 100836
rect 263008 100824 263014 100836
rect 265342 100824 265348 100836
rect 263008 100796 265348 100824
rect 263008 100784 263014 100796
rect 265342 100784 265348 100796
rect 265400 100784 265406 100836
rect 176010 100716 176016 100768
rect 176068 100756 176074 100768
rect 213914 100756 213920 100768
rect 176068 100728 213920 100756
rect 176068 100716 176074 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 249242 100716 249248 100768
rect 249300 100756 249306 100768
rect 264974 100756 264980 100768
rect 249300 100728 264980 100756
rect 249300 100716 249306 100728
rect 264974 100716 264980 100728
rect 265032 100716 265038 100768
rect 231578 100648 231584 100700
rect 231636 100688 231642 100700
rect 263134 100688 263140 100700
rect 231636 100660 263140 100688
rect 231636 100648 231642 100660
rect 263134 100648 263140 100660
rect 263192 100648 263198 100700
rect 281718 100648 281724 100700
rect 281776 100688 281782 100700
rect 291378 100688 291384 100700
rect 281776 100660 291384 100688
rect 281776 100648 281782 100660
rect 291378 100648 291384 100660
rect 291436 100648 291442 100700
rect 231118 100580 231124 100632
rect 231176 100620 231182 100632
rect 238202 100620 238208 100632
rect 231176 100592 238208 100620
rect 231176 100580 231182 100592
rect 238202 100580 238208 100592
rect 238260 100580 238266 100632
rect 230658 99968 230664 100020
rect 230716 100008 230722 100020
rect 240962 100008 240968 100020
rect 230716 99980 240968 100008
rect 230716 99968 230722 99980
rect 240962 99968 240968 99980
rect 241020 99968 241026 100020
rect 169294 99424 169300 99476
rect 169352 99464 169358 99476
rect 214006 99464 214012 99476
rect 169352 99436 214012 99464
rect 169352 99424 169358 99436
rect 214006 99424 214012 99436
rect 214064 99424 214070 99476
rect 250530 99424 250536 99476
rect 250588 99464 250594 99476
rect 265066 99464 265072 99476
rect 250588 99436 265072 99464
rect 250588 99424 250594 99436
rect 265066 99424 265072 99436
rect 265124 99424 265130 99476
rect 166534 99356 166540 99408
rect 166592 99396 166598 99408
rect 213914 99396 213920 99408
rect 166592 99368 213920 99396
rect 166592 99356 166598 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 242158 99356 242164 99408
rect 242216 99396 242222 99408
rect 264974 99396 264980 99408
rect 242216 99368 264980 99396
rect 242216 99356 242222 99368
rect 264974 99356 264980 99368
rect 265032 99356 265038 99408
rect 231118 99288 231124 99340
rect 231176 99328 231182 99340
rect 233878 99328 233884 99340
rect 231176 99300 233884 99328
rect 231176 99288 231182 99300
rect 233878 99288 233884 99300
rect 233936 99288 233942 99340
rect 282822 99288 282828 99340
rect 282880 99328 282886 99340
rect 309226 99328 309232 99340
rect 282880 99300 309232 99328
rect 282880 99288 282886 99300
rect 309226 99288 309232 99300
rect 309284 99288 309290 99340
rect 203610 98064 203616 98116
rect 203668 98104 203674 98116
rect 213914 98104 213920 98116
rect 203668 98076 213920 98104
rect 203668 98064 203674 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 245102 98064 245108 98116
rect 245160 98104 245166 98116
rect 264974 98104 264980 98116
rect 245160 98076 264980 98104
rect 245160 98064 245166 98076
rect 264974 98064 264980 98076
rect 265032 98064 265038 98116
rect 164878 97996 164884 98048
rect 164936 98036 164942 98048
rect 214006 98036 214012 98048
rect 164936 98008 214012 98036
rect 164936 97996 164942 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 231210 97996 231216 98048
rect 231268 98036 231274 98048
rect 265066 98036 265072 98048
rect 231268 98008 265072 98036
rect 231268 97996 231274 98008
rect 265066 97996 265072 98008
rect 265124 97996 265130 98048
rect 282178 97928 282184 97980
rect 282236 97968 282242 97980
rect 294138 97968 294144 97980
rect 282236 97940 294144 97968
rect 282236 97928 282242 97940
rect 294138 97928 294144 97940
rect 294196 97928 294202 97980
rect 282822 97860 282828 97912
rect 282880 97900 282886 97912
rect 287146 97900 287152 97912
rect 282880 97872 287152 97900
rect 282880 97860 282886 97872
rect 287146 97860 287152 97872
rect 287204 97860 287210 97912
rect 229186 97248 229192 97300
rect 229244 97288 229250 97300
rect 264974 97288 264980 97300
rect 229244 97260 264980 97288
rect 229244 97248 229250 97260
rect 264974 97248 264980 97260
rect 265032 97248 265038 97300
rect 206554 96908 206560 96960
rect 206612 96948 206618 96960
rect 213914 96948 213920 96960
rect 206612 96920 213920 96948
rect 206612 96908 206618 96920
rect 213914 96908 213920 96920
rect 213972 96908 213978 96960
rect 196618 96840 196624 96892
rect 196676 96880 196682 96892
rect 229186 96880 229192 96892
rect 196676 96852 229192 96880
rect 196676 96840 196682 96852
rect 229186 96840 229192 96852
rect 229244 96880 229250 96892
rect 234062 96880 234068 96892
rect 229244 96852 234068 96880
rect 229244 96840 229250 96852
rect 234062 96840 234068 96852
rect 234120 96840 234126 96892
rect 209314 96772 209320 96824
rect 209372 96812 209378 96824
rect 214006 96812 214012 96824
rect 209372 96784 214012 96812
rect 209372 96772 209378 96784
rect 214006 96772 214012 96784
rect 214064 96772 214070 96824
rect 215938 96772 215944 96824
rect 215996 96812 216002 96824
rect 264974 96812 264980 96824
rect 215996 96784 264980 96812
rect 215996 96772 216002 96784
rect 264974 96772 264980 96784
rect 265032 96772 265038 96824
rect 214650 96704 214656 96756
rect 214708 96744 214714 96756
rect 265158 96744 265164 96756
rect 214708 96716 265164 96744
rect 214708 96704 214714 96716
rect 265158 96704 265164 96716
rect 265216 96704 265222 96756
rect 173158 96636 173164 96688
rect 173216 96676 173222 96688
rect 265066 96676 265072 96688
rect 173216 96648 265072 96676
rect 173216 96636 173222 96648
rect 265066 96636 265072 96648
rect 265124 96636 265130 96688
rect 205542 96364 205548 96416
rect 205600 96404 205606 96416
rect 279326 96404 279332 96416
rect 205600 96376 279332 96404
rect 205600 96364 205606 96376
rect 279326 96364 279332 96376
rect 279384 96364 279390 96416
rect 206278 96296 206284 96348
rect 206336 96336 206342 96348
rect 279234 96336 279240 96348
rect 206336 96308 279240 96336
rect 206336 96296 206342 96308
rect 279234 96296 279240 96308
rect 279292 96296 279298 96348
rect 231118 95820 231124 95872
rect 231176 95860 231182 95872
rect 233878 95860 233884 95872
rect 231176 95832 233884 95860
rect 231176 95820 231182 95832
rect 233878 95820 233884 95832
rect 233936 95820 233942 95872
rect 211890 95208 211896 95260
rect 211948 95248 211954 95260
rect 214098 95248 214104 95260
rect 211948 95220 214104 95248
rect 211948 95208 211954 95220
rect 214098 95208 214104 95220
rect 214156 95208 214162 95260
rect 220170 95208 220176 95260
rect 220228 95248 220234 95260
rect 264974 95248 264980 95260
rect 220228 95220 264980 95248
rect 220228 95208 220234 95220
rect 264974 95208 264980 95220
rect 265032 95208 265038 95260
rect 212442 95140 212448 95192
rect 212500 95180 212506 95192
rect 229094 95180 229100 95192
rect 212500 95152 229100 95180
rect 212500 95140 212506 95152
rect 229094 95140 229100 95152
rect 229152 95180 229158 95192
rect 230658 95180 230664 95192
rect 229152 95152 230664 95180
rect 229152 95140 229158 95152
rect 230658 95140 230664 95152
rect 230716 95140 230722 95192
rect 225598 94732 225604 94784
rect 225656 94772 225662 94784
rect 234154 94772 234160 94784
rect 225656 94744 234160 94772
rect 225656 94732 225662 94744
rect 234154 94732 234160 94744
rect 234212 94732 234218 94784
rect 221550 94664 221556 94716
rect 221608 94704 221614 94716
rect 249334 94704 249340 94716
rect 221608 94676 249340 94704
rect 221608 94664 221614 94676
rect 249334 94664 249340 94676
rect 249392 94664 249398 94716
rect 228358 94596 228364 94648
rect 228416 94636 228422 94648
rect 256326 94636 256332 94648
rect 228416 94608 256332 94636
rect 228416 94596 228422 94608
rect 256326 94596 256332 94608
rect 256384 94596 256390 94648
rect 224310 94528 224316 94580
rect 224368 94568 224374 94580
rect 261294 94568 261300 94580
rect 224368 94540 261300 94568
rect 224368 94528 224374 94540
rect 261294 94528 261300 94540
rect 261352 94528 261358 94580
rect 222838 94460 222844 94512
rect 222896 94500 222902 94512
rect 265710 94500 265716 94512
rect 222896 94472 265716 94500
rect 222896 94460 222902 94472
rect 265710 94460 265716 94472
rect 265768 94460 265774 94512
rect 267642 94460 267648 94512
rect 267700 94500 267706 94512
rect 269114 94500 269120 94512
rect 267700 94472 269120 94500
rect 267700 94460 267706 94472
rect 269114 94460 269120 94472
rect 269172 94460 269178 94512
rect 151630 94120 151636 94172
rect 151688 94160 151694 94172
rect 166258 94160 166264 94172
rect 151688 94132 166264 94160
rect 151688 94120 151694 94132
rect 166258 94120 166264 94132
rect 166316 94120 166322 94172
rect 110690 94052 110696 94104
rect 110748 94092 110754 94104
rect 173342 94092 173348 94104
rect 110748 94064 173348 94092
rect 110748 94052 110754 94064
rect 173342 94052 173348 94064
rect 173400 94052 173406 94104
rect 119430 93984 119436 94036
rect 119488 94024 119494 94036
rect 185578 94024 185584 94036
rect 119488 93996 185584 94024
rect 119488 93984 119494 93996
rect 185578 93984 185584 93996
rect 185636 93984 185642 94036
rect 109034 93916 109040 93968
rect 109092 93956 109098 93968
rect 181530 93956 181536 93968
rect 109092 93928 181536 93956
rect 109092 93916 109098 93928
rect 181530 93916 181536 93928
rect 181588 93916 181594 93968
rect 115842 93848 115848 93900
rect 115900 93888 115906 93900
rect 196802 93888 196808 93900
rect 115900 93860 196808 93888
rect 115900 93848 115906 93860
rect 196802 93848 196808 93860
rect 196860 93848 196866 93900
rect 213178 93780 213184 93832
rect 213236 93820 213242 93832
rect 281810 93820 281816 93832
rect 213236 93792 281816 93820
rect 213236 93780 213242 93792
rect 281810 93780 281816 93792
rect 281868 93780 281874 93832
rect 230658 93712 230664 93764
rect 230716 93752 230722 93764
rect 276934 93752 276940 93764
rect 230716 93724 276940 93752
rect 230716 93712 230722 93724
rect 276934 93712 276940 93724
rect 276992 93712 276998 93764
rect 234062 93644 234068 93696
rect 234120 93684 234126 93696
rect 270954 93684 270960 93696
rect 234120 93656 270960 93684
rect 234120 93644 234126 93656
rect 270954 93644 270960 93656
rect 271012 93644 271018 93696
rect 151538 93440 151544 93492
rect 151596 93480 151602 93492
rect 170398 93480 170404 93492
rect 151596 93452 170404 93480
rect 151596 93440 151602 93452
rect 170398 93440 170404 93452
rect 170456 93440 170462 93492
rect 152090 93372 152096 93424
rect 152148 93412 152154 93424
rect 184290 93412 184296 93424
rect 152148 93384 184296 93412
rect 152148 93372 152154 93384
rect 184290 93372 184296 93384
rect 184348 93372 184354 93424
rect 125410 93304 125416 93356
rect 125468 93344 125474 93356
rect 193950 93344 193956 93356
rect 125468 93316 193956 93344
rect 125468 93304 125474 93316
rect 193950 93304 193956 93316
rect 194008 93304 194014 93356
rect 213270 93304 213276 93356
rect 213328 93344 213334 93356
rect 230014 93344 230020 93356
rect 213328 93316 230020 93344
rect 213328 93304 213334 93316
rect 230014 93304 230020 93316
rect 230072 93304 230078 93356
rect 100570 93236 100576 93288
rect 100628 93276 100634 93288
rect 169110 93276 169116 93288
rect 100628 93248 169116 93276
rect 100628 93236 100634 93248
rect 169110 93236 169116 93248
rect 169168 93236 169174 93288
rect 204898 93236 204904 93288
rect 204956 93276 204962 93288
rect 236914 93276 236920 93288
rect 204956 93248 236920 93276
rect 204956 93236 204962 93248
rect 236914 93236 236920 93248
rect 236972 93236 236978 93288
rect 105538 93168 105544 93220
rect 105596 93208 105602 93220
rect 177574 93208 177580 93220
rect 105596 93180 177580 93208
rect 105596 93168 105602 93180
rect 177574 93168 177580 93180
rect 177632 93168 177638 93220
rect 195330 93168 195336 93220
rect 195388 93208 195394 93220
rect 238294 93208 238300 93220
rect 195388 93180 238300 93208
rect 195388 93168 195394 93180
rect 238294 93168 238300 93180
rect 238352 93168 238358 93220
rect 118234 93100 118240 93152
rect 118292 93140 118298 93152
rect 206462 93140 206468 93152
rect 118292 93112 206468 93140
rect 118292 93100 118298 93112
rect 206462 93100 206468 93112
rect 206520 93100 206526 93152
rect 226978 93100 226984 93152
rect 227036 93140 227042 93152
rect 258902 93140 258908 93152
rect 227036 93112 258908 93140
rect 227036 93100 227042 93112
rect 258902 93100 258908 93112
rect 258960 93100 258966 93152
rect 230658 92556 230664 92608
rect 230716 92596 230722 92608
rect 231210 92596 231216 92608
rect 230716 92568 231216 92596
rect 230716 92556 230722 92568
rect 231210 92556 231216 92568
rect 231268 92556 231274 92608
rect 109586 92420 109592 92472
rect 109644 92460 109650 92472
rect 213362 92460 213368 92472
rect 109644 92432 213368 92460
rect 109644 92420 109650 92432
rect 213362 92420 213368 92432
rect 213420 92420 213426 92472
rect 113266 92352 113272 92404
rect 113324 92392 113330 92404
rect 216030 92392 216036 92404
rect 113324 92364 216036 92392
rect 113324 92352 113330 92364
rect 216030 92352 216036 92364
rect 216088 92352 216094 92404
rect 123018 92284 123024 92336
rect 123076 92324 123082 92336
rect 195422 92324 195428 92336
rect 123076 92296 195428 92324
rect 123076 92284 123082 92296
rect 195422 92284 195428 92296
rect 195480 92284 195486 92336
rect 115750 92216 115756 92268
rect 115808 92256 115814 92268
rect 182818 92256 182824 92268
rect 115808 92228 182824 92256
rect 115808 92216 115814 92228
rect 182818 92216 182824 92228
rect 182876 92216 182882 92268
rect 105722 92148 105728 92200
rect 105780 92188 105786 92200
rect 169202 92188 169208 92200
rect 105780 92160 169208 92188
rect 105780 92148 105786 92160
rect 169202 92148 169208 92160
rect 169260 92148 169266 92200
rect 125778 92080 125784 92132
rect 125836 92120 125842 92132
rect 177298 92120 177304 92132
rect 125836 92092 177304 92120
rect 125836 92080 125842 92092
rect 177298 92080 177304 92092
rect 177356 92080 177362 92132
rect 200758 91944 200764 91996
rect 200816 91984 200822 91996
rect 235442 91984 235448 91996
rect 200816 91956 235448 91984
rect 200816 91944 200822 91956
rect 235442 91944 235448 91956
rect 235500 91944 235506 91996
rect 206278 91876 206284 91928
rect 206336 91916 206342 91928
rect 242526 91916 242532 91928
rect 206336 91888 242532 91916
rect 206336 91876 206342 91888
rect 242526 91876 242532 91888
rect 242584 91876 242590 91928
rect 216122 91808 216128 91860
rect 216180 91848 216186 91860
rect 260374 91848 260380 91860
rect 216180 91820 260380 91848
rect 216180 91808 216186 91820
rect 260374 91808 260380 91820
rect 260432 91808 260438 91860
rect 218698 91740 218704 91792
rect 218756 91780 218762 91792
rect 263042 91780 263048 91792
rect 218756 91752 263048 91780
rect 218756 91740 218762 91752
rect 263042 91740 263048 91752
rect 263100 91740 263106 91792
rect 85850 91128 85856 91180
rect 85908 91168 85914 91180
rect 116578 91168 116584 91180
rect 85908 91140 116584 91168
rect 85908 91128 85914 91140
rect 116578 91128 116584 91140
rect 116636 91128 116642 91180
rect 74810 91060 74816 91112
rect 74868 91100 74874 91112
rect 115198 91100 115204 91112
rect 74868 91072 115204 91100
rect 74868 91060 74874 91072
rect 115198 91060 115204 91072
rect 115256 91060 115262 91112
rect 104434 90992 104440 91044
rect 104492 91032 104498 91044
rect 200850 91032 200856 91044
rect 104492 91004 200856 91032
rect 104492 90992 104498 91004
rect 200850 90992 200856 91004
rect 200908 90992 200914 91044
rect 91462 90924 91468 90976
rect 91520 90964 91526 90976
rect 182910 90964 182916 90976
rect 91520 90936 182916 90964
rect 91520 90924 91526 90936
rect 182910 90924 182916 90936
rect 182968 90924 182974 90976
rect 99006 90856 99012 90908
rect 99064 90896 99070 90908
rect 178862 90896 178868 90908
rect 99064 90868 178868 90896
rect 99064 90856 99070 90868
rect 178862 90856 178868 90868
rect 178920 90856 178926 90908
rect 106734 90788 106740 90840
rect 106792 90828 106798 90840
rect 185670 90828 185676 90840
rect 106792 90800 185676 90828
rect 106792 90788 106798 90800
rect 185670 90788 185676 90800
rect 185728 90788 185734 90840
rect 121178 90720 121184 90772
rect 121236 90760 121242 90772
rect 171778 90760 171784 90772
rect 121236 90732 171784 90760
rect 121236 90720 121242 90732
rect 171778 90720 171784 90732
rect 171836 90720 171842 90772
rect 136174 90652 136180 90704
rect 136232 90692 136238 90704
rect 166350 90692 166356 90704
rect 136232 90664 166356 90692
rect 136232 90652 136238 90664
rect 166350 90652 166356 90664
rect 166408 90652 166414 90704
rect 220078 90448 220084 90500
rect 220136 90488 220142 90500
rect 254670 90488 254676 90500
rect 220136 90460 254676 90488
rect 220136 90448 220142 90460
rect 254670 90448 254676 90460
rect 254728 90448 254734 90500
rect 187050 90380 187056 90432
rect 187108 90420 187114 90432
rect 258994 90420 259000 90432
rect 187108 90392 259000 90420
rect 187108 90380 187114 90392
rect 258994 90380 259000 90392
rect 259052 90380 259058 90432
rect 177298 90312 177304 90364
rect 177356 90352 177362 90364
rect 265802 90352 265808 90364
rect 177356 90324 265808 90352
rect 177356 90312 177362 90324
rect 265802 90312 265808 90324
rect 265860 90312 265866 90364
rect 101858 89632 101864 89684
rect 101916 89672 101922 89684
rect 211798 89672 211804 89684
rect 101916 89644 211804 89672
rect 101916 89632 101922 89644
rect 211798 89632 211804 89644
rect 211856 89632 211862 89684
rect 97350 89564 97356 89616
rect 97408 89604 97414 89616
rect 198182 89604 198188 89616
rect 97408 89576 198188 89604
rect 97408 89564 97414 89576
rect 198182 89564 198188 89576
rect 198240 89564 198246 89616
rect 117130 89496 117136 89548
rect 117188 89536 117194 89548
rect 207658 89536 207664 89548
rect 117188 89508 207664 89536
rect 117188 89496 117194 89508
rect 207658 89496 207664 89508
rect 207716 89496 207722 89548
rect 86770 89428 86776 89480
rect 86828 89468 86834 89480
rect 164878 89468 164884 89480
rect 86828 89440 164884 89468
rect 86828 89428 86834 89440
rect 164878 89428 164884 89440
rect 164936 89428 164942 89480
rect 110138 89360 110144 89412
rect 110196 89400 110202 89412
rect 171870 89400 171876 89412
rect 110196 89372 171876 89400
rect 110196 89360 110202 89372
rect 171870 89360 171876 89372
rect 171928 89360 171934 89412
rect 126606 89292 126612 89344
rect 126664 89332 126670 89344
rect 167638 89332 167644 89344
rect 126664 89304 167644 89332
rect 126664 89292 126670 89304
rect 167638 89292 167644 89304
rect 167696 89292 167702 89344
rect 197998 89088 198004 89140
rect 198056 89128 198062 89140
rect 232682 89128 232688 89140
rect 198056 89100 232688 89128
rect 198056 89088 198062 89100
rect 232682 89088 232688 89100
rect 232740 89088 232746 89140
rect 217318 89020 217324 89072
rect 217376 89060 217382 89072
rect 257430 89060 257436 89072
rect 217376 89032 257436 89060
rect 217376 89020 217382 89032
rect 257430 89020 257436 89032
rect 257488 89020 257494 89072
rect 202230 88952 202236 89004
rect 202288 88992 202294 89004
rect 253474 88992 253480 89004
rect 202288 88964 253480 88992
rect 202288 88952 202294 88964
rect 253474 88952 253480 88964
rect 253532 88952 253538 89004
rect 107930 88272 107936 88324
rect 107988 88312 107994 88324
rect 216214 88312 216220 88324
rect 107988 88284 216220 88312
rect 107988 88272 107994 88284
rect 216214 88272 216220 88284
rect 216272 88272 216278 88324
rect 102870 88204 102876 88256
rect 102928 88244 102934 88256
rect 196710 88244 196716 88256
rect 102928 88216 196716 88244
rect 102928 88204 102934 88216
rect 196710 88204 196716 88216
rect 196768 88204 196774 88256
rect 113818 88136 113824 88188
rect 113876 88176 113882 88188
rect 192478 88176 192484 88188
rect 113876 88148 192484 88176
rect 113876 88136 113882 88148
rect 192478 88136 192484 88148
rect 192536 88136 192542 88188
rect 94406 88068 94412 88120
rect 94464 88108 94470 88120
rect 167822 88108 167828 88120
rect 94464 88080 167828 88108
rect 94464 88068 94470 88080
rect 167822 88068 167828 88080
rect 167880 88068 167886 88120
rect 96338 88000 96344 88052
rect 96396 88040 96402 88052
rect 166442 88040 166448 88052
rect 96396 88012 166448 88040
rect 96396 88000 96402 88012
rect 166442 88000 166448 88012
rect 166500 88000 166506 88052
rect 124122 87932 124128 87984
rect 124180 87972 124186 87984
rect 178770 87972 178776 87984
rect 124180 87944 178776 87972
rect 124180 87932 124186 87944
rect 178770 87932 178776 87944
rect 178828 87932 178834 87984
rect 209038 87728 209044 87780
rect 209096 87768 209102 87780
rect 247862 87768 247868 87780
rect 209096 87740 247868 87768
rect 209096 87728 209102 87740
rect 247862 87728 247868 87740
rect 247920 87728 247926 87780
rect 221458 87660 221464 87712
rect 221516 87700 221522 87712
rect 264514 87700 264520 87712
rect 221516 87672 264520 87700
rect 221516 87660 221522 87672
rect 264514 87660 264520 87672
rect 264572 87660 264578 87712
rect 191190 87592 191196 87644
rect 191248 87632 191254 87644
rect 250714 87632 250720 87644
rect 191248 87604 250720 87632
rect 191248 87592 191254 87604
rect 250714 87592 250720 87604
rect 250772 87592 250778 87644
rect 112714 86912 112720 86964
rect 112772 86952 112778 86964
rect 209222 86952 209228 86964
rect 112772 86924 209228 86952
rect 112772 86912 112778 86924
rect 209222 86912 209228 86924
rect 209280 86912 209286 86964
rect 89162 86844 89168 86896
rect 89220 86884 89226 86896
rect 169294 86884 169300 86896
rect 89220 86856 169300 86884
rect 89220 86844 89226 86856
rect 169294 86844 169300 86856
rect 169352 86844 169358 86896
rect 111334 86776 111340 86828
rect 111392 86816 111398 86828
rect 189810 86816 189816 86828
rect 111392 86788 189816 86816
rect 111392 86776 111398 86788
rect 189810 86776 189816 86788
rect 189868 86776 189874 86828
rect 100202 86708 100208 86760
rect 100260 86748 100266 86760
rect 177482 86748 177488 86760
rect 100260 86720 177488 86748
rect 100260 86708 100266 86720
rect 177482 86708 177488 86720
rect 177540 86708 177546 86760
rect 112070 86640 112076 86692
rect 112128 86680 112134 86692
rect 181438 86680 181444 86692
rect 112128 86652 181444 86680
rect 112128 86640 112134 86652
rect 181438 86640 181444 86652
rect 181496 86640 181502 86692
rect 121914 86572 121920 86624
rect 121972 86612 121978 86624
rect 173434 86612 173440 86624
rect 121972 86584 173440 86612
rect 121972 86572 121978 86584
rect 173434 86572 173440 86584
rect 173492 86572 173498 86624
rect 184290 86232 184296 86284
rect 184348 86272 184354 86284
rect 252186 86272 252192 86284
rect 184348 86244 252192 86272
rect 184348 86232 184354 86244
rect 252186 86232 252192 86244
rect 252244 86232 252250 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 18598 85524 18604 85536
rect 3200 85496 18604 85524
rect 3200 85484 3206 85496
rect 18598 85484 18604 85496
rect 18656 85484 18662 85536
rect 93118 85484 93124 85536
rect 93176 85524 93182 85536
rect 199378 85524 199384 85536
rect 93176 85496 199384 85524
rect 93176 85484 93182 85496
rect 199378 85484 199384 85496
rect 199436 85484 199442 85536
rect 97810 85416 97816 85468
rect 97868 85456 97874 85468
rect 202322 85456 202328 85468
rect 97868 85428 202328 85456
rect 97868 85416 97874 85428
rect 202322 85416 202328 85428
rect 202380 85416 202386 85468
rect 119706 85348 119712 85400
rect 119764 85388 119770 85400
rect 203518 85388 203524 85400
rect 119764 85360 203524 85388
rect 119764 85348 119770 85360
rect 203518 85348 203524 85360
rect 203576 85348 203582 85400
rect 88058 85280 88064 85332
rect 88116 85320 88122 85332
rect 166534 85320 166540 85332
rect 88116 85292 166540 85320
rect 88116 85280 88122 85292
rect 166534 85280 166540 85292
rect 166592 85280 166598 85332
rect 115014 85212 115020 85264
rect 115072 85252 115078 85264
rect 193858 85252 193864 85264
rect 115072 85224 193864 85252
rect 115072 85212 115078 85224
rect 193858 85212 193864 85224
rect 193916 85212 193922 85264
rect 98730 85144 98736 85196
rect 98788 85184 98794 85196
rect 174538 85184 174544 85196
rect 98788 85156 174544 85184
rect 98788 85144 98794 85156
rect 174538 85144 174544 85156
rect 174596 85144 174602 85196
rect 211798 84804 211804 84856
rect 211856 84844 211862 84856
rect 261662 84844 261668 84856
rect 211856 84816 261668 84844
rect 211856 84804 211862 84816
rect 261662 84804 261668 84816
rect 261720 84804 261726 84856
rect 102042 84124 102048 84176
rect 102100 84164 102106 84176
rect 210418 84164 210424 84176
rect 102100 84136 210424 84164
rect 102100 84124 102106 84136
rect 210418 84124 210424 84136
rect 210476 84124 210482 84176
rect 95142 84056 95148 84108
rect 95200 84096 95206 84108
rect 191282 84096 191288 84108
rect 95200 84068 191288 84096
rect 95200 84056 95206 84068
rect 191282 84056 191288 84068
rect 191340 84056 191346 84108
rect 114462 83988 114468 84040
rect 114520 84028 114526 84040
rect 209130 84028 209136 84040
rect 114520 84000 209136 84028
rect 114520 83988 114526 84000
rect 209130 83988 209136 84000
rect 209188 83988 209194 84040
rect 101950 83920 101956 83972
rect 102008 83960 102014 83972
rect 170490 83960 170496 83972
rect 102008 83932 170496 83960
rect 102008 83920 102014 83932
rect 170490 83920 170496 83932
rect 170548 83920 170554 83972
rect 132402 83852 132408 83904
rect 132460 83892 132466 83904
rect 184198 83892 184204 83904
rect 132460 83864 184204 83892
rect 132460 83852 132466 83864
rect 184198 83852 184204 83864
rect 184256 83852 184262 83904
rect 37182 83444 37188 83496
rect 37240 83484 37246 83496
rect 246482 83484 246488 83496
rect 37240 83456 246488 83484
rect 37240 83444 37246 83456
rect 246482 83444 246488 83456
rect 246540 83444 246546 83496
rect 67634 82764 67640 82816
rect 67692 82804 67698 82816
rect 209314 82804 209320 82816
rect 67692 82776 209320 82804
rect 67692 82764 67698 82776
rect 209314 82764 209320 82776
rect 209372 82764 209378 82816
rect 99098 82696 99104 82748
rect 99156 82736 99162 82748
rect 204990 82736 204996 82748
rect 99156 82708 204996 82736
rect 99156 82696 99162 82708
rect 204990 82696 204996 82708
rect 205048 82696 205054 82748
rect 122742 82628 122748 82680
rect 122800 82668 122806 82680
rect 206370 82668 206376 82680
rect 122800 82640 206376 82668
rect 122800 82628 122806 82640
rect 206370 82628 206376 82640
rect 206428 82628 206434 82680
rect 121270 82560 121276 82612
rect 121328 82600 121334 82612
rect 187142 82600 187148 82612
rect 121328 82572 187148 82600
rect 121328 82560 121334 82572
rect 187142 82560 187148 82572
rect 187200 82560 187206 82612
rect 151722 82492 151728 82544
rect 151780 82532 151786 82544
rect 180058 82532 180064 82544
rect 151780 82504 180064 82532
rect 151780 82492 151786 82504
rect 180058 82492 180064 82504
rect 180116 82492 180122 82544
rect 106182 82084 106188 82136
rect 106240 82124 106246 82136
rect 229830 82124 229836 82136
rect 106240 82096 229836 82124
rect 106240 82084 106246 82096
rect 229830 82084 229836 82096
rect 229888 82084 229894 82136
rect 63402 81336 63408 81388
rect 63460 81376 63466 81388
rect 195514 81376 195520 81388
rect 63460 81348 195520 81376
rect 63460 81336 63466 81348
rect 195514 81336 195520 81348
rect 195572 81336 195578 81388
rect 129642 81268 129648 81320
rect 129700 81308 129706 81320
rect 198090 81308 198096 81320
rect 129700 81280 198096 81308
rect 129700 81268 129706 81280
rect 198090 81268 198096 81280
rect 198148 81268 198154 81320
rect 108942 81200 108948 81252
rect 109000 81240 109006 81252
rect 175918 81240 175924 81252
rect 109000 81212 175924 81240
rect 109000 81200 109006 81212
rect 175918 81200 175924 81212
rect 175976 81200 175982 81252
rect 113082 80724 113088 80776
rect 113140 80764 113146 80776
rect 239582 80764 239588 80776
rect 113140 80736 239588 80764
rect 113140 80724 113146 80736
rect 239582 80724 239588 80736
rect 239640 80724 239646 80776
rect 79318 80656 79324 80708
rect 79376 80696 79382 80708
rect 265618 80696 265624 80708
rect 79376 80668 265624 80696
rect 79376 80656 79382 80668
rect 265618 80656 265624 80668
rect 265676 80656 265682 80708
rect 66162 79976 66168 80028
rect 66220 80016 66226 80028
rect 170582 80016 170588 80028
rect 66220 79988 170588 80016
rect 66220 79976 66226 79988
rect 170582 79976 170588 79988
rect 170640 79976 170646 80028
rect 128262 79908 128268 79960
rect 128320 79948 128326 79960
rect 188338 79948 188344 79960
rect 128320 79920 188344 79948
rect 128320 79908 128326 79920
rect 188338 79908 188344 79920
rect 188396 79908 188402 79960
rect 124122 79432 124128 79484
rect 124180 79472 124186 79484
rect 254762 79472 254768 79484
rect 124180 79444 254768 79472
rect 124180 79432 124186 79444
rect 254762 79432 254768 79444
rect 254820 79432 254826 79484
rect 108942 79364 108948 79416
rect 109000 79404 109006 79416
rect 256142 79404 256148 79416
rect 109000 79376 256148 79404
rect 109000 79364 109006 79376
rect 256142 79364 256148 79376
rect 256200 79364 256206 79416
rect 71038 79296 71044 79348
rect 71096 79336 71102 79348
rect 221550 79336 221556 79348
rect 71096 79308 221556 79336
rect 71096 79296 71102 79308
rect 221550 79296 221556 79308
rect 221608 79296 221614 79348
rect 67542 78616 67548 78668
rect 67600 78656 67606 78668
rect 213454 78656 213460 78668
rect 67600 78628 213460 78656
rect 67600 78616 67606 78628
rect 213454 78616 213460 78628
rect 213512 78616 213518 78668
rect 135162 78548 135168 78600
rect 135220 78588 135226 78600
rect 202138 78588 202144 78600
rect 135220 78560 202144 78588
rect 135220 78548 135226 78560
rect 202138 78548 202144 78560
rect 202196 78548 202202 78600
rect 126882 78480 126888 78532
rect 126940 78520 126946 78532
rect 186958 78520 186964 78532
rect 126940 78492 186964 78520
rect 126940 78480 126946 78492
rect 186958 78480 186964 78492
rect 187016 78480 187022 78532
rect 102042 78004 102048 78056
rect 102100 78044 102106 78056
rect 253290 78044 253296 78056
rect 102100 78016 253296 78044
rect 102100 78004 102106 78016
rect 253290 78004 253296 78016
rect 253348 78004 253354 78056
rect 50982 77936 50988 77988
rect 51040 77976 51046 77988
rect 267182 77976 267188 77988
rect 51040 77948 267188 77976
rect 51040 77936 51046 77948
rect 267182 77936 267188 77948
rect 267240 77936 267246 77988
rect 107562 77188 107568 77240
rect 107620 77228 107626 77240
rect 173250 77228 173256 77240
rect 107620 77200 173256 77228
rect 107620 77188 107626 77200
rect 173250 77188 173256 77200
rect 173308 77188 173314 77240
rect 131022 77120 131028 77172
rect 131080 77160 131086 77172
rect 191098 77160 191104 77172
rect 131080 77132 191104 77160
rect 131080 77120 131086 77132
rect 191098 77120 191104 77132
rect 191156 77120 191162 77172
rect 125502 76644 125508 76696
rect 125560 76684 125566 76696
rect 243538 76684 243544 76696
rect 125560 76656 243544 76684
rect 125560 76644 125566 76656
rect 243538 76644 243544 76656
rect 243596 76644 243602 76696
rect 73062 76576 73068 76628
rect 73120 76616 73126 76628
rect 264422 76616 264428 76628
rect 73120 76588 264428 76616
rect 73120 76576 73126 76588
rect 264422 76576 264428 76588
rect 264480 76576 264486 76628
rect 30282 76508 30288 76560
rect 30340 76548 30346 76560
rect 249242 76548 249248 76560
rect 30340 76520 249248 76548
rect 30340 76508 30346 76520
rect 249242 76508 249248 76520
rect 249300 76508 249306 76560
rect 115198 75828 115204 75880
rect 115256 75868 115262 75880
rect 211890 75868 211896 75880
rect 115256 75840 211896 75868
rect 115256 75828 115262 75840
rect 211890 75828 211896 75840
rect 211948 75828 211954 75880
rect 133782 75760 133788 75812
rect 133840 75800 133846 75812
rect 195238 75800 195244 75812
rect 133840 75772 195244 75800
rect 133840 75760 133846 75772
rect 195238 75760 195244 75772
rect 195296 75760 195302 75812
rect 91002 75216 91008 75268
rect 91060 75256 91066 75268
rect 241146 75256 241152 75268
rect 91060 75228 241152 75256
rect 91060 75216 91066 75228
rect 241146 75216 241152 75228
rect 241204 75216 241210 75268
rect 34422 75148 34428 75200
rect 34480 75188 34486 75200
rect 262950 75188 262956 75200
rect 34480 75160 262956 75188
rect 34480 75148 34486 75160
rect 262950 75148 262956 75160
rect 263008 75148 263014 75200
rect 116578 74468 116584 74520
rect 116636 74508 116642 74520
rect 203610 74508 203616 74520
rect 116636 74480 203616 74508
rect 116636 74468 116642 74480
rect 203610 74468 203616 74480
rect 203668 74468 203674 74520
rect 95142 73992 95148 74044
rect 95200 74032 95206 74044
rect 243722 74032 243728 74044
rect 95200 74004 243728 74032
rect 95200 73992 95206 74004
rect 243722 73992 243728 74004
rect 243780 73992 243786 74044
rect 75822 73924 75828 73976
rect 75880 73964 75886 73976
rect 239490 73964 239496 73976
rect 75880 73936 239496 73964
rect 75880 73924 75886 73936
rect 239490 73924 239496 73936
rect 239548 73924 239554 73976
rect 41322 73856 41328 73908
rect 41380 73896 41386 73908
rect 242434 73896 242440 73908
rect 41380 73868 242440 73896
rect 41380 73856 41386 73868
rect 242434 73856 242440 73868
rect 242492 73856 242498 73908
rect 15102 73788 15108 73840
rect 15160 73828 15166 73840
rect 261570 73828 261576 73840
rect 15160 73800 261576 73828
rect 15160 73788 15166 73800
rect 261570 73788 261576 73800
rect 261628 73788 261634 73840
rect 574738 73108 574744 73160
rect 574796 73148 574802 73160
rect 580166 73148 580172 73160
rect 574796 73120 580172 73148
rect 574796 73108 574802 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 115842 72564 115848 72616
rect 115900 72604 115906 72616
rect 236730 72604 236736 72616
rect 115900 72576 236736 72604
rect 115900 72564 115906 72576
rect 236730 72564 236736 72576
rect 236788 72564 236794 72616
rect 89622 72496 89628 72548
rect 89680 72536 89686 72548
rect 245010 72536 245016 72548
rect 89680 72508 245016 72536
rect 89680 72496 89686 72508
rect 245010 72496 245016 72508
rect 245068 72496 245074 72548
rect 70302 72428 70308 72480
rect 70360 72468 70366 72480
rect 258810 72468 258816 72480
rect 70360 72440 258816 72468
rect 70360 72428 70366 72440
rect 258810 72428 258816 72440
rect 258868 72428 258874 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 57238 71720 57244 71732
rect 3476 71692 57244 71720
rect 3476 71680 3482 71692
rect 57238 71680 57244 71692
rect 57296 71680 57302 71732
rect 65978 71680 65984 71732
rect 66036 71720 66042 71732
rect 206554 71720 206560 71732
rect 66036 71692 206560 71720
rect 66036 71680 66042 71692
rect 206554 71680 206560 71692
rect 206612 71680 206618 71732
rect 122742 71068 122748 71120
rect 122800 71108 122806 71120
rect 251818 71108 251824 71120
rect 122800 71080 251824 71108
rect 122800 71068 122806 71080
rect 251818 71068 251824 71080
rect 251876 71068 251882 71120
rect 86862 71000 86868 71052
rect 86920 71040 86926 71052
rect 264330 71040 264336 71052
rect 86920 71012 264336 71040
rect 86920 71000 86926 71012
rect 264330 71000 264336 71012
rect 264388 71000 264394 71052
rect 107562 69776 107568 69828
rect 107620 69816 107626 69828
rect 233970 69816 233976 69828
rect 107620 69788 233976 69816
rect 107620 69776 107626 69788
rect 233970 69776 233976 69788
rect 234028 69776 234034 69828
rect 111702 69708 111708 69760
rect 111760 69748 111766 69760
rect 239398 69748 239404 69760
rect 111760 69720 239404 69748
rect 111760 69708 111766 69720
rect 239398 69708 239404 69720
rect 239456 69708 239462 69760
rect 68922 69640 68928 69692
rect 68980 69680 68986 69692
rect 260190 69680 260196 69692
rect 68980 69652 260196 69680
rect 68980 69640 68986 69652
rect 260190 69640 260196 69652
rect 260248 69640 260254 69692
rect 117222 68348 117228 68400
rect 117280 68388 117286 68400
rect 235258 68388 235264 68400
rect 117280 68360 235264 68388
rect 117280 68348 117286 68360
rect 235258 68348 235264 68360
rect 235316 68348 235322 68400
rect 88242 68280 88248 68332
rect 88300 68320 88306 68332
rect 243630 68320 243636 68332
rect 88300 68292 243636 68320
rect 88300 68280 88306 68292
rect 243630 68280 243636 68292
rect 243688 68280 243694 68332
rect 77202 66852 77208 66904
rect 77260 66892 77266 66904
rect 242342 66892 242348 66904
rect 77260 66864 242348 66892
rect 77260 66852 77266 66864
rect 242342 66852 242348 66864
rect 242400 66852 242406 66904
rect 84102 65492 84108 65544
rect 84160 65532 84166 65544
rect 246574 65532 246580 65544
rect 84160 65504 246580 65532
rect 84160 65492 84166 65504
rect 246574 65492 246580 65504
rect 246632 65492 246638 65544
rect 47578 64200 47584 64252
rect 47636 64240 47642 64252
rect 222930 64240 222936 64252
rect 47636 64212 222936 64240
rect 47636 64200 47642 64212
rect 222930 64200 222936 64212
rect 222988 64200 222994 64252
rect 35802 64132 35808 64184
rect 35860 64172 35866 64184
rect 249150 64172 249156 64184
rect 35860 64144 249156 64172
rect 35860 64132 35866 64144
rect 249150 64132 249156 64144
rect 249208 64132 249214 64184
rect 97902 62840 97908 62892
rect 97960 62880 97966 62892
rect 260282 62880 260288 62892
rect 97960 62852 260288 62880
rect 97960 62840 97966 62852
rect 260282 62840 260288 62852
rect 260340 62840 260346 62892
rect 53742 62772 53748 62824
rect 53800 62812 53806 62824
rect 267090 62812 267096 62824
rect 53800 62784 267096 62812
rect 53800 62772 53806 62784
rect 267090 62772 267096 62784
rect 267148 62772 267154 62824
rect 93762 61344 93768 61396
rect 93820 61384 93826 61396
rect 229738 61384 229744 61396
rect 93820 61356 229744 61384
rect 93820 61344 93826 61356
rect 229738 61344 229744 61356
rect 229796 61344 229802 61396
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 17218 59344 17224 59356
rect 3108 59316 17224 59344
rect 3108 59304 3114 59316
rect 17218 59304 17224 59316
rect 17276 59304 17282 59356
rect 119890 58692 119896 58744
rect 119948 58732 119954 58744
rect 226978 58732 226984 58744
rect 119948 58704 226984 58732
rect 119948 58692 119954 58704
rect 226978 58692 226984 58704
rect 227036 58692 227042 58744
rect 86770 58624 86776 58676
rect 86828 58664 86834 58676
rect 221458 58664 221464 58676
rect 86828 58636 221464 58664
rect 86828 58624 86834 58636
rect 221458 58624 221464 58636
rect 221516 58624 221522 58676
rect 17862 57196 17868 57248
rect 17920 57236 17926 57248
rect 250530 57236 250536 57248
rect 17920 57208 250536 57236
rect 17920 57196 17926 57208
rect 250530 57196 250536 57208
rect 250588 57196 250594 57248
rect 111610 55904 111616 55956
rect 111668 55944 111674 55956
rect 216122 55944 216128 55956
rect 111668 55916 216128 55944
rect 111668 55904 111674 55916
rect 216122 55904 216128 55916
rect 216180 55904 216186 55956
rect 44082 55836 44088 55888
rect 44140 55876 44146 55888
rect 254578 55876 254584 55888
rect 44140 55848 254584 55876
rect 44140 55836 44146 55848
rect 254578 55836 254584 55848
rect 254636 55836 254642 55888
rect 39942 54476 39948 54528
rect 40000 54516 40006 54528
rect 257338 54516 257344 54528
rect 40000 54488 257344 54516
rect 40000 54476 40006 54488
rect 257338 54476 257344 54488
rect 257396 54476 257402 54528
rect 27522 53116 27528 53168
rect 27580 53156 27586 53168
rect 224310 53156 224316 53168
rect 27580 53128 224316 53156
rect 27580 53116 27586 53128
rect 224310 53116 224316 53128
rect 224368 53116 224374 53168
rect 26142 53048 26148 53100
rect 26200 53088 26206 53100
rect 245102 53088 245108 53100
rect 26200 53060 245108 53088
rect 26200 53048 26206 53060
rect 245102 53048 245108 53060
rect 245160 53048 245166 53100
rect 55122 51756 55128 51808
rect 55180 51796 55186 51808
rect 256050 51796 256056 51808
rect 55180 51768 256056 51796
rect 55180 51756 55186 51768
rect 256050 51756 256056 51768
rect 256108 51756 256114 51808
rect 5442 51688 5448 51740
rect 5500 51728 5506 51740
rect 220170 51728 220176 51740
rect 5500 51700 220176 51728
rect 5500 51688 5506 51700
rect 220170 51688 220176 51700
rect 220228 51688 220234 51740
rect 104158 50328 104164 50380
rect 104216 50368 104222 50380
rect 206278 50368 206284 50380
rect 104216 50340 206284 50368
rect 104216 50328 104222 50340
rect 206278 50328 206284 50340
rect 206336 50328 206342 50380
rect 3418 48968 3424 49020
rect 3476 49008 3482 49020
rect 54478 49008 54484 49020
rect 3476 48980 54484 49008
rect 3476 48968 3482 48980
rect 54478 48968 54484 48980
rect 54536 48968 54542 49020
rect 65518 48968 65524 49020
rect 65576 49008 65582 49020
rect 231118 49008 231124 49020
rect 65576 48980 231124 49008
rect 65576 48968 65582 48980
rect 231118 48968 231124 48980
rect 231176 48968 231182 49020
rect 58618 47608 58624 47660
rect 58676 47648 58682 47660
rect 231210 47648 231216 47660
rect 58676 47620 231216 47648
rect 58676 47608 58682 47620
rect 231210 47608 231216 47620
rect 231268 47608 231274 47660
rect 13722 47540 13728 47592
rect 13780 47580 13786 47592
rect 269114 47580 269120 47592
rect 13780 47552 269120 47580
rect 13780 47540 13786 47552
rect 269114 47540 269120 47552
rect 269172 47540 269178 47592
rect 70210 46180 70216 46232
rect 70268 46220 70274 46232
rect 218698 46220 218704 46232
rect 70268 46192 218704 46220
rect 70268 46180 70274 46192
rect 218698 46180 218704 46192
rect 218756 46180 218762 46232
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4798 45540 4804 45552
rect 2832 45512 4804 45540
rect 2832 45500 2838 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 92382 44888 92388 44940
rect 92440 44928 92446 44940
rect 228358 44928 228364 44940
rect 92440 44900 228364 44928
rect 92440 44888 92446 44900
rect 228358 44888 228364 44900
rect 228416 44888 228422 44940
rect 71682 44820 71688 44872
rect 71740 44860 71746 44872
rect 225598 44860 225604 44872
rect 71740 44832 225604 44860
rect 71740 44820 71746 44832
rect 225598 44820 225604 44832
rect 225656 44820 225662 44872
rect 42702 43392 42708 43444
rect 42760 43432 42766 43444
rect 200758 43432 200764 43444
rect 42760 43404 200764 43432
rect 42760 43392 42766 43404
rect 200758 43392 200764 43404
rect 200816 43392 200822 43444
rect 110322 42100 110328 42152
rect 110380 42140 110386 42152
rect 184290 42140 184296 42152
rect 110380 42112 184296 42140
rect 110380 42100 110386 42112
rect 184290 42100 184296 42112
rect 184348 42100 184354 42152
rect 38562 42032 38568 42084
rect 38620 42072 38626 42084
rect 258718 42072 258724 42084
rect 38620 42044 258724 42072
rect 38620 42032 38626 42044
rect 258718 42032 258724 42044
rect 258776 42032 258782 42084
rect 99282 40672 99288 40724
rect 99340 40712 99346 40724
rect 191190 40712 191196 40724
rect 99340 40684 191196 40712
rect 99340 40672 99346 40684
rect 191190 40672 191196 40684
rect 191248 40672 191254 40724
rect 12342 39312 12348 39364
rect 12400 39352 12406 39364
rect 214650 39352 214656 39364
rect 12400 39324 214656 39352
rect 12400 39312 12406 39324
rect 214650 39312 214656 39324
rect 214708 39312 214714 39364
rect 103422 37952 103428 38004
rect 103480 37992 103486 38004
rect 240778 37992 240784 38004
rect 103480 37964 240784 37992
rect 103480 37952 103486 37964
rect 240778 37952 240784 37964
rect 240836 37952 240842 38004
rect 45462 37884 45468 37936
rect 45520 37924 45526 37936
rect 202230 37924 202236 37936
rect 45520 37896 202236 37924
rect 45520 37884 45526 37896
rect 202230 37884 202236 37896
rect 202288 37884 202294 37936
rect 100662 36524 100668 36576
rect 100720 36564 100726 36576
rect 236638 36564 236644 36576
rect 100720 36536 236644 36564
rect 100720 36524 100726 36536
rect 236638 36524 236644 36536
rect 236696 36524 236702 36576
rect 82722 35232 82728 35284
rect 82780 35272 82786 35284
rect 238110 35272 238116 35284
rect 82780 35244 238116 35272
rect 82780 35232 82786 35244
rect 238110 35232 238116 35244
rect 238168 35232 238174 35284
rect 10962 35164 10968 35216
rect 11020 35204 11026 35216
rect 204898 35204 204904 35216
rect 11020 35176 204904 35204
rect 11020 35164 11026 35176
rect 204898 35164 204904 35176
rect 204956 35164 204962 35216
rect 78582 33736 78588 33788
rect 78640 33776 78646 33788
rect 247678 33776 247684 33788
rect 78640 33748 247684 33776
rect 78640 33736 78646 33748
rect 247678 33736 247684 33748
rect 247736 33736 247742 33788
rect 96522 32444 96528 32496
rect 96580 32484 96586 32496
rect 217318 32484 217324 32496
rect 96580 32456 217324 32484
rect 96580 32444 96586 32456
rect 217318 32444 217324 32456
rect 217376 32444 217382 32496
rect 62022 32376 62028 32428
rect 62080 32416 62086 32428
rect 187050 32416 187056 32428
rect 62080 32388 187056 32416
rect 62080 32376 62086 32388
rect 187050 32376 187056 32388
rect 187108 32376 187114 32428
rect 114462 29656 114468 29708
rect 114520 29696 114526 29708
rect 213270 29696 213276 29708
rect 114520 29668 213276 29696
rect 114520 29656 114526 29668
rect 213270 29656 213276 29668
rect 213328 29656 213334 29708
rect 4062 29588 4068 29640
rect 4120 29628 4126 29640
rect 224218 29628 224224 29640
rect 4120 29600 224224 29628
rect 4120 29588 4126 29600
rect 224218 29588 224224 29600
rect 224276 29588 224282 29640
rect 81342 28296 81348 28348
rect 81400 28336 81406 28348
rect 195330 28336 195336 28348
rect 81400 28308 195336 28336
rect 81400 28296 81406 28308
rect 195330 28296 195336 28308
rect 195388 28296 195394 28348
rect 24762 28228 24768 28280
rect 24820 28268 24826 28280
rect 270586 28268 270592 28280
rect 24820 28240 270592 28268
rect 24820 28228 24826 28240
rect 270586 28228 270592 28240
rect 270644 28228 270650 28280
rect 118602 26936 118608 26988
rect 118660 26976 118666 26988
rect 220078 26976 220084 26988
rect 118660 26948 220084 26976
rect 118660 26936 118666 26948
rect 220078 26936 220084 26948
rect 220136 26936 220142 26988
rect 53650 26868 53656 26920
rect 53708 26908 53714 26920
rect 261478 26908 261484 26920
rect 53708 26880 261484 26908
rect 53708 26868 53714 26880
rect 261478 26868 261484 26880
rect 261536 26868 261542 26920
rect 3970 25508 3976 25560
rect 4028 25548 4034 25560
rect 215938 25548 215944 25560
rect 4028 25520 215944 25548
rect 4028 25508 4034 25520
rect 215938 25508 215944 25520
rect 215996 25508 216002 25560
rect 46842 24080 46848 24132
rect 46900 24120 46906 24132
rect 211798 24120 211804 24132
rect 46900 24092 211804 24120
rect 46900 24080 46906 24092
rect 211798 24080 211804 24092
rect 211856 24080 211862 24132
rect 37090 22720 37096 22772
rect 37148 22760 37154 22772
rect 255958 22760 255964 22772
rect 37148 22732 255964 22760
rect 37148 22720 37154 22732
rect 255958 22720 255964 22732
rect 256016 22720 256022 22772
rect 56502 21360 56508 21412
rect 56560 21400 56566 21412
rect 266998 21400 267004 21412
rect 56560 21372 267004 21400
rect 56560 21360 56566 21372
rect 266998 21360 267004 21372
rect 267056 21360 267062 21412
rect 106 19932 112 19984
rect 164 19972 170 19984
rect 196618 19972 196624 19984
rect 164 19944 196624 19972
rect 164 19932 170 19944
rect 196618 19932 196624 19944
rect 196676 19932 196682 19984
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 244918 18612 244924 18624
rect 9640 18584 244924 18612
rect 9640 18572 9646 18584
rect 244918 18572 244924 18584
rect 244976 18572 244982 18624
rect 49602 17212 49608 17264
rect 49660 17252 49666 17264
rect 260098 17252 260104 17264
rect 49660 17224 260104 17252
rect 49660 17212 49666 17224
rect 260098 17212 260104 17224
rect 260156 17212 260162 17264
rect 66162 15852 66168 15904
rect 66220 15892 66226 15904
rect 250438 15892 250444 15904
rect 66220 15864 250444 15892
rect 66220 15852 66226 15864
rect 250438 15852 250444 15864
rect 250496 15852 250502 15904
rect 59262 14424 59268 14476
rect 59320 14464 59326 14476
rect 253198 14464 253204 14476
rect 59320 14436 253204 14464
rect 59320 14424 59326 14436
rect 253198 14424 253204 14436
rect 253256 14424 253262 14476
rect 60642 13064 60648 13116
rect 60700 13104 60706 13116
rect 209038 13104 209044 13116
rect 60700 13076 209044 13104
rect 60700 13064 60706 13076
rect 209038 13064 209044 13076
rect 209096 13064 209102 13116
rect 85482 11772 85488 11824
rect 85540 11812 85546 11824
rect 246298 11812 246304 11824
rect 85540 11784 246304 11812
rect 85540 11772 85546 11784
rect 246298 11772 246304 11784
rect 246356 11772 246362 11824
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4062 11744 4068 11756
rect 3936 11716 4068 11744
rect 3936 11704 3942 11716
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 47854 11704 47860 11756
rect 47912 11744 47918 11756
rect 262858 11744 262864 11756
rect 47912 11716 262864 11744
rect 47912 11704 47918 11716
rect 262858 11704 262864 11716
rect 262916 11704 262922 11756
rect 79686 10276 79692 10328
rect 79744 10316 79750 10328
rect 249058 10316 249064 10328
rect 79744 10288 249064 10316
rect 79744 10276 79750 10288
rect 249058 10276 249064 10288
rect 249116 10276 249122 10328
rect 104526 8916 104532 8968
rect 104584 8956 104590 8968
rect 238018 8956 238024 8968
rect 104584 8928 238024 8956
rect 104584 8916 104590 8928
rect 238018 8916 238024 8928
rect 238076 8916 238082 8968
rect 44266 7624 44272 7676
rect 44324 7664 44330 7676
rect 240870 7664 240876 7676
rect 44324 7636 240876 7664
rect 44324 7624 44330 7636
rect 240870 7624 240876 7636
rect 240928 7624 240934 7676
rect 12250 7556 12256 7608
rect 12308 7596 12314 7608
rect 242158 7596 242164 7608
rect 12308 7568 242164 7596
rect 12308 7556 12314 7568
rect 242158 7556 242164 7568
rect 242216 7556 242222 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 51718 6848 51724 6860
rect 3476 6820 51724 6848
rect 3476 6808 3482 6820
rect 51718 6808 51724 6820
rect 51776 6808 51782 6860
rect 102226 6196 102232 6248
rect 102284 6236 102290 6248
rect 197998 6236 198004 6248
rect 102284 6208 198004 6236
rect 102284 6196 102290 6208
rect 197998 6196 198004 6208
rect 198056 6196 198062 6248
rect 60826 6128 60832 6180
rect 60884 6168 60890 6180
rect 214558 6168 214564 6180
rect 60884 6140 214564 6168
rect 60884 6128 60890 6140
rect 214558 6128 214564 6140
rect 214616 6128 214622 6180
rect 73798 4836 73804 4888
rect 73856 4876 73862 4888
rect 232498 4876 232504 4888
rect 73856 4848 232504 4876
rect 73856 4836 73862 4848
rect 232498 4836 232504 4848
rect 232556 4836 232562 4888
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 173158 4808 173164 4820
rect 6512 4780 173164 4808
rect 6512 4768 6518 4780
rect 173158 4768 173164 4780
rect 173216 4768 173222 4820
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 71038 3720 71044 3732
rect 51408 3692 71044 3720
rect 51408 3680 51414 3692
rect 71038 3680 71044 3692
rect 71096 3680 71102 3732
rect 35986 3612 35992 3664
rect 36044 3652 36050 3664
rect 37090 3652 37096 3664
rect 36044 3624 37096 3652
rect 36044 3612 36050 3624
rect 37090 3612 37096 3624
rect 37148 3612 37154 3664
rect 58618 3652 58624 3664
rect 55876 3624 58624 3652
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12342 3584 12348 3596
rect 11204 3556 12348 3584
rect 11204 3544 11210 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 47578 3584 47584 3596
rect 19484 3556 47584 3584
rect 19484 3544 19490 3556
rect 47578 3544 47584 3556
rect 47636 3544 47642 3596
rect 48958 3544 48964 3596
rect 49016 3584 49022 3596
rect 49602 3584 49608 3596
rect 49016 3556 49608 3584
rect 49016 3544 49022 3556
rect 49602 3544 49608 3556
rect 49660 3544 49666 3596
rect 50154 3544 50160 3596
rect 50212 3584 50218 3596
rect 50982 3584 50988 3596
rect 50212 3556 50988 3584
rect 50212 3544 50218 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53650 3584 53656 3596
rect 52604 3556 53656 3584
rect 52604 3544 52610 3556
rect 53650 3544 53656 3556
rect 53708 3544 53714 3596
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3878 3516 3884 3528
rect 2924 3488 3884 3516
rect 2924 3476 2930 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 55876 3516 55904 3624
rect 58618 3612 58624 3624
rect 58676 3612 58682 3664
rect 85666 3612 85672 3664
rect 85724 3652 85730 3664
rect 86770 3652 86776 3664
rect 85724 3624 86776 3652
rect 85724 3612 85730 3624
rect 86770 3612 86776 3624
rect 86828 3612 86834 3664
rect 79318 3584 79324 3596
rect 64846 3556 79324 3584
rect 6886 3488 55904 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 6886 3448 6914 3488
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64846 3516 64874 3556
rect 79318 3544 79324 3556
rect 79376 3544 79382 3596
rect 104158 3584 104164 3596
rect 79428 3556 104164 3584
rect 64380 3488 64874 3516
rect 64380 3476 64386 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 77386 3476 77392 3528
rect 77444 3516 77450 3528
rect 79428 3516 79456 3556
rect 104158 3544 104164 3556
rect 104216 3544 104222 3596
rect 105722 3544 105728 3596
rect 105780 3584 105786 3596
rect 106182 3584 106188 3596
rect 105780 3556 106188 3584
rect 105780 3544 105786 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 106918 3544 106924 3596
rect 106976 3584 106982 3596
rect 107562 3584 107568 3596
rect 106976 3556 107568 3584
rect 106976 3544 106982 3556
rect 107562 3544 107568 3556
rect 107620 3544 107626 3596
rect 108114 3544 108120 3596
rect 108172 3584 108178 3596
rect 108942 3584 108948 3596
rect 108172 3556 108948 3584
rect 108172 3544 108178 3556
rect 108942 3544 108948 3556
rect 109000 3544 109006 3596
rect 109310 3544 109316 3596
rect 109368 3584 109374 3596
rect 110322 3584 110328 3596
rect 109368 3556 110328 3584
rect 109368 3544 109374 3556
rect 110322 3544 110328 3556
rect 110380 3544 110386 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 114462 3584 114468 3596
rect 114060 3556 114468 3584
rect 114060 3544 114066 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 115842 3584 115848 3596
rect 115256 3556 115848 3584
rect 115256 3544 115262 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 117222 3584 117228 3596
rect 116452 3556 117228 3584
rect 116452 3544 116458 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 117590 3544 117596 3596
rect 117648 3584 117654 3596
rect 118602 3584 118608 3596
rect 117648 3556 118608 3584
rect 117648 3544 117654 3556
rect 118602 3544 118608 3556
rect 118660 3544 118666 3596
rect 118786 3544 118792 3596
rect 118844 3584 118850 3596
rect 119798 3584 119804 3596
rect 118844 3556 119804 3584
rect 118844 3544 118850 3556
rect 119798 3544 119804 3556
rect 119856 3544 119862 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 122742 3584 122748 3596
rect 122340 3556 122748 3584
rect 122340 3544 122346 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 124122 3584 124128 3596
rect 123536 3556 124128 3584
rect 123536 3544 123542 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 124674 3544 124680 3596
rect 124732 3584 124738 3596
rect 125502 3584 125508 3596
rect 124732 3556 125508 3584
rect 124732 3544 124738 3556
rect 125502 3544 125508 3556
rect 125560 3544 125566 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 178678 3584 178684 3596
rect 125928 3556 178684 3584
rect 125928 3544 125934 3556
rect 178678 3544 178684 3556
rect 178736 3544 178742 3596
rect 77444 3488 79456 3516
rect 77444 3476 77450 3488
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95142 3516 95148 3528
rect 94004 3488 95148 3516
rect 94004 3476 94010 3488
rect 95142 3476 95148 3488
rect 95200 3476 95206 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 222838 3516 222844 3528
rect 100864 3488 222844 3516
rect 1728 3420 6914 3448
rect 1728 3408 1734 3420
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 9582 3448 9588 3460
rect 8812 3420 9588 3448
rect 8812 3408 8818 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 10962 3448 10968 3460
rect 10008 3420 10968 3448
rect 10008 3408 10014 3420
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16482 3448 16488 3460
rect 15988 3420 16488 3448
rect 15988 3408 15994 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17862 3448 17868 3460
rect 17092 3420 17868 3448
rect 17092 3408 17098 3420
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 19242 3448 19248 3460
rect 18288 3420 19248 3448
rect 18288 3408 18294 3420
rect 19242 3408 19248 3420
rect 19300 3408 19306 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 24762 3448 24768 3460
rect 24268 3420 24768 3448
rect 24268 3408 24274 3420
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 26142 3448 26148 3460
rect 25372 3420 26148 3448
rect 25372 3408 25378 3420
rect 26142 3408 26148 3420
rect 26200 3408 26206 3460
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 27522 3448 27528 3460
rect 26568 3420 27528 3448
rect 26568 3408 26574 3420
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 33042 3448 33048 3460
rect 32456 3420 33048 3448
rect 32456 3408 32462 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 34422 3448 34428 3460
rect 33652 3420 34428 3448
rect 33652 3408 33658 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 34532 3420 84194 3448
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 34532 3380 34560 3420
rect 27764 3352 34560 3380
rect 27764 3340 27770 3352
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42702 3380 42708 3392
rect 41932 3352 42708 3380
rect 41932 3340 41938 3352
rect 42702 3340 42708 3352
rect 42760 3340 42766 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 44082 3380 44088 3392
rect 43128 3352 44088 3380
rect 43128 3340 43134 3352
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 84166 3312 84194 3420
rect 84470 3408 84476 3460
rect 84528 3448 84534 3460
rect 85482 3448 85488 3460
rect 84528 3420 85488 3448
rect 84528 3408 84534 3420
rect 85482 3408 85488 3420
rect 85540 3408 85546 3460
rect 95142 3340 95148 3392
rect 95200 3380 95206 3392
rect 100864 3380 100892 3488
rect 222838 3476 222844 3488
rect 222896 3476 222902 3528
rect 177298 3448 177304 3460
rect 95200 3352 100892 3380
rect 103486 3420 177304 3448
rect 95200 3340 95206 3352
rect 103486 3312 103514 3420
rect 177298 3408 177304 3420
rect 177356 3408 177362 3460
rect 84166 3284 103514 3312
rect 101030 3136 101036 3188
rect 101088 3176 101094 3188
rect 102042 3176 102048 3188
rect 101088 3148 102048 3176
rect 101088 3136 101094 3148
rect 102042 3136 102048 3148
rect 102100 3136 102106 3188
rect 110506 3136 110512 3188
rect 110564 3176 110570 3188
rect 111702 3176 111708 3188
rect 110564 3148 111708 3176
rect 110564 3136 110570 3148
rect 111702 3136 111708 3148
rect 111760 3136 111766 3188
rect 233878 3000 233884 3052
rect 233936 3040 233942 3052
rect 235810 3040 235816 3052
rect 233936 3012 235816 3040
rect 233936 3000 233942 3012
rect 235810 3000 235816 3012
rect 235868 3000 235874 3052
rect 92750 2864 92756 2916
rect 92808 2904 92814 2916
rect 93762 2904 93768 2916
rect 92808 2876 93768 2904
rect 92808 2864 92814 2876
rect 93762 2864 93768 2876
rect 93820 2864 93826 2916
rect 7650 2116 7656 2168
rect 7708 2156 7714 2168
rect 65426 2156 65432 2168
rect 7708 2128 65432 2156
rect 7708 2116 7714 2128
rect 65426 2116 65432 2128
rect 65484 2116 65490 2168
rect 63218 2048 63224 2100
rect 63276 2088 63282 2100
rect 264238 2088 264244 2100
rect 63276 2060 264244 2088
rect 63276 2048 63282 2060
rect 264238 2048 264244 2060
rect 264296 2048 264302 2100
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 235172 700340 235224 700392
rect 252560 700340 252612 700392
rect 269764 700340 269816 700392
rect 283840 700340 283892 700392
rect 395344 700340 395396 700392
rect 494796 700340 494848 700392
rect 24308 700272 24360 700324
rect 215944 700272 215996 700324
rect 238024 700272 238076 700324
rect 413652 700272 413704 700324
rect 453304 700272 453356 700324
rect 462320 700272 462372 700324
rect 497464 700272 497516 700324
rect 559656 700272 559708 700324
rect 154120 700068 154172 700120
rect 155224 700068 155276 700120
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 363604 699660 363656 699712
rect 364984 699660 365036 699712
rect 475384 699660 475436 699712
rect 478512 699660 478564 699712
rect 249064 698912 249116 698964
rect 527180 698912 527232 698964
rect 266360 697620 266412 697672
rect 267648 697620 267700 697672
rect 180708 697552 180760 697604
rect 397460 697552 397512 697604
rect 222844 696192 222896 696244
rect 348792 696192 348844 696244
rect 3516 670692 3568 670744
rect 196624 670692 196676 670744
rect 73068 665796 73120 665848
rect 240508 665796 240560 665848
rect 202144 660288 202196 660340
rect 331220 660288 331272 660340
rect 3516 656888 3568 656940
rect 112444 656888 112496 656940
rect 3516 632068 3568 632120
rect 166264 632068 166316 632120
rect 191748 623024 191800 623076
rect 299480 623024 299532 623076
rect 2780 619080 2832 619132
rect 4804 619080 4856 619132
rect 3516 605820 3568 605872
rect 220084 605820 220136 605872
rect 3332 579640 3384 579692
rect 226984 579640 227036 579692
rect 3240 565836 3292 565888
rect 68284 565836 68336 565888
rect 3332 553392 3384 553444
rect 35164 553392 35216 553444
rect 2964 527144 3016 527196
rect 71044 527144 71096 527196
rect 3516 514768 3568 514820
rect 162124 514768 162176 514820
rect 3056 500964 3108 501016
rect 233884 500964 233936 501016
rect 3056 474716 3108 474768
rect 244924 474716 244976 474768
rect 3424 462952 3476 463004
rect 258080 462952 258132 463004
rect 188988 456764 189040 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 204904 448536 204956 448588
rect 309784 430584 309836 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 21364 422288 21416 422340
rect 2872 409844 2924 409896
rect 29644 409844 29696 409896
rect 206284 404336 206336 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 177304 397468 177356 397520
rect 21364 382916 21416 382968
rect 209044 382916 209096 382968
rect 198648 380128 198700 380180
rect 583576 380128 583628 380180
rect 3424 371220 3476 371272
rect 21364 371220 21416 371272
rect 305644 364352 305696 364404
rect 579620 364352 579672 364404
rect 3148 357416 3200 357468
rect 15844 357416 15896 357468
rect 246304 356668 246356 356720
rect 583024 356668 583076 356720
rect 3332 345040 3384 345092
rect 232504 345040 232556 345092
rect 15844 338716 15896 338768
rect 228364 338716 228416 338768
rect 3332 318792 3384 318844
rect 224224 318792 224276 318844
rect 566464 311856 566516 311908
rect 579988 311856 580040 311908
rect 3424 304988 3476 305040
rect 249984 304988 250036 305040
rect 260196 302200 260248 302252
rect 266360 302200 266412 302252
rect 226248 300092 226300 300144
rect 583300 300092 583352 300144
rect 214564 298732 214616 298784
rect 580264 298732 580316 298784
rect 209688 296692 209740 296744
rect 264244 296692 264296 296744
rect 235724 295944 235776 295996
rect 475384 295944 475436 295996
rect 202788 294652 202840 294704
rect 244280 294652 244332 294704
rect 213828 294584 213880 294636
rect 582380 294584 582432 294636
rect 227628 293972 227680 294024
rect 273904 293972 273956 294024
rect 195796 293224 195848 293276
rect 429200 293224 429252 293276
rect 219348 292680 219400 292732
rect 251180 292680 251232 292732
rect 232596 292612 232648 292664
rect 305000 292612 305052 292664
rect 3424 292544 3476 292596
rect 11704 292544 11756 292596
rect 236920 292544 236972 292596
rect 583668 292544 583720 292596
rect 224224 291932 224276 291984
rect 240140 291932 240192 291984
rect 112444 291864 112496 291916
rect 245660 291864 245712 291916
rect 211068 291796 211120 291848
rect 583024 291796 583076 291848
rect 224868 291252 224920 291304
rect 247040 291252 247092 291304
rect 242716 291184 242768 291236
rect 271144 291184 271196 291236
rect 89628 290504 89680 290556
rect 232780 290504 232832 290556
rect 232504 290436 232556 290488
rect 243820 290436 243872 290488
rect 20 290096 72 290148
rect 242900 290096 242952 290148
rect 216496 290028 216548 290080
rect 253940 290028 253992 290080
rect 215208 289960 215260 290012
rect 260840 289960 260892 290012
rect 235816 289892 235868 289944
rect 260104 289892 260156 289944
rect 239956 289824 240008 289876
rect 574744 289824 574796 289876
rect 215944 289756 215996 289808
rect 218244 289756 218296 289808
rect 200396 289144 200448 289196
rect 206284 289144 206336 289196
rect 155224 289076 155276 289128
rect 204260 289076 204312 289128
rect 233884 289076 233936 289128
rect 245844 289076 245896 289128
rect 236644 288600 236696 288652
rect 249800 288600 249852 288652
rect 240876 288532 240928 288584
rect 255964 288532 256016 288584
rect 237380 288464 237432 288516
rect 265624 288464 265676 288516
rect 206652 288396 206704 288448
rect 583024 288396 583076 288448
rect 220084 288328 220136 288380
rect 225420 288328 225472 288380
rect 235908 288328 235960 288380
rect 238024 288328 238076 288380
rect 229836 287376 229888 287428
rect 255320 287376 255372 287428
rect 239588 287308 239640 287360
rect 267004 287308 267056 287360
rect 57244 287240 57296 287292
rect 230388 287240 230440 287292
rect 233148 287240 233200 287292
rect 302884 287240 302936 287292
rect 201316 287172 201368 287224
rect 309140 287172 309192 287224
rect 201684 287104 201736 287156
rect 334624 287104 334676 287156
rect 196624 287036 196676 287088
rect 202788 287036 202840 287088
rect 222108 287036 222160 287088
rect 302240 287036 302292 287088
rect 218612 286424 218664 286476
rect 222844 286424 222896 286476
rect 208492 286356 208544 286408
rect 232596 286356 232648 286408
rect 210884 286288 210936 286340
rect 236644 286288 236696 286340
rect 195888 286016 195940 286068
rect 203156 286016 203208 286068
rect 231676 286016 231728 286068
rect 244004 286016 244056 286068
rect 182088 285948 182140 286000
rect 204628 285948 204680 286000
rect 236092 285948 236144 286000
rect 253204 285948 253256 286000
rect 43444 285880 43496 285932
rect 206100 285880 206152 285932
rect 232228 285880 232280 285932
rect 262864 285880 262916 285932
rect 194508 285812 194560 285864
rect 203708 285812 203760 285864
rect 200028 285744 200080 285796
rect 207020 285812 207072 285864
rect 227812 285812 227864 285864
rect 276664 285812 276716 285864
rect 199936 285676 199988 285728
rect 205548 285744 205600 285796
rect 213460 285744 213512 285796
rect 214564 285744 214616 285796
rect 214748 285744 214800 285796
rect 221188 285744 221240 285796
rect 221556 285744 221608 285796
rect 204904 285676 204956 285728
rect 208124 285676 208176 285728
rect 209964 285676 210016 285728
rect 211068 285676 211120 285728
rect 212908 285676 212960 285728
rect 213828 285676 213880 285728
rect 214380 285676 214432 285728
rect 215208 285676 215260 285728
rect 215300 285676 215352 285728
rect 216588 285676 216640 285728
rect 223580 285676 223632 285728
rect 224868 285676 224920 285728
rect 226524 285676 226576 285728
rect 227628 285676 227680 285728
rect 234620 285744 234672 285796
rect 235724 285744 235776 285796
rect 239036 285744 239088 285796
rect 239956 285744 240008 285796
rect 241980 285744 242032 285796
rect 291200 285744 291252 285796
rect 303620 285676 303672 285728
rect 240140 285268 240192 285320
rect 241060 285268 241112 285320
rect 215852 284928 215904 284980
rect 237380 284928 237432 284980
rect 221188 284656 221240 284708
rect 264336 284656 264388 284708
rect 237012 284588 237064 284640
rect 249892 284588 249944 284640
rect 212356 284520 212408 284572
rect 249156 284520 249208 284572
rect 173164 284452 173216 284504
rect 223948 284452 224000 284504
rect 238116 284452 238168 284504
rect 261484 284452 261536 284504
rect 65524 284384 65576 284436
rect 213828 284384 213880 284436
rect 237564 284384 237616 284436
rect 244096 284384 244148 284436
rect 17224 284316 17276 284368
rect 227444 284316 227496 284368
rect 239956 284316 240008 284368
rect 299480 284316 299532 284368
rect 201500 284180 201552 284232
rect 202144 284180 202196 284232
rect 234528 283908 234580 283960
rect 284300 283840 284352 283892
rect 244096 283568 244148 283620
rect 282920 283568 282972 283620
rect 246028 282820 246080 282872
rect 583576 282820 583628 282872
rect 183468 281596 183520 281648
rect 197452 281596 197504 281648
rect 51724 281528 51776 281580
rect 197360 281528 197412 281580
rect 245936 281528 245988 281580
rect 254032 281528 254084 281580
rect 246028 280236 246080 280288
rect 268384 280236 268436 280288
rect 245936 280168 245988 280220
rect 271236 280168 271288 280220
rect 188896 278740 188948 278792
rect 197360 278740 197412 278792
rect 245936 278740 245988 278792
rect 583576 278740 583628 278792
rect 245936 278128 245988 278180
rect 249984 278128 250036 278180
rect 194416 277720 194468 277772
rect 197360 277720 197412 277772
rect 245936 277380 245988 277432
rect 583484 277380 583536 277432
rect 191656 276020 191708 276072
rect 197452 276020 197504 276072
rect 246028 276020 246080 276072
rect 280804 276020 280856 276072
rect 4804 275952 4856 276004
rect 197360 275952 197412 276004
rect 245936 275952 245988 276004
rect 583852 275952 583904 276004
rect 245936 275340 245988 275392
rect 249064 275340 249116 275392
rect 187608 274660 187660 274712
rect 197360 274660 197412 274712
rect 8208 273912 8260 273964
rect 178040 273912 178092 273964
rect 190368 273300 190420 273352
rect 197452 273300 197504 273352
rect 245936 273300 245988 273352
rect 256700 273300 256752 273352
rect 184848 273232 184900 273284
rect 197360 273232 197412 273284
rect 246028 273232 246080 273284
rect 295340 273232 295392 273284
rect 171048 273164 171100 273216
rect 197452 273164 197504 273216
rect 246028 271940 246080 271992
rect 255412 271940 255464 271992
rect 245936 271872 245988 271924
rect 267096 271872 267148 271924
rect 304264 271872 304316 271924
rect 579804 271872 579856 271924
rect 300124 271124 300176 271176
rect 580356 271124 580408 271176
rect 187516 270580 187568 270632
rect 197360 270580 197412 270632
rect 246028 270580 246080 270632
rect 258172 270580 258224 270632
rect 186228 270512 186280 270564
rect 197452 270512 197504 270564
rect 245936 270512 245988 270564
rect 276756 270512 276808 270564
rect 193128 269152 193180 269204
rect 197452 269152 197504 269204
rect 54484 269084 54536 269136
rect 197360 269084 197412 269136
rect 245936 269084 245988 269136
rect 285680 269084 285732 269136
rect 68284 269016 68336 269068
rect 197452 269016 197504 269068
rect 178040 268948 178092 269000
rect 197360 268948 197412 269000
rect 246028 267792 246080 267844
rect 268476 267792 268528 267844
rect 245936 267724 245988 267776
rect 583852 267724 583904 267776
rect 166264 267656 166316 267708
rect 197360 267656 197412 267708
rect 3056 266364 3108 266416
rect 170404 266364 170456 266416
rect 195612 266364 195664 266416
rect 197912 266364 197964 266416
rect 246028 266364 246080 266416
rect 269856 266364 269908 266416
rect 245936 266296 245988 266348
rect 566464 266296 566516 266348
rect 15844 264936 15896 264988
rect 197452 264936 197504 264988
rect 245844 264936 245896 264988
rect 251272 264936 251324 264988
rect 35164 264868 35216 264920
rect 197360 264868 197412 264920
rect 184756 263576 184808 263628
rect 197360 263576 197412 263628
rect 245936 263576 245988 263628
rect 248420 263576 248472 263628
rect 193036 262216 193088 262268
rect 197452 262216 197504 262268
rect 245936 262216 245988 262268
rect 259460 262216 259512 262268
rect 71044 262148 71096 262200
rect 197360 262148 197412 262200
rect 245844 260856 245896 260908
rect 258264 260856 258316 260908
rect 244924 260720 244976 260772
rect 245844 260720 245896 260772
rect 187424 259428 187476 259480
rect 197360 259428 197412 259480
rect 245936 259428 245988 259480
rect 300860 259428 300912 259480
rect 249156 259360 249208 259412
rect 580172 259360 580224 259412
rect 191564 258544 191616 258596
rect 197452 258544 197504 258596
rect 246028 258136 246080 258188
rect 287060 258136 287112 258188
rect 32404 258068 32456 258120
rect 197360 258068 197412 258120
rect 245936 258068 245988 258120
rect 294052 258068 294104 258120
rect 3516 257320 3568 257372
rect 178684 257320 178736 257372
rect 246396 257320 246448 257372
rect 583300 257320 583352 257372
rect 195704 256776 195756 256828
rect 197544 256776 197596 256828
rect 188804 256708 188856 256760
rect 197360 256708 197412 256760
rect 245936 256708 245988 256760
rect 272524 256708 272576 256760
rect 195796 256640 195848 256692
rect 197912 256640 197964 256692
rect 245752 256640 245804 256692
rect 583392 256640 583444 256692
rect 192944 255280 192996 255332
rect 197360 255280 197412 255332
rect 137928 254532 137980 254584
rect 147680 254532 147732 254584
rect 246488 254532 246540 254584
rect 582748 254532 582800 254584
rect 191472 253988 191524 254040
rect 197452 253988 197504 254040
rect 18604 253920 18656 253972
rect 197360 253920 197412 253972
rect 245936 253920 245988 253972
rect 252652 253920 252704 253972
rect 186136 253172 186188 253224
rect 198004 253172 198056 253224
rect 194324 252968 194376 253020
rect 198096 252968 198148 253020
rect 245936 252628 245988 252680
rect 306380 252628 306432 252680
rect 180616 252560 180668 252612
rect 197360 252560 197412 252612
rect 245844 252560 245896 252612
rect 306472 252560 306524 252612
rect 245936 252492 245988 252544
rect 258080 252492 258132 252544
rect 245936 251200 245988 251252
rect 583392 251200 583444 251252
rect 147680 251132 147732 251184
rect 197360 251132 197412 251184
rect 255964 250452 256016 250504
rect 582748 250452 582800 250504
rect 245844 249772 245896 249824
rect 307760 249772 307812 249824
rect 245936 249704 245988 249756
rect 252560 249704 252612 249756
rect 190276 248480 190328 248532
rect 197360 248480 197412 248532
rect 188712 248412 188764 248464
rect 197452 248412 197504 248464
rect 180708 248344 180760 248396
rect 197360 248344 197412 248396
rect 245844 248344 245896 248396
rect 583760 248344 583812 248396
rect 245936 248276 245988 248328
rect 309784 248276 309836 248328
rect 195796 247052 195848 247104
rect 197636 247052 197688 247104
rect 29644 246984 29696 247036
rect 197360 246984 197412 247036
rect 245936 245624 245988 245676
rect 305184 245624 305236 245676
rect 245936 244264 245988 244316
rect 251364 244264 251416 244316
rect 11704 244196 11756 244248
rect 197360 244196 197412 244248
rect 191748 244128 191800 244180
rect 197452 244128 197504 244180
rect 583852 243584 583904 243636
rect 582748 243516 582800 243568
rect 583760 243516 583812 243568
rect 583852 243380 583904 243432
rect 245844 242904 245896 242956
rect 273996 242904 274048 242956
rect 188988 242836 189040 242888
rect 197360 242836 197412 242888
rect 3424 242156 3476 242208
rect 180064 242156 180116 242208
rect 245844 241544 245896 241596
rect 269948 241544 270000 241596
rect 191748 241476 191800 241528
rect 197452 241476 197504 241528
rect 244096 241476 244148 241528
rect 579620 241476 579672 241528
rect 199108 240184 199160 240236
rect 246028 240388 246080 240440
rect 245936 240320 245988 240372
rect 255504 240320 255556 240372
rect 269764 240252 269816 240304
rect 453304 240184 453356 240236
rect 3424 240116 3476 240168
rect 213184 240116 213236 240168
rect 240508 240116 240560 240168
rect 240600 240116 240652 240168
rect 240968 240116 241020 240168
rect 225236 240048 225288 240100
rect 235908 240048 235960 240100
rect 582472 240116 582524 240168
rect 241152 240048 241204 240100
rect 582564 240048 582616 240100
rect 170404 239980 170456 240032
rect 212724 239980 212776 240032
rect 238852 239980 238904 240032
rect 234988 239912 235040 239964
rect 240968 239912 241020 239964
rect 497464 239980 497516 240032
rect 162124 239844 162176 239896
rect 242716 239844 242768 239896
rect 232596 239776 232648 239828
rect 395344 239912 395396 239964
rect 199844 239504 199896 239556
rect 209136 239504 209188 239556
rect 207940 239436 207992 239488
rect 288624 239436 288676 239488
rect 106188 239368 106240 239420
rect 209780 239368 209832 239420
rect 209780 238688 209832 238740
rect 214564 238688 214616 238740
rect 239220 238688 239272 238740
rect 244096 238688 244148 238740
rect 180064 238620 180116 238672
rect 231492 238620 231544 238672
rect 236460 238620 236512 238672
rect 582932 238620 582984 238672
rect 177304 238552 177356 238604
rect 209228 238552 209280 238604
rect 216036 238552 216088 238604
rect 304264 238552 304316 238604
rect 216588 238484 216640 238536
rect 300124 238484 300176 238536
rect 21364 238416 21416 238468
rect 221924 238416 221976 238468
rect 227628 238416 227680 238468
rect 260196 238416 260248 238468
rect 233516 238348 233568 238400
rect 583116 238348 583168 238400
rect 223764 238280 223816 238332
rect 224776 238280 224828 238332
rect 234068 238280 234120 238332
rect 234528 238280 234580 238332
rect 206468 238212 206520 238264
rect 206928 238212 206980 238264
rect 211252 238076 211304 238128
rect 220084 238076 220136 238128
rect 214196 238008 214248 238060
rect 215024 238008 215076 238060
rect 220452 238008 220504 238060
rect 238760 238008 238812 238060
rect 222844 237940 222896 237992
rect 223488 237940 223540 237992
rect 230572 237804 230624 237856
rect 231768 237804 231820 237856
rect 201500 237736 201552 237788
rect 202696 237736 202748 237788
rect 200212 237668 200264 237720
rect 201316 237668 201368 237720
rect 205916 237668 205968 237720
rect 206744 237668 206796 237720
rect 207388 237668 207440 237720
rect 208216 237668 208268 237720
rect 201132 237532 201184 237584
rect 209044 237532 209096 237584
rect 202972 237464 203024 237516
rect 203892 237464 203944 237516
rect 218060 237464 218112 237516
rect 220176 237464 220228 237516
rect 200580 237396 200632 237448
rect 201408 237396 201460 237448
rect 203524 237396 203576 237448
rect 203984 237396 204036 237448
rect 208400 237396 208452 237448
rect 210332 237396 210384 237448
rect 211804 237396 211856 237448
rect 212448 237396 212500 237448
rect 213092 237396 213144 237448
rect 213736 237396 213788 237448
rect 215668 237396 215720 237448
rect 216588 237396 216640 237448
rect 218428 237396 218480 237448
rect 219256 237396 219308 237448
rect 219900 237396 219952 237448
rect 220728 237396 220780 237448
rect 221004 237396 221056 237448
rect 222016 237396 222068 237448
rect 225788 237396 225840 237448
rect 226248 237396 226300 237448
rect 226708 237396 226760 237448
rect 227628 237396 227680 237448
rect 232044 237396 232096 237448
rect 233148 237396 233200 237448
rect 236828 237396 236880 237448
rect 237288 237396 237340 237448
rect 237380 237396 237432 237448
rect 238668 237396 238720 237448
rect 240324 237396 240376 237448
rect 241428 237396 241480 237448
rect 41328 237328 41380 237380
rect 219532 237328 219584 237380
rect 221372 237328 221424 237380
rect 363604 237328 363656 237380
rect 235264 236784 235316 236836
rect 243268 236784 243320 236836
rect 217140 236648 217192 236700
rect 232136 236648 232188 236700
rect 235356 236648 235408 236700
rect 582656 236648 582708 236700
rect 240508 236104 240560 236156
rect 240968 236104 241020 236156
rect 202052 235900 202104 235952
rect 305644 235900 305696 235952
rect 22744 235288 22796 235340
rect 230204 235356 230256 235408
rect 229100 235288 229152 235340
rect 295432 235288 295484 235340
rect 212172 235220 212224 235272
rect 582472 235220 582524 235272
rect 243636 234064 243688 234116
rect 293960 234064 294012 234116
rect 227260 233996 227312 234048
rect 289820 233996 289872 234048
rect 170404 233928 170456 233980
rect 245752 233928 245804 233980
rect 3424 233860 3476 233912
rect 208400 233860 208452 233912
rect 209872 233860 209924 233912
rect 582748 233860 582800 233912
rect 239404 233520 239456 233572
rect 242164 233520 242216 233572
rect 231124 233180 231176 233232
rect 233332 233180 233384 233232
rect 195612 232568 195664 232620
rect 303712 232568 303764 232620
rect 4804 232500 4856 232552
rect 229652 232500 229704 232552
rect 222292 231140 222344 231192
rect 278044 231140 278096 231192
rect 204996 231072 205048 231124
rect 582564 231072 582616 231124
rect 178684 229848 178736 229900
rect 245660 229848 245712 229900
rect 218980 229780 219032 229832
rect 288716 229780 288768 229832
rect 194324 229712 194376 229764
rect 298284 229712 298336 229764
rect 241336 228420 241388 228472
rect 291292 228420 291344 228472
rect 196992 228352 197044 228404
rect 276848 228352 276900 228404
rect 222016 227060 222068 227112
rect 302332 227060 302384 227112
rect 203984 226992 204036 227044
rect 292580 226992 292632 227044
rect 226156 225564 226208 225616
rect 305092 225564 305144 225616
rect 220728 224204 220780 224256
rect 282184 224204 282236 224256
rect 352564 224204 352616 224256
rect 580264 224204 580316 224256
rect 202696 221416 202748 221468
rect 285772 221416 285824 221468
rect 224684 218696 224736 218748
rect 299664 218696 299716 218748
rect 201316 215908 201368 215960
rect 296812 215908 296864 215960
rect 3332 215228 3384 215280
rect 15844 215228 15896 215280
rect 233148 213188 233200 213240
rect 288532 213188 288584 213240
rect 188804 211760 188856 211812
rect 296720 211760 296772 211812
rect 208216 210400 208268 210452
rect 280160 210400 280212 210452
rect 191472 209040 191524 209092
rect 582840 209040 582892 209092
rect 302884 206932 302936 206984
rect 579804 206932 579856 206984
rect 219256 204892 219308 204944
rect 284392 204892 284444 204944
rect 209136 203600 209188 203652
rect 214564 203600 214616 203652
rect 205456 203532 205508 203584
rect 289912 203532 289964 203584
rect 3056 202784 3108 202836
rect 170404 202784 170456 202836
rect 215024 202104 215076 202156
rect 307852 202104 307904 202156
rect 233884 201832 233936 201884
rect 237932 201832 237984 201884
rect 204904 200744 204956 200796
rect 299572 200744 299624 200796
rect 220176 199384 220228 199436
rect 230756 199384 230808 199436
rect 227628 197956 227680 198008
rect 291384 197956 291436 198008
rect 198464 196596 198516 196648
rect 279056 196596 279108 196648
rect 199844 195304 199896 195356
rect 245660 195304 245712 195356
rect 217876 195236 217928 195288
rect 300952 195236 301004 195288
rect 180616 193808 180668 193860
rect 271328 193808 271380 193860
rect 334624 193128 334676 193180
rect 580172 193128 580224 193180
rect 187608 192516 187660 192568
rect 242900 192516 242952 192568
rect 220084 192448 220136 192500
rect 292764 192448 292816 192500
rect 214564 189932 214616 189984
rect 240416 189932 240468 189984
rect 182088 189864 182140 189916
rect 228364 189864 228416 189916
rect 197176 189796 197228 189848
rect 278780 189796 278832 189848
rect 192944 189728 192996 189780
rect 302424 189728 302476 189780
rect 3516 188980 3568 189032
rect 173164 188980 173216 189032
rect 195704 188368 195756 188420
rect 230572 188368 230624 188420
rect 203892 188300 203944 188352
rect 285864 188300 285916 188352
rect 204168 187076 204220 187128
rect 244464 187076 244516 187128
rect 188712 187008 188764 187060
rect 248512 187008 248564 187060
rect 193036 186940 193088 186992
rect 287244 186940 287296 186992
rect 261484 185648 261536 185700
rect 291476 185648 291528 185700
rect 226248 185580 226300 185632
rect 282184 185580 282236 185632
rect 285956 185580 286008 185632
rect 284484 185512 284536 185564
rect 213828 184492 213880 184544
rect 242992 184492 243044 184544
rect 206836 184424 206888 184476
rect 236000 184424 236052 184476
rect 197084 184356 197136 184408
rect 240140 184356 240192 184408
rect 240416 184356 240468 184408
rect 278136 184356 278188 184408
rect 199936 184288 199988 184340
rect 245752 184288 245804 184340
rect 229008 184220 229060 184272
rect 302516 184220 302568 184272
rect 191656 184152 191708 184204
rect 290096 184152 290148 184204
rect 272524 182860 272576 182912
rect 298376 182860 298428 182912
rect 246396 182792 246448 182844
rect 287152 182792 287204 182844
rect 262864 181704 262916 181756
rect 281540 181704 281592 181756
rect 183468 181636 183520 181688
rect 241612 181636 241664 181688
rect 267004 181636 267056 181688
rect 296904 181636 296956 181688
rect 187424 181568 187476 181620
rect 247224 181568 247276 181620
rect 253204 181568 253256 181620
rect 295616 181568 295668 181620
rect 234528 181500 234580 181552
rect 303804 181500 303856 181552
rect 202604 181432 202656 181484
rect 283472 181432 283524 181484
rect 130936 181024 130988 181076
rect 173256 181024 173308 181076
rect 128176 180956 128228 181008
rect 184388 180956 184440 181008
rect 102048 180888 102100 180940
rect 169024 180888 169076 180940
rect 99472 180820 99524 180872
rect 203524 180820 203576 180872
rect 273904 180276 273956 180328
rect 294144 180276 294196 180328
rect 215208 180208 215260 180260
rect 237564 180208 237616 180260
rect 260104 180208 260156 180260
rect 292672 180208 292724 180260
rect 200028 180140 200080 180192
rect 230664 180140 230716 180192
rect 237288 180140 237340 180192
rect 283196 180140 283248 180192
rect 201408 180072 201460 180124
rect 292856 180072 292908 180124
rect 129464 179732 129516 179784
rect 168380 179732 168432 179784
rect 123300 179664 123352 179716
rect 175924 179664 175976 179716
rect 121276 179596 121328 179648
rect 177396 179596 177448 179648
rect 110696 179528 110748 179580
rect 182824 179528 182876 179580
rect 108120 179460 108172 179512
rect 181444 179460 181496 179512
rect 114560 179392 114612 179444
rect 214564 179392 214616 179444
rect 224776 178984 224828 179036
rect 231952 178984 232004 179036
rect 269948 178984 270000 179036
rect 284576 178984 284628 179036
rect 212448 178916 212500 178968
rect 229468 178916 229520 178968
rect 268384 178916 268436 178968
rect 290004 178916 290056 178968
rect 206928 178848 206980 178900
rect 237472 178848 237524 178900
rect 271236 178848 271288 178900
rect 296996 178848 297048 178900
rect 195796 178780 195848 178832
rect 236092 178780 236144 178832
rect 267096 178780 267148 178832
rect 295524 178780 295576 178832
rect 186136 178712 186188 178764
rect 229192 178712 229244 178764
rect 241428 178712 241480 178764
rect 279240 178712 279292 178764
rect 184756 178644 184808 178696
rect 236184 178644 236236 178696
rect 238668 178644 238720 178696
rect 283380 178644 283432 178696
rect 132408 178372 132460 178424
rect 165344 178372 165396 178424
rect 112260 178304 112312 178356
rect 166356 178304 166408 178356
rect 116952 178236 117004 178288
rect 174544 178236 174596 178288
rect 125968 178168 126020 178220
rect 186964 178168 187016 178220
rect 109592 178100 109644 178152
rect 180064 178100 180116 178152
rect 119528 178032 119580 178084
rect 200764 178032 200816 178084
rect 223396 177964 223448 178016
rect 229376 177964 229428 178016
rect 271328 177556 271380 177608
rect 288440 177556 288492 177608
rect 278136 177488 278188 177540
rect 301044 177488 301096 177540
rect 219348 177420 219400 177472
rect 234804 177420 234856 177472
rect 269856 177420 269908 177472
rect 294236 177420 294288 177472
rect 208308 177352 208360 177404
rect 279148 177352 279200 177404
rect 198648 177284 198700 177336
rect 280344 177284 280396 177336
rect 105728 177080 105780 177132
rect 191104 177080 191156 177132
rect 134432 177012 134484 177064
rect 165436 177012 165488 177064
rect 127164 176944 127216 176996
rect 167736 176944 167788 176996
rect 158904 176876 158956 176928
rect 207664 176876 207716 176928
rect 148232 176808 148284 176860
rect 198096 176808 198148 176860
rect 107016 176740 107068 176792
rect 170496 176740 170548 176792
rect 136088 176672 136140 176724
rect 213920 176604 213972 176656
rect 276848 176604 276900 176656
rect 283012 176604 283064 176656
rect 191564 176536 191616 176588
rect 241520 176536 241572 176588
rect 280804 176536 280856 176588
rect 287336 176536 287388 176588
rect 278044 176468 278096 176520
rect 280252 176468 280304 176520
rect 133144 176196 133196 176248
rect 165528 176196 165580 176248
rect 124496 176128 124548 176180
rect 166448 176128 166500 176180
rect 276756 176128 276808 176180
rect 279332 176128 279384 176180
rect 121920 176060 121972 176112
rect 169116 176060 169168 176112
rect 224868 176060 224920 176112
rect 231860 176060 231912 176112
rect 276664 176060 276716 176112
rect 280436 176060 280488 176112
rect 118424 175992 118476 176044
rect 173164 175992 173216 176044
rect 223488 175992 223540 176044
rect 232044 175992 232096 176044
rect 273996 175992 274048 176044
rect 281632 175992 281684 176044
rect 115756 175924 115808 175976
rect 184296 175924 184348 175976
rect 188896 175924 188948 175976
rect 230940 175924 230992 175976
rect 268476 175924 268528 175976
rect 281816 175924 281868 175976
rect 220912 175788 220964 175840
rect 224224 175788 224276 175840
rect 165436 175176 165488 175228
rect 213920 175176 213972 175228
rect 165528 175108 165580 175160
rect 214012 175108 214064 175160
rect 246396 175244 246448 175296
rect 264980 175244 265032 175296
rect 229284 175176 229336 175228
rect 231124 175176 231176 175228
rect 256700 175176 256752 175228
rect 229008 175108 229060 175160
rect 231768 175108 231820 175160
rect 255504 175108 255556 175160
rect 194508 175040 194560 175092
rect 230480 174972 230532 175024
rect 209044 174496 209096 174548
rect 237656 174496 237708 174548
rect 257436 174020 257488 174072
rect 264980 174020 265032 174072
rect 229008 173952 229060 174004
rect 256148 173952 256200 174004
rect 265072 173952 265124 174004
rect 236276 173884 236328 173936
rect 252100 173884 252152 173936
rect 265256 173884 265308 173936
rect 165344 173816 165396 173868
rect 213920 173816 213972 173868
rect 231584 173816 231636 173868
rect 247132 173816 247184 173868
rect 173256 173748 173308 173800
rect 214012 173748 214064 173800
rect 229192 173612 229244 173664
rect 229376 173612 229428 173664
rect 281724 173544 281776 173596
rect 284300 173544 284352 173596
rect 229100 173204 229152 173256
rect 229468 173204 229520 173256
rect 247960 173136 248012 173188
rect 265164 173136 265216 173188
rect 240968 172660 241020 172712
rect 264980 172660 265032 172712
rect 260380 172524 260432 172576
rect 265072 172524 265124 172576
rect 168380 172456 168432 172508
rect 213920 172456 213972 172508
rect 231676 172456 231728 172508
rect 259460 172456 259512 172508
rect 184388 172388 184440 172440
rect 214012 172388 214064 172440
rect 231768 172388 231820 172440
rect 248420 172388 248472 172440
rect 282644 172388 282696 172440
rect 285956 172388 286008 172440
rect 231492 172184 231544 172236
rect 235264 172184 235316 172236
rect 262956 171504 263008 171556
rect 264980 171504 265032 171556
rect 250444 171164 250496 171216
rect 265072 171164 265124 171216
rect 167920 171096 167972 171148
rect 184204 171096 184256 171148
rect 249156 171096 249208 171148
rect 264980 171096 265032 171148
rect 167736 171028 167788 171080
rect 213920 171028 213972 171080
rect 231768 171028 231820 171080
rect 251180 171028 251232 171080
rect 186964 170960 187016 171012
rect 214012 170960 214064 171012
rect 231492 170960 231544 171012
rect 240232 170960 240284 171012
rect 231216 170756 231268 170808
rect 236092 170756 236144 170808
rect 281724 170620 281776 170672
rect 283472 170620 283524 170672
rect 258816 169872 258868 169924
rect 265164 169872 265216 169924
rect 257344 169804 257396 169856
rect 264980 169804 265032 169856
rect 239496 169736 239548 169788
rect 265072 169736 265124 169788
rect 166448 169668 166500 169720
rect 213920 169668 213972 169720
rect 231124 169668 231176 169720
rect 233424 169668 233476 169720
rect 175924 169600 175976 169652
rect 214012 169600 214064 169652
rect 231768 169532 231820 169584
rect 238760 169532 238812 169584
rect 282736 168716 282788 168768
rect 288624 168716 288676 168768
rect 282828 168648 282880 168700
rect 287244 168648 287296 168700
rect 260288 168580 260340 168632
rect 265256 168580 265308 168632
rect 254768 168512 254820 168564
rect 265072 168512 265124 168564
rect 253480 168444 253532 168496
rect 264980 168444 265032 168496
rect 244924 168376 244976 168428
rect 265164 168376 265216 168428
rect 169116 168308 169168 168360
rect 213920 168308 213972 168360
rect 231768 168308 231820 168360
rect 251364 168308 251416 168360
rect 282736 168308 282788 168360
rect 301044 168308 301096 168360
rect 177396 168240 177448 168292
rect 214012 168240 214064 168292
rect 231400 168240 231452 168292
rect 247040 168240 247092 168292
rect 282828 168240 282880 168292
rect 288440 168240 288492 168292
rect 231676 168036 231728 168088
rect 234804 168036 234856 168088
rect 261760 167084 261812 167136
rect 265164 167084 265216 167136
rect 241152 167016 241204 167068
rect 264980 167016 265032 167068
rect 173164 166948 173216 167000
rect 214104 166948 214156 167000
rect 174544 166880 174596 166932
rect 214012 166880 214064 166932
rect 200764 166812 200816 166864
rect 213920 166812 213972 166864
rect 231032 166676 231084 166728
rect 233884 166676 233936 166728
rect 231308 166540 231360 166592
rect 236184 166540 236236 166592
rect 251824 166336 251876 166388
rect 265072 166336 265124 166388
rect 231124 166268 231176 166320
rect 252652 166268 252704 166320
rect 230480 165860 230532 165912
rect 232136 165860 232188 165912
rect 253296 165656 253348 165708
rect 264980 165656 265032 165708
rect 242440 165588 242492 165640
rect 265072 165588 265124 165640
rect 171784 165520 171836 165572
rect 214012 165520 214064 165572
rect 231400 165520 231452 165572
rect 249892 165520 249944 165572
rect 282000 165520 282052 165572
rect 299664 165520 299716 165572
rect 184296 165452 184348 165504
rect 213920 165452 213972 165504
rect 282828 165452 282880 165504
rect 296812 165452 296864 165504
rect 231308 165112 231360 165164
rect 237564 165112 237616 165164
rect 250720 164840 250772 164892
rect 265164 164840 265216 164892
rect 261484 164296 261536 164348
rect 265072 164296 265124 164348
rect 236828 164228 236880 164280
rect 264980 164228 265032 164280
rect 3240 164160 3292 164212
rect 65524 164160 65576 164212
rect 166356 164160 166408 164212
rect 213920 164160 213972 164212
rect 231400 164160 231452 164212
rect 238852 164160 238904 164212
rect 178776 163480 178828 163532
rect 214932 163480 214984 163532
rect 235540 163072 235592 163124
rect 265164 163072 265216 163124
rect 246304 163004 246356 163056
rect 265072 163004 265124 163056
rect 242348 162936 242400 162988
rect 264980 162936 265032 162988
rect 180064 162800 180116 162852
rect 214012 162800 214064 162852
rect 231400 162800 231452 162852
rect 258264 162800 258316 162852
rect 282092 162800 282144 162852
rect 295616 162800 295668 162852
rect 182824 162732 182876 162784
rect 213920 162732 213972 162784
rect 230940 162732 230992 162784
rect 241612 162732 241664 162784
rect 231400 161848 231452 161900
rect 237472 161848 237524 161900
rect 247868 161508 247920 161560
rect 264980 161508 265032 161560
rect 238024 161440 238076 161492
rect 265164 161440 265216 161492
rect 170496 161372 170548 161424
rect 214012 161372 214064 161424
rect 230940 161372 230992 161424
rect 234436 161372 234488 161424
rect 181444 161304 181496 161356
rect 213920 161304 213972 161356
rect 231400 161168 231452 161220
rect 236276 161168 236328 161220
rect 282460 161168 282512 161220
rect 287336 161168 287388 161220
rect 229836 160760 229888 160812
rect 240140 160760 240192 160812
rect 234160 160692 234212 160744
rect 264980 160692 265032 160744
rect 260104 160216 260156 160268
rect 265164 160216 265216 160268
rect 243728 160148 243780 160200
rect 265072 160148 265124 160200
rect 240876 160080 240928 160132
rect 264980 160080 265032 160132
rect 170404 160012 170456 160064
rect 214012 160012 214064 160064
rect 231400 160012 231452 160064
rect 255412 160012 255464 160064
rect 282092 160012 282144 160064
rect 292856 160012 292908 160064
rect 191104 159944 191156 159996
rect 213920 159944 213972 159996
rect 230940 159944 230992 159996
rect 254032 159944 254084 159996
rect 258724 158856 258776 158908
rect 265164 158856 265216 158908
rect 257620 158788 257672 158840
rect 265072 158788 265124 158840
rect 236736 158720 236788 158772
rect 264980 158720 265032 158772
rect 167644 158652 167696 158704
rect 213920 158652 213972 158704
rect 282828 158652 282880 158704
rect 294052 158652 294104 158704
rect 169024 158584 169076 158636
rect 214012 158584 214064 158636
rect 231216 157972 231268 158024
rect 240968 157972 241020 158024
rect 258908 157496 258960 157548
rect 265164 157496 265216 157548
rect 254860 157428 254912 157480
rect 265072 157428 265124 157480
rect 238300 157360 238352 157412
rect 264980 157360 265032 157412
rect 203524 157292 203576 157344
rect 213920 157292 213972 157344
rect 231768 157292 231820 157344
rect 255320 157292 255372 157344
rect 231124 157224 231176 157276
rect 244372 157224 244424 157276
rect 255964 156068 256016 156120
rect 265072 156068 265124 156120
rect 241244 156000 241296 156052
rect 264980 156000 265032 156052
rect 234068 155932 234120 155984
rect 265164 155932 265216 155984
rect 166264 155864 166316 155916
rect 213920 155864 213972 155916
rect 230940 155864 230992 155916
rect 234712 155864 234764 155916
rect 177304 155796 177356 155848
rect 214012 155796 214064 155848
rect 232504 155184 232556 155236
rect 265624 155184 265676 155236
rect 249340 154640 249392 154692
rect 265072 154640 265124 154692
rect 239680 154572 239732 154624
rect 264980 154572 265032 154624
rect 231768 154504 231820 154556
rect 242992 154504 243044 154556
rect 281724 154504 281776 154556
rect 307852 154504 307904 154556
rect 231492 153960 231544 154012
rect 237656 153960 237708 154012
rect 253388 153824 253440 153876
rect 265164 153824 265216 153876
rect 180064 153280 180116 153332
rect 214012 153280 214064 153332
rect 252008 153280 252060 153332
rect 265072 153280 265124 153332
rect 166264 153212 166316 153264
rect 213920 153212 213972 153264
rect 232780 153212 232832 153264
rect 264980 153212 265032 153264
rect 231400 153144 231452 153196
rect 251272 153144 251324 153196
rect 231768 153076 231820 153128
rect 245752 153076 245804 153128
rect 229744 152532 229796 152584
rect 248512 152532 248564 152584
rect 229928 152464 229980 152516
rect 265348 152464 265400 152516
rect 184296 151852 184348 151904
rect 213920 151852 213972 151904
rect 251916 151852 251968 151904
rect 265072 151852 265124 151904
rect 170404 151784 170456 151836
rect 214012 151784 214064 151836
rect 245108 151784 245160 151836
rect 264980 151784 265032 151836
rect 282828 151716 282880 151768
rect 302516 151716 302568 151768
rect 231216 151580 231268 151632
rect 233332 151580 233384 151632
rect 282644 151240 282696 151292
rect 285864 151240 285916 151292
rect 250628 151104 250680 151156
rect 265164 151104 265216 151156
rect 200764 151036 200816 151088
rect 214472 151036 214524 151088
rect 231216 151036 231268 151088
rect 252100 151036 252152 151088
rect 198004 150424 198056 150476
rect 213920 150424 213972 150476
rect 249064 150424 249116 150476
rect 264980 150424 265032 150476
rect 3516 150356 3568 150408
rect 43444 150356 43496 150408
rect 184204 150356 184256 150408
rect 214012 150356 214064 150408
rect 230940 150356 230992 150408
rect 253940 150356 253992 150408
rect 282828 150356 282880 150408
rect 290096 150356 290148 150408
rect 198096 150288 198148 150340
rect 213920 150288 213972 150340
rect 230848 150288 230900 150340
rect 240784 150288 240836 150340
rect 234252 149744 234304 149796
rect 249800 149744 249852 149796
rect 246580 149676 246632 149728
rect 265256 149676 265308 149728
rect 281724 149608 281776 149660
rect 284576 149608 284628 149660
rect 263048 149200 263100 149252
rect 265440 149200 265492 149252
rect 253204 149132 253256 149184
rect 264980 149132 265032 149184
rect 235448 149064 235500 149116
rect 265072 149064 265124 149116
rect 207664 148996 207716 149048
rect 213920 148996 213972 149048
rect 231768 148996 231820 149048
rect 244464 148996 244516 149048
rect 282736 148996 282788 149048
rect 292764 148996 292816 149048
rect 282828 148928 282880 148980
rect 287060 148928 287112 148980
rect 231124 148316 231176 148368
rect 234620 148316 234672 148368
rect 231400 148248 231452 148300
rect 257436 148316 257488 148368
rect 262864 147840 262916 147892
rect 265348 147840 265400 147892
rect 260472 147772 260524 147824
rect 265072 147772 265124 147824
rect 264428 147704 264480 147756
rect 266084 147704 266136 147756
rect 166356 147636 166408 147688
rect 213920 147636 213972 147688
rect 250536 147636 250588 147688
rect 264980 147636 265032 147688
rect 256056 146888 256108 146940
rect 265164 146888 265216 146940
rect 202144 146344 202196 146396
rect 214012 146344 214064 146396
rect 245200 146344 245252 146396
rect 265072 146344 265124 146396
rect 195244 146276 195296 146328
rect 213920 146276 213972 146328
rect 232596 146276 232648 146328
rect 264980 146276 265032 146328
rect 231768 146208 231820 146260
rect 247224 146208 247276 146260
rect 282000 146208 282052 146260
rect 302424 146208 302476 146260
rect 282828 146140 282880 146192
rect 291200 146140 291252 146192
rect 231676 145392 231728 145444
rect 236000 145392 236052 145444
rect 247776 145052 247828 145104
rect 265072 145052 265124 145104
rect 191104 144984 191156 145036
rect 213920 144984 213972 145036
rect 242164 144984 242216 145036
rect 264980 144984 265032 145036
rect 184204 144916 184256 144968
rect 214012 144916 214064 144968
rect 235356 144916 235408 144968
rect 265164 144916 265216 144968
rect 231308 144848 231360 144900
rect 244280 144848 244332 144900
rect 282828 144848 282880 144900
rect 294236 144848 294288 144900
rect 231492 144780 231544 144832
rect 239404 144780 239456 144832
rect 237380 144168 237432 144220
rect 241796 144168 241848 144220
rect 249248 144168 249300 144220
rect 265256 144168 265308 144220
rect 198096 143624 198148 143676
rect 214012 143624 214064 143676
rect 242256 143624 242308 143676
rect 265072 143624 265124 143676
rect 188344 143556 188396 143608
rect 213920 143556 213972 143608
rect 239588 143556 239640 143608
rect 264980 143556 265032 143608
rect 281632 143488 281684 143540
rect 296996 143488 297048 143540
rect 231308 143352 231360 143404
rect 237380 143352 237432 143404
rect 256240 142264 256292 142316
rect 264980 142264 265032 142316
rect 241060 142196 241112 142248
rect 265164 142196 265216 142248
rect 186964 142128 187016 142180
rect 213920 142128 213972 142180
rect 238208 142128 238260 142180
rect 265072 142128 265124 142180
rect 231768 142060 231820 142112
rect 258172 142060 258224 142112
rect 282736 142060 282788 142112
rect 299756 142060 299808 142112
rect 282828 141992 282880 142044
rect 298376 141992 298428 142044
rect 282828 141380 282880 141432
rect 291476 141380 291528 141432
rect 252100 140904 252152 140956
rect 264980 140904 265032 140956
rect 189724 140836 189776 140888
rect 213920 140836 213972 140888
rect 240968 140836 241020 140888
rect 265072 140836 265124 140888
rect 177396 140768 177448 140820
rect 214012 140768 214064 140820
rect 233884 140768 233936 140820
rect 265164 140768 265216 140820
rect 231676 140700 231728 140752
rect 260840 140700 260892 140752
rect 281908 140700 281960 140752
rect 290004 140700 290056 140752
rect 231768 140632 231820 140684
rect 242900 140632 242952 140684
rect 206376 139476 206428 139528
rect 214012 139476 214064 139528
rect 187148 139408 187200 139460
rect 213920 139408 213972 139460
rect 243544 139408 243596 139460
rect 264980 139408 265032 139460
rect 231768 139340 231820 139392
rect 245660 139340 245712 139392
rect 583392 139340 583444 139392
rect 583852 139340 583904 139392
rect 177304 138660 177356 138712
rect 214932 138660 214984 138712
rect 231308 138660 231360 138712
rect 239496 138660 239548 138712
rect 254676 138048 254728 138100
rect 265072 138048 265124 138100
rect 185584 137980 185636 138032
rect 214012 137980 214064 138032
rect 239404 137980 239456 138032
rect 264980 137980 265032 138032
rect 3516 137912 3568 137964
rect 32404 137912 32456 137964
rect 282828 137912 282880 137964
rect 306472 137912 306524 137964
rect 231676 137844 231728 137896
rect 234252 137844 234304 137896
rect 240784 136756 240836 136808
rect 265072 136756 265124 136808
rect 236644 136688 236696 136740
rect 264980 136688 265032 136740
rect 169024 136620 169076 136672
rect 213920 136620 213972 136672
rect 233976 136620 234028 136672
rect 265256 136620 265308 136672
rect 282368 136552 282420 136604
rect 305000 136552 305052 136604
rect 282552 136348 282604 136400
rect 285772 136348 285824 136400
rect 182824 135872 182876 135924
rect 214104 135872 214156 135924
rect 231124 135872 231176 135924
rect 264520 135872 264572 135924
rect 229744 135464 229796 135516
rect 265072 135464 265124 135516
rect 257436 135396 257488 135448
rect 265164 135396 265216 135448
rect 209136 135328 209188 135380
rect 214012 135328 214064 135380
rect 245016 135328 245068 135380
rect 264980 135328 265032 135380
rect 181444 135260 181496 135312
rect 213920 135260 213972 135312
rect 231768 135192 231820 135244
rect 256148 135192 256200 135244
rect 231676 135124 231728 135176
rect 247960 135124 248012 135176
rect 247684 134036 247736 134088
rect 265072 134036 265124 134088
rect 239496 133968 239548 134020
rect 264980 133968 265032 134020
rect 173348 133900 173400 133952
rect 213920 133900 213972 133952
rect 238116 133900 238168 133952
rect 265164 133900 265216 133952
rect 231676 133832 231728 133884
rect 262956 133832 263008 133884
rect 231768 133764 231820 133816
rect 260380 133764 260432 133816
rect 231216 133560 231268 133612
rect 238300 133560 238352 133612
rect 260196 132812 260248 132864
rect 265072 132812 265124 132864
rect 261852 132744 261904 132796
rect 264980 132744 265032 132796
rect 263140 132608 263192 132660
rect 265900 132608 265952 132660
rect 175924 132540 175976 132592
rect 214012 132540 214064 132592
rect 173256 132472 173308 132524
rect 213920 132472 213972 132524
rect 231768 132404 231820 132456
rect 250444 132404 250496 132456
rect 282736 132404 282788 132456
rect 296904 132404 296956 132456
rect 231676 132336 231728 132388
rect 249156 132336 249208 132388
rect 282828 132336 282880 132388
rect 295340 132336 295392 132388
rect 250812 131724 250864 131776
rect 265808 131724 265860 131776
rect 167736 131112 167788 131164
rect 213920 131112 213972 131164
rect 231768 131044 231820 131096
rect 258816 131044 258868 131096
rect 282828 131044 282880 131096
rect 307760 131044 307812 131096
rect 231676 130976 231728 131028
rect 257344 130976 257396 131028
rect 282184 130976 282236 131028
rect 300952 130976 301004 131028
rect 231584 130908 231636 130960
rect 254768 130908 254820 130960
rect 210424 129820 210476 129872
rect 214012 129820 214064 129872
rect 261668 129820 261720 129872
rect 265072 129820 265124 129872
rect 174636 129752 174688 129804
rect 213920 129752 213972 129804
rect 254584 129752 254636 129804
rect 264980 129752 265032 129804
rect 231768 129684 231820 129736
rect 253480 129684 253532 129736
rect 231676 129616 231728 129668
rect 244924 129616 244976 129668
rect 231124 129072 231176 129124
rect 242440 129072 242492 129124
rect 231584 129004 231636 129056
rect 246304 129004 246356 129056
rect 204996 128392 205048 128444
rect 213920 128392 213972 128444
rect 257344 128392 257396 128444
rect 265072 128392 265124 128444
rect 59268 128324 59320 128376
rect 66168 128324 66220 128376
rect 170496 128324 170548 128376
rect 214012 128324 214064 128376
rect 246488 128324 246540 128376
rect 264980 128324 265032 128376
rect 230848 128256 230900 128308
rect 261760 128256 261812 128308
rect 281724 128256 281776 128308
rect 295432 128256 295484 128308
rect 231768 128188 231820 128240
rect 260288 128188 260340 128240
rect 282828 128188 282880 128240
rect 289912 128188 289964 128240
rect 231032 127576 231084 127628
rect 239588 127576 239640 127628
rect 253572 127576 253624 127628
rect 265716 127576 265768 127628
rect 202328 127032 202380 127084
rect 213920 127032 213972 127084
rect 174544 126964 174596 127016
rect 214012 126964 214064 127016
rect 261576 126964 261628 127016
rect 264980 126964 265032 127016
rect 231768 126896 231820 126948
rect 251824 126896 251876 126948
rect 281908 126896 281960 126948
rect 285680 126896 285732 126948
rect 231676 126828 231728 126880
rect 250720 126828 250772 126880
rect 257528 125740 257580 125792
rect 264980 125740 265032 125792
rect 193956 125672 194008 125724
rect 213920 125672 213972 125724
rect 254768 125672 254820 125724
rect 265072 125672 265124 125724
rect 167644 125604 167696 125656
rect 214012 125604 214064 125656
rect 236920 125604 236972 125656
rect 265164 125604 265216 125656
rect 231492 125536 231544 125588
rect 261484 125536 261536 125588
rect 282828 125536 282880 125588
rect 305184 125536 305236 125588
rect 231768 125468 231820 125520
rect 253296 125468 253348 125520
rect 282736 125468 282788 125520
rect 298192 125468 298244 125520
rect 231768 125060 231820 125112
rect 236828 125060 236880 125112
rect 230940 124584 230992 124636
rect 235540 124584 235592 124636
rect 252192 124312 252244 124364
rect 264980 124312 265032 124364
rect 195428 124244 195480 124296
rect 213920 124244 213972 124296
rect 239588 124244 239640 124296
rect 265072 124244 265124 124296
rect 178776 124176 178828 124228
rect 214012 124176 214064 124228
rect 235264 124176 235316 124228
rect 265164 124176 265216 124228
rect 230756 124108 230808 124160
rect 232504 124108 232556 124160
rect 282644 124108 282696 124160
rect 306380 124108 306432 124160
rect 282828 124040 282880 124092
rect 295524 124040 295576 124092
rect 230756 123564 230808 123616
rect 238024 123564 238076 123616
rect 282736 123428 282788 123480
rect 303620 123428 303672 123480
rect 250720 122952 250772 123004
rect 264980 122952 265032 123004
rect 173440 122884 173492 122936
rect 214012 122884 214064 122936
rect 232688 122884 232740 122936
rect 265072 122884 265124 122936
rect 171784 122816 171836 122868
rect 213920 122816 213972 122868
rect 229836 122816 229888 122868
rect 265164 122816 265216 122868
rect 231676 122748 231728 122800
rect 264244 122748 264296 122800
rect 282828 122748 282880 122800
rect 292580 122748 292632 122800
rect 231768 122680 231820 122732
rect 242348 122680 242400 122732
rect 231676 122068 231728 122120
rect 243728 122068 243780 122120
rect 256332 121592 256384 121644
rect 265072 121592 265124 121644
rect 206468 121524 206520 121576
rect 213920 121524 213972 121576
rect 246304 121524 246356 121576
rect 264980 121524 265032 121576
rect 63408 121456 63460 121508
rect 65984 121456 66036 121508
rect 203524 121456 203576 121508
rect 214012 121456 214064 121508
rect 243636 121456 243688 121508
rect 265164 121456 265216 121508
rect 231768 121388 231820 121440
rect 247868 121388 247920 121440
rect 281540 121320 281592 121372
rect 284392 121320 284444 121372
rect 231584 121252 231636 121304
rect 234160 121252 234212 121304
rect 230756 120708 230808 120760
rect 257620 120708 257672 120760
rect 242532 120232 242584 120284
rect 264980 120232 265032 120284
rect 207664 120164 207716 120216
rect 214012 120164 214064 120216
rect 238300 120164 238352 120216
rect 265164 120164 265216 120216
rect 62028 120096 62080 120148
rect 65892 120096 65944 120148
rect 196808 120096 196860 120148
rect 213920 120096 213972 120148
rect 232504 120096 232556 120148
rect 265072 120096 265124 120148
rect 230940 120028 230992 120080
rect 260104 120028 260156 120080
rect 282092 120028 282144 120080
rect 291292 120028 291344 120080
rect 231400 119960 231452 120012
rect 240876 119960 240928 120012
rect 209228 118804 209280 118856
rect 213920 118804 213972 118856
rect 193864 118736 193916 118788
rect 214104 118736 214156 118788
rect 192484 118668 192536 118720
rect 214012 118668 214064 118720
rect 231308 118668 231360 118720
rect 232780 118668 232832 118720
rect 258816 118668 258868 118720
rect 264980 118668 265032 118720
rect 231492 118600 231544 118652
rect 258908 118600 258960 118652
rect 282828 118600 282880 118652
rect 289820 118600 289872 118652
rect 231768 118532 231820 118584
rect 258724 118532 258776 118584
rect 282736 118532 282788 118584
rect 288716 118532 288768 118584
rect 231676 118396 231728 118448
rect 236736 118396 236788 118448
rect 189816 117376 189868 117428
rect 214012 117376 214064 117428
rect 261484 117376 261536 117428
rect 265072 117376 265124 117428
rect 171876 117308 171928 117360
rect 213920 117308 213972 117360
rect 247868 117308 247920 117360
rect 264980 117308 265032 117360
rect 231768 117240 231820 117292
rect 254860 117240 254912 117292
rect 282828 117240 282880 117292
rect 298284 117240 298336 117292
rect 282736 117172 282788 117224
rect 288532 117172 288584 117224
rect 230664 116968 230716 117020
rect 234068 116968 234120 117020
rect 234160 116560 234212 116612
rect 261852 116560 261904 116612
rect 253480 116152 253532 116204
rect 264980 116152 265032 116204
rect 260104 116084 260156 116136
rect 265164 116084 265216 116136
rect 258724 116016 258776 116068
rect 264980 116016 265032 116068
rect 181536 115948 181588 116000
rect 213920 115948 213972 116000
rect 262956 115948 263008 116000
rect 265072 115948 265124 116000
rect 231768 115880 231820 115932
rect 255964 115880 256016 115932
rect 281724 115880 281776 115932
rect 309140 115880 309192 115932
rect 231676 115812 231728 115864
rect 249340 115812 249392 115864
rect 282092 115812 282144 115864
rect 296720 115812 296772 115864
rect 231768 115268 231820 115320
rect 239680 115268 239732 115320
rect 230020 115200 230072 115252
rect 267280 115200 267332 115252
rect 185676 114588 185728 114640
rect 214012 114588 214064 114640
rect 177580 114520 177632 114572
rect 213920 114520 213972 114572
rect 249156 114520 249208 114572
rect 264980 114520 265032 114572
rect 231492 114452 231544 114504
rect 253388 114452 253440 114504
rect 282828 114452 282880 114504
rect 302332 114452 302384 114504
rect 282736 114384 282788 114436
rect 299572 114384 299624 114436
rect 230848 113772 230900 113824
rect 263048 113772 263100 113824
rect 200856 113228 200908 113280
rect 214012 113228 214064 113280
rect 196716 113160 196768 113212
rect 213920 113160 213972 113212
rect 231768 113092 231820 113144
rect 252008 113092 252060 113144
rect 282092 113092 282144 113144
rect 300860 113092 300912 113144
rect 231676 113024 231728 113076
rect 250628 113024 250680 113076
rect 258908 111936 258960 111988
rect 265164 111936 265216 111988
rect 211804 111868 211856 111920
rect 214012 111868 214064 111920
rect 251824 111868 251876 111920
rect 264980 111868 265032 111920
rect 169116 111800 169168 111852
rect 213920 111800 213972 111852
rect 244924 111800 244976 111852
rect 265072 111800 265124 111852
rect 3148 111732 3200 111784
rect 22744 111732 22796 111784
rect 167828 111732 167880 111784
rect 198004 111732 198056 111784
rect 231768 111732 231820 111784
rect 251916 111732 251968 111784
rect 282736 111732 282788 111784
rect 303712 111732 303764 111784
rect 230572 111664 230624 111716
rect 246580 111664 246632 111716
rect 282828 111664 282880 111716
rect 298100 111664 298152 111716
rect 231308 111052 231360 111104
rect 260472 111052 260524 111104
rect 260380 110576 260432 110628
rect 265164 110576 265216 110628
rect 178868 110508 178920 110560
rect 213920 110508 213972 110560
rect 256148 110508 256200 110560
rect 264980 110508 265032 110560
rect 177488 110440 177540 110492
rect 214012 110440 214064 110492
rect 236736 110440 236788 110492
rect 265072 110440 265124 110492
rect 167828 110372 167880 110424
rect 215300 110372 215352 110424
rect 231676 110372 231728 110424
rect 264428 110372 264480 110424
rect 282092 110372 282144 110424
rect 302240 110372 302292 110424
rect 230572 110304 230624 110356
rect 262864 110304 262916 110356
rect 282276 110304 282328 110356
rect 292672 110304 292724 110356
rect 231768 110236 231820 110288
rect 245108 110236 245160 110288
rect 260288 109148 260340 109200
rect 265164 109148 265216 109200
rect 198188 109080 198240 109132
rect 214012 109080 214064 109132
rect 253296 109080 253348 109132
rect 264980 109080 265032 109132
rect 166448 109012 166500 109064
rect 213920 109012 213972 109064
rect 238024 109012 238076 109064
rect 265072 109012 265124 109064
rect 167828 108944 167880 108996
rect 200764 108944 200816 108996
rect 231768 108944 231820 108996
rect 249064 108944 249116 108996
rect 281724 108944 281776 108996
rect 303804 108944 303856 108996
rect 282092 108876 282144 108928
rect 293960 108876 294012 108928
rect 231492 108604 231544 108656
rect 235448 108604 235500 108656
rect 231400 108264 231452 108316
rect 241060 108264 241112 108316
rect 241152 107856 241204 107908
rect 265072 107856 265124 107908
rect 246580 107788 246632 107840
rect 264980 107788 265032 107840
rect 191288 107720 191340 107772
rect 214012 107720 214064 107772
rect 243728 107720 243780 107772
rect 265164 107720 265216 107772
rect 167828 107652 167880 107704
rect 213920 107652 213972 107704
rect 231492 107584 231544 107636
rect 256056 107584 256108 107636
rect 231768 107516 231820 107568
rect 253204 107516 253256 107568
rect 169208 106904 169260 106956
rect 214656 106904 214708 106956
rect 231216 106904 231268 106956
rect 246396 106904 246448 106956
rect 242348 106428 242400 106480
rect 264980 106428 265032 106480
rect 199384 106360 199436 106412
rect 214012 106360 214064 106412
rect 249064 106360 249116 106412
rect 265072 106360 265124 106412
rect 182916 106292 182968 106344
rect 213920 106292 213972 106344
rect 231676 106224 231728 106276
rect 250812 106224 250864 106276
rect 281540 106224 281592 106276
rect 284484 106224 284536 106276
rect 231768 106156 231820 106208
rect 250536 106156 250588 106208
rect 230572 106088 230624 106140
rect 245200 106088 245252 106140
rect 259000 105000 259052 105052
rect 265072 105000 265124 105052
rect 184388 104932 184440 104984
rect 214012 104932 214064 104984
rect 263048 104932 263100 104984
rect 265440 104932 265492 104984
rect 180156 104864 180208 104916
rect 213920 104864 213972 104916
rect 250444 104864 250496 104916
rect 264980 104864 265032 104916
rect 282828 104796 282880 104848
rect 305092 104796 305144 104848
rect 230848 104728 230900 104780
rect 232596 104728 232648 104780
rect 231768 104660 231820 104712
rect 249248 104660 249300 104712
rect 230756 104184 230808 104236
rect 256240 104184 256292 104236
rect 235448 104116 235500 104168
rect 262956 104116 263008 104168
rect 231492 103844 231544 103896
rect 235356 103844 235408 103896
rect 256056 103640 256108 103692
rect 265072 103640 265124 103692
rect 253204 103572 253256 103624
rect 265164 103572 265216 103624
rect 170588 103504 170640 103556
rect 213920 103504 213972 103556
rect 249340 103504 249392 103556
rect 264980 103504 265032 103556
rect 231768 103436 231820 103488
rect 247776 103436 247828 103488
rect 282828 103436 282880 103488
rect 299480 103436 299532 103488
rect 231676 103368 231728 103420
rect 242164 103368 242216 103420
rect 231584 103300 231636 103352
rect 242256 103300 242308 103352
rect 240876 102348 240928 102400
rect 265072 102348 265124 102400
rect 255964 102280 256016 102332
rect 264980 102280 265032 102332
rect 242440 102212 242492 102264
rect 265164 102212 265216 102264
rect 195520 102144 195572 102196
rect 213920 102144 213972 102196
rect 262864 102144 262916 102196
rect 265256 102144 265308 102196
rect 231768 102076 231820 102128
rect 253572 102076 253624 102128
rect 231676 101396 231728 101448
rect 252100 101396 252152 101448
rect 261300 100852 261352 100904
rect 265072 100852 265124 100904
rect 262956 100784 263008 100836
rect 265348 100784 265400 100836
rect 176016 100716 176068 100768
rect 213920 100716 213972 100768
rect 249248 100716 249300 100768
rect 264980 100716 265032 100768
rect 231584 100648 231636 100700
rect 263140 100648 263192 100700
rect 281724 100648 281776 100700
rect 291384 100648 291436 100700
rect 231124 100580 231176 100632
rect 238208 100580 238260 100632
rect 230664 99968 230716 100020
rect 240968 99968 241020 100020
rect 169300 99424 169352 99476
rect 214012 99424 214064 99476
rect 250536 99424 250588 99476
rect 265072 99424 265124 99476
rect 166540 99356 166592 99408
rect 213920 99356 213972 99408
rect 242164 99356 242216 99408
rect 264980 99356 265032 99408
rect 231124 99288 231176 99340
rect 233884 99288 233936 99340
rect 282828 99288 282880 99340
rect 309232 99288 309284 99340
rect 203616 98064 203668 98116
rect 213920 98064 213972 98116
rect 245108 98064 245160 98116
rect 264980 98064 265032 98116
rect 164884 97996 164936 98048
rect 214012 97996 214064 98048
rect 231216 97996 231268 98048
rect 265072 97996 265124 98048
rect 282184 97928 282236 97980
rect 294144 97928 294196 97980
rect 282828 97860 282880 97912
rect 287152 97860 287204 97912
rect 229192 97248 229244 97300
rect 264980 97248 265032 97300
rect 206560 96908 206612 96960
rect 213920 96908 213972 96960
rect 196624 96840 196676 96892
rect 229192 96840 229244 96892
rect 234068 96840 234120 96892
rect 209320 96772 209372 96824
rect 214012 96772 214064 96824
rect 215944 96772 215996 96824
rect 264980 96772 265032 96824
rect 214656 96704 214708 96756
rect 265164 96704 265216 96756
rect 173164 96636 173216 96688
rect 265072 96636 265124 96688
rect 205548 96364 205600 96416
rect 279332 96364 279384 96416
rect 206284 96296 206336 96348
rect 279240 96296 279292 96348
rect 231124 95820 231176 95872
rect 233884 95820 233936 95872
rect 211896 95208 211948 95260
rect 214104 95208 214156 95260
rect 220176 95208 220228 95260
rect 264980 95208 265032 95260
rect 212448 95140 212500 95192
rect 229100 95140 229152 95192
rect 230664 95140 230716 95192
rect 225604 94732 225656 94784
rect 234160 94732 234212 94784
rect 221556 94664 221608 94716
rect 249340 94664 249392 94716
rect 228364 94596 228416 94648
rect 256332 94596 256384 94648
rect 224316 94528 224368 94580
rect 261300 94528 261352 94580
rect 222844 94460 222896 94512
rect 265716 94460 265768 94512
rect 267648 94460 267700 94512
rect 269120 94460 269172 94512
rect 151636 94120 151688 94172
rect 166264 94120 166316 94172
rect 110696 94052 110748 94104
rect 173348 94052 173400 94104
rect 119436 93984 119488 94036
rect 185584 93984 185636 94036
rect 109040 93916 109092 93968
rect 181536 93916 181588 93968
rect 115848 93848 115900 93900
rect 196808 93848 196860 93900
rect 213184 93780 213236 93832
rect 281816 93780 281868 93832
rect 230664 93712 230716 93764
rect 276940 93712 276992 93764
rect 234068 93644 234120 93696
rect 270960 93644 271012 93696
rect 151544 93440 151596 93492
rect 170404 93440 170456 93492
rect 152096 93372 152148 93424
rect 184296 93372 184348 93424
rect 125416 93304 125468 93356
rect 193956 93304 194008 93356
rect 213276 93304 213328 93356
rect 230020 93304 230072 93356
rect 100576 93236 100628 93288
rect 169116 93236 169168 93288
rect 204904 93236 204956 93288
rect 236920 93236 236972 93288
rect 105544 93168 105596 93220
rect 177580 93168 177632 93220
rect 195336 93168 195388 93220
rect 238300 93168 238352 93220
rect 118240 93100 118292 93152
rect 206468 93100 206520 93152
rect 226984 93100 227036 93152
rect 258908 93100 258960 93152
rect 230664 92556 230716 92608
rect 231216 92556 231268 92608
rect 109592 92420 109644 92472
rect 213368 92420 213420 92472
rect 113272 92352 113324 92404
rect 216036 92352 216088 92404
rect 123024 92284 123076 92336
rect 195428 92284 195480 92336
rect 115756 92216 115808 92268
rect 182824 92216 182876 92268
rect 105728 92148 105780 92200
rect 169208 92148 169260 92200
rect 125784 92080 125836 92132
rect 177304 92080 177356 92132
rect 200764 91944 200816 91996
rect 235448 91944 235500 91996
rect 206284 91876 206336 91928
rect 242532 91876 242584 91928
rect 216128 91808 216180 91860
rect 260380 91808 260432 91860
rect 218704 91740 218756 91792
rect 263048 91740 263100 91792
rect 85856 91128 85908 91180
rect 116584 91128 116636 91180
rect 74816 91060 74868 91112
rect 115204 91060 115256 91112
rect 104440 90992 104492 91044
rect 200856 90992 200908 91044
rect 91468 90924 91520 90976
rect 182916 90924 182968 90976
rect 99012 90856 99064 90908
rect 178868 90856 178920 90908
rect 106740 90788 106792 90840
rect 185676 90788 185728 90840
rect 121184 90720 121236 90772
rect 171784 90720 171836 90772
rect 136180 90652 136232 90704
rect 166356 90652 166408 90704
rect 220084 90448 220136 90500
rect 254676 90448 254728 90500
rect 187056 90380 187108 90432
rect 259000 90380 259052 90432
rect 177304 90312 177356 90364
rect 265808 90312 265860 90364
rect 101864 89632 101916 89684
rect 211804 89632 211856 89684
rect 97356 89564 97408 89616
rect 198188 89564 198240 89616
rect 117136 89496 117188 89548
rect 207664 89496 207716 89548
rect 86776 89428 86828 89480
rect 164884 89428 164936 89480
rect 110144 89360 110196 89412
rect 171876 89360 171928 89412
rect 126612 89292 126664 89344
rect 167644 89292 167696 89344
rect 198004 89088 198056 89140
rect 232688 89088 232740 89140
rect 217324 89020 217376 89072
rect 257436 89020 257488 89072
rect 202236 88952 202288 89004
rect 253480 88952 253532 89004
rect 107936 88272 107988 88324
rect 216220 88272 216272 88324
rect 102876 88204 102928 88256
rect 196716 88204 196768 88256
rect 113824 88136 113876 88188
rect 192484 88136 192536 88188
rect 94412 88068 94464 88120
rect 167828 88068 167880 88120
rect 96344 88000 96396 88052
rect 166448 88000 166500 88052
rect 124128 87932 124180 87984
rect 178776 87932 178828 87984
rect 209044 87728 209096 87780
rect 247868 87728 247920 87780
rect 221464 87660 221516 87712
rect 264520 87660 264572 87712
rect 191196 87592 191248 87644
rect 250720 87592 250772 87644
rect 112720 86912 112772 86964
rect 209228 86912 209280 86964
rect 89168 86844 89220 86896
rect 169300 86844 169352 86896
rect 111340 86776 111392 86828
rect 189816 86776 189868 86828
rect 100208 86708 100260 86760
rect 177488 86708 177540 86760
rect 112076 86640 112128 86692
rect 181444 86640 181496 86692
rect 121920 86572 121972 86624
rect 173440 86572 173492 86624
rect 184296 86232 184348 86284
rect 252192 86232 252244 86284
rect 3148 85484 3200 85536
rect 18604 85484 18656 85536
rect 93124 85484 93176 85536
rect 199384 85484 199436 85536
rect 97816 85416 97868 85468
rect 202328 85416 202380 85468
rect 119712 85348 119764 85400
rect 203524 85348 203576 85400
rect 88064 85280 88116 85332
rect 166540 85280 166592 85332
rect 115020 85212 115072 85264
rect 193864 85212 193916 85264
rect 98736 85144 98788 85196
rect 174544 85144 174596 85196
rect 211804 84804 211856 84856
rect 261668 84804 261720 84856
rect 102048 84124 102100 84176
rect 210424 84124 210476 84176
rect 95148 84056 95200 84108
rect 191288 84056 191340 84108
rect 114468 83988 114520 84040
rect 209136 83988 209188 84040
rect 101956 83920 102008 83972
rect 170496 83920 170548 83972
rect 132408 83852 132460 83904
rect 184204 83852 184256 83904
rect 37188 83444 37240 83496
rect 246488 83444 246540 83496
rect 67640 82764 67692 82816
rect 209320 82764 209372 82816
rect 99104 82696 99156 82748
rect 204996 82696 205048 82748
rect 122748 82628 122800 82680
rect 206376 82628 206428 82680
rect 121276 82560 121328 82612
rect 187148 82560 187200 82612
rect 151728 82492 151780 82544
rect 180064 82492 180116 82544
rect 106188 82084 106240 82136
rect 229836 82084 229888 82136
rect 63408 81336 63460 81388
rect 195520 81336 195572 81388
rect 129648 81268 129700 81320
rect 198096 81268 198148 81320
rect 108948 81200 109000 81252
rect 175924 81200 175976 81252
rect 113088 80724 113140 80776
rect 239588 80724 239640 80776
rect 79324 80656 79376 80708
rect 265624 80656 265676 80708
rect 66168 79976 66220 80028
rect 170588 79976 170640 80028
rect 128268 79908 128320 79960
rect 188344 79908 188396 79960
rect 124128 79432 124180 79484
rect 254768 79432 254820 79484
rect 108948 79364 109000 79416
rect 256148 79364 256200 79416
rect 71044 79296 71096 79348
rect 221556 79296 221608 79348
rect 67548 78616 67600 78668
rect 213460 78616 213512 78668
rect 135168 78548 135220 78600
rect 202144 78548 202196 78600
rect 126888 78480 126940 78532
rect 186964 78480 187016 78532
rect 102048 78004 102100 78056
rect 253296 78004 253348 78056
rect 50988 77936 51040 77988
rect 267188 77936 267240 77988
rect 107568 77188 107620 77240
rect 173256 77188 173308 77240
rect 131028 77120 131080 77172
rect 191104 77120 191156 77172
rect 125508 76644 125560 76696
rect 243544 76644 243596 76696
rect 73068 76576 73120 76628
rect 264428 76576 264480 76628
rect 30288 76508 30340 76560
rect 249248 76508 249300 76560
rect 115204 75828 115256 75880
rect 211896 75828 211948 75880
rect 133788 75760 133840 75812
rect 195244 75760 195296 75812
rect 91008 75216 91060 75268
rect 241152 75216 241204 75268
rect 34428 75148 34480 75200
rect 262956 75148 263008 75200
rect 116584 74468 116636 74520
rect 203616 74468 203668 74520
rect 95148 73992 95200 74044
rect 243728 73992 243780 74044
rect 75828 73924 75880 73976
rect 239496 73924 239548 73976
rect 41328 73856 41380 73908
rect 242440 73856 242492 73908
rect 15108 73788 15160 73840
rect 261576 73788 261628 73840
rect 574744 73108 574796 73160
rect 580172 73108 580224 73160
rect 115848 72564 115900 72616
rect 236736 72564 236788 72616
rect 89628 72496 89680 72548
rect 245016 72496 245068 72548
rect 70308 72428 70360 72480
rect 258816 72428 258868 72480
rect 3424 71680 3476 71732
rect 57244 71680 57296 71732
rect 65984 71680 66036 71732
rect 206560 71680 206612 71732
rect 122748 71068 122800 71120
rect 251824 71068 251876 71120
rect 86868 71000 86920 71052
rect 264336 71000 264388 71052
rect 107568 69776 107620 69828
rect 233976 69776 234028 69828
rect 111708 69708 111760 69760
rect 239404 69708 239456 69760
rect 68928 69640 68980 69692
rect 260196 69640 260248 69692
rect 117228 68348 117280 68400
rect 235264 68348 235316 68400
rect 88248 68280 88300 68332
rect 243636 68280 243688 68332
rect 77208 66852 77260 66904
rect 242348 66852 242400 66904
rect 84108 65492 84160 65544
rect 246580 65492 246632 65544
rect 47584 64200 47636 64252
rect 222936 64200 222988 64252
rect 35808 64132 35860 64184
rect 249156 64132 249208 64184
rect 97908 62840 97960 62892
rect 260288 62840 260340 62892
rect 53748 62772 53800 62824
rect 267096 62772 267148 62824
rect 93768 61344 93820 61396
rect 229744 61344 229796 61396
rect 3056 59304 3108 59356
rect 17224 59304 17276 59356
rect 119896 58692 119948 58744
rect 226984 58692 227036 58744
rect 86776 58624 86828 58676
rect 221464 58624 221516 58676
rect 17868 57196 17920 57248
rect 250536 57196 250588 57248
rect 111616 55904 111668 55956
rect 216128 55904 216180 55956
rect 44088 55836 44140 55888
rect 254584 55836 254636 55888
rect 39948 54476 40000 54528
rect 257344 54476 257396 54528
rect 27528 53116 27580 53168
rect 224316 53116 224368 53168
rect 26148 53048 26200 53100
rect 245108 53048 245160 53100
rect 55128 51756 55180 51808
rect 256056 51756 256108 51808
rect 5448 51688 5500 51740
rect 220176 51688 220228 51740
rect 104164 50328 104216 50380
rect 206284 50328 206336 50380
rect 3424 48968 3476 49020
rect 54484 48968 54536 49020
rect 65524 48968 65576 49020
rect 231124 48968 231176 49020
rect 58624 47608 58676 47660
rect 231216 47608 231268 47660
rect 13728 47540 13780 47592
rect 269120 47540 269172 47592
rect 70216 46180 70268 46232
rect 218704 46180 218756 46232
rect 2780 45500 2832 45552
rect 4804 45500 4856 45552
rect 92388 44888 92440 44940
rect 228364 44888 228416 44940
rect 71688 44820 71740 44872
rect 225604 44820 225656 44872
rect 42708 43392 42760 43444
rect 200764 43392 200816 43444
rect 110328 42100 110380 42152
rect 184296 42100 184348 42152
rect 38568 42032 38620 42084
rect 258724 42032 258776 42084
rect 99288 40672 99340 40724
rect 191196 40672 191248 40724
rect 12348 39312 12400 39364
rect 214656 39312 214708 39364
rect 103428 37952 103480 38004
rect 240784 37952 240836 38004
rect 45468 37884 45520 37936
rect 202236 37884 202288 37936
rect 100668 36524 100720 36576
rect 236644 36524 236696 36576
rect 82728 35232 82780 35284
rect 238116 35232 238168 35284
rect 10968 35164 11020 35216
rect 204904 35164 204956 35216
rect 78588 33736 78640 33788
rect 247684 33736 247736 33788
rect 96528 32444 96580 32496
rect 217324 32444 217376 32496
rect 62028 32376 62080 32428
rect 187056 32376 187108 32428
rect 114468 29656 114520 29708
rect 213276 29656 213328 29708
rect 4068 29588 4120 29640
rect 224224 29588 224276 29640
rect 81348 28296 81400 28348
rect 195336 28296 195388 28348
rect 24768 28228 24820 28280
rect 270592 28228 270644 28280
rect 118608 26936 118660 26988
rect 220084 26936 220136 26988
rect 53656 26868 53708 26920
rect 261484 26868 261536 26920
rect 3976 25508 4028 25560
rect 215944 25508 215996 25560
rect 46848 24080 46900 24132
rect 211804 24080 211856 24132
rect 37096 22720 37148 22772
rect 255964 22720 256016 22772
rect 56508 21360 56560 21412
rect 267004 21360 267056 21412
rect 112 19932 164 19984
rect 196624 19932 196676 19984
rect 9588 18572 9640 18624
rect 244924 18572 244976 18624
rect 49608 17212 49660 17264
rect 260104 17212 260156 17264
rect 66168 15852 66220 15904
rect 250444 15852 250496 15904
rect 59268 14424 59320 14476
rect 253204 14424 253256 14476
rect 60648 13064 60700 13116
rect 209044 13064 209096 13116
rect 85488 11772 85540 11824
rect 246304 11772 246356 11824
rect 3884 11704 3936 11756
rect 4068 11704 4120 11756
rect 47860 11704 47912 11756
rect 262864 11704 262916 11756
rect 79692 10276 79744 10328
rect 249064 10276 249116 10328
rect 104532 8916 104584 8968
rect 238024 8916 238076 8968
rect 44272 7624 44324 7676
rect 240876 7624 240928 7676
rect 12256 7556 12308 7608
rect 242164 7556 242216 7608
rect 3424 6808 3476 6860
rect 51724 6808 51776 6860
rect 102232 6196 102284 6248
rect 198004 6196 198056 6248
rect 60832 6128 60884 6180
rect 214564 6128 214616 6180
rect 73804 4836 73856 4888
rect 232504 4836 232556 4888
rect 6460 4768 6512 4820
rect 173164 4768 173216 4820
rect 51356 3680 51408 3732
rect 71044 3680 71096 3732
rect 35992 3612 36044 3664
rect 37096 3612 37148 3664
rect 11152 3544 11204 3596
rect 12348 3544 12400 3596
rect 19432 3544 19484 3596
rect 47584 3544 47636 3596
rect 48964 3544 49016 3596
rect 49608 3544 49660 3596
rect 50160 3544 50212 3596
rect 50988 3544 51040 3596
rect 52552 3544 52604 3596
rect 53656 3544 53708 3596
rect 2872 3476 2924 3528
rect 3884 3476 3936 3528
rect 58624 3612 58676 3664
rect 85672 3612 85724 3664
rect 86776 3612 86828 3664
rect 1676 3408 1728 3460
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 64328 3476 64380 3528
rect 79324 3544 79376 3596
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 77392 3476 77444 3528
rect 104164 3544 104216 3596
rect 105728 3544 105780 3596
rect 106188 3544 106240 3596
rect 106924 3544 106976 3596
rect 107568 3544 107620 3596
rect 108120 3544 108172 3596
rect 108948 3544 109000 3596
rect 109316 3544 109368 3596
rect 110328 3544 110380 3596
rect 114008 3544 114060 3596
rect 114468 3544 114520 3596
rect 115204 3544 115256 3596
rect 115848 3544 115900 3596
rect 116400 3544 116452 3596
rect 117228 3544 117280 3596
rect 117596 3544 117648 3596
rect 118608 3544 118660 3596
rect 118792 3544 118844 3596
rect 119804 3544 119856 3596
rect 122288 3544 122340 3596
rect 122748 3544 122800 3596
rect 123484 3544 123536 3596
rect 124128 3544 124180 3596
rect 124680 3544 124732 3596
rect 125508 3544 125560 3596
rect 125876 3544 125928 3596
rect 178684 3544 178736 3596
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 93952 3476 94004 3528
rect 95148 3476 95200 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 8760 3408 8812 3460
rect 9588 3408 9640 3460
rect 9956 3408 10008 3460
rect 10968 3408 11020 3460
rect 15936 3408 15988 3460
rect 16488 3408 16540 3460
rect 17040 3408 17092 3460
rect 17868 3408 17920 3460
rect 18236 3408 18288 3460
rect 19248 3408 19300 3460
rect 24216 3408 24268 3460
rect 24768 3408 24820 3460
rect 25320 3408 25372 3460
rect 26148 3408 26200 3460
rect 26516 3408 26568 3460
rect 27528 3408 27580 3460
rect 32404 3408 32456 3460
rect 33048 3408 33100 3460
rect 33600 3408 33652 3460
rect 34428 3408 34480 3460
rect 27712 3340 27764 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 41880 3340 41932 3392
rect 42708 3340 42760 3392
rect 43076 3340 43128 3392
rect 44088 3340 44140 3392
rect 84476 3408 84528 3460
rect 85488 3408 85540 3460
rect 95148 3340 95200 3392
rect 222844 3476 222896 3528
rect 177304 3408 177356 3460
rect 101036 3136 101088 3188
rect 102048 3136 102100 3188
rect 110512 3136 110564 3188
rect 111708 3136 111760 3188
rect 233884 3000 233936 3052
rect 235816 3000 235868 3052
rect 92756 2864 92808 2916
rect 93768 2864 93820 2916
rect 7656 2116 7708 2168
rect 65432 2116 65484 2168
rect 63224 2048 63276 2100
rect 264244 2048 264296 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 619168 2834 619177
rect 2778 619103 2780 619112
rect 2832 619103 2834 619112
rect 2780 619074 2832 619080
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3436 463010 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 4804 619132 4856 619138
rect 4804 619074 4856 619080
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3424 463004 3476 463010
rect 3424 462946 3476 462952
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305046 3464 306167
rect 3424 305040 3476 305046
rect 3424 304982 3476 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 20 290148 72 290154
rect 20 290090 72 290096
rect 32 19961 60 290090
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3528 257378 3556 462567
rect 4816 276010 4844 619074
rect 4804 276004 4856 276010
rect 4804 275946 4856 275952
rect 8220 273970 8248 702406
rect 24320 700330 24348 703520
rect 40512 700466 40540 703520
rect 72988 702434 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72988 702406 73108 702434
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 35164 553444 35216 553450
rect 35164 553386 35216 553392
rect 21364 422340 21416 422346
rect 21364 422282 21416 422288
rect 21376 382974 21404 422282
rect 29644 409896 29696 409902
rect 29644 409838 29696 409844
rect 21364 382968 21416 382974
rect 21364 382910 21416 382916
rect 21364 371272 21416 371278
rect 21364 371214 21416 371220
rect 15844 357468 15896 357474
rect 15844 357410 15896 357416
rect 15856 338774 15884 357410
rect 15844 338768 15896 338774
rect 15844 338710 15896 338716
rect 11704 292596 11756 292602
rect 11704 292538 11756 292544
rect 8208 273964 8260 273970
rect 8208 273906 8260 273912
rect 3516 257372 3568 257378
rect 3516 257314 3568 257320
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 242214 3464 254079
rect 11716 244254 11744 292538
rect 17224 284368 17276 284374
rect 17224 284310 17276 284316
rect 15844 264988 15896 264994
rect 15844 264930 15896 264936
rect 11704 244248 11756 244254
rect 11704 244190 11756 244196
rect 3424 242208 3476 242214
rect 3424 242150 3476 242156
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240174 3464 241023
rect 3424 240168 3476 240174
rect 3424 240110 3476 240116
rect 3424 233912 3476 233918
rect 3424 233854 3476 233860
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 97617 3464 233854
rect 4804 232552 4856 232558
rect 4804 232494 4856 232500
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 49020 3476 49026
rect 3424 48962 3476 48968
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 2832 45520 2834 45529
rect 2778 45455 2834 45464
rect 3436 32473 3464 48962
rect 4816 45558 4844 232494
rect 15856 215286 15884 264930
rect 15844 215280 15896 215286
rect 15844 215222 15896 215228
rect 15108 73840 15160 73846
rect 15108 73782 15160 73788
rect 5448 51740 5500 51746
rect 5448 51682 5500 51688
rect 4804 45552 4856 45558
rect 4804 45494 4856 45500
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 3976 25560 4028 25566
rect 3976 25502 4028 25508
rect 112 19984 164 19990
rect 18 19952 74 19961
rect 112 19926 164 19932
rect 18 19887 74 19896
rect 124 16574 152 19926
rect 124 16546 612 16574
rect 584 480 612 16546
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3896 3534 3924 11698
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3470
rect 3988 1578 4016 25502
rect 4080 11762 4108 29582
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 5460 6914 5488 51682
rect 13728 47592 13780 47598
rect 13728 47534 13780 47540
rect 12348 39364 12400 39370
rect 12348 39306 12400 39312
rect 10968 35216 11020 35222
rect 10968 35158 11020 35164
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 5276 6886 5488 6914
rect 3988 1550 4108 1578
rect 4080 480 4108 1550
rect 5276 480 5304 6886
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6472 480 6500 4762
rect 9600 3466 9628 18566
rect 10980 3466 11008 35158
rect 12256 7608 12308 7614
rect 12256 7550 12308 7556
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 7656 2168 7708 2174
rect 7656 2110 7708 2116
rect 7668 480 7696 2110
rect 8772 480 8800 3402
rect 9968 480 9996 3402
rect 11164 480 11192 3538
rect 12268 3482 12296 7550
rect 12360 3602 12388 39306
rect 13740 6914 13768 47534
rect 15120 6914 15148 73782
rect 17236 59362 17264 284310
rect 18604 253972 18656 253978
rect 18604 253914 18656 253920
rect 18616 85542 18644 253914
rect 21376 238474 21404 371214
rect 29656 247042 29684 409838
rect 35176 264926 35204 553386
rect 35164 264920 35216 264926
rect 35164 264862 35216 264868
rect 32404 258120 32456 258126
rect 32404 258062 32456 258068
rect 29644 247036 29696 247042
rect 29644 246978 29696 246984
rect 21364 238468 21416 238474
rect 21364 238410 21416 238416
rect 22744 235340 22796 235346
rect 22744 235282 22796 235288
rect 22756 111790 22784 235282
rect 32416 137970 32444 258062
rect 41340 237386 41368 700402
rect 73080 665854 73108 702406
rect 73068 665848 73120 665854
rect 73068 665790 73120 665796
rect 68284 565888 68336 565894
rect 68284 565830 68336 565836
rect 57244 287292 57296 287298
rect 57244 287234 57296 287240
rect 43444 285932 43496 285938
rect 43444 285874 43496 285880
rect 41328 237380 41380 237386
rect 41328 237322 41380 237328
rect 43456 150414 43484 285874
rect 51724 281580 51776 281586
rect 51724 281522 51776 281528
rect 43444 150408 43496 150414
rect 43444 150350 43496 150356
rect 32404 137964 32456 137970
rect 32404 137906 32456 137912
rect 22744 111784 22796 111790
rect 22744 111726 22796 111732
rect 18604 85536 18656 85542
rect 18604 85478 18656 85484
rect 37188 83496 37240 83502
rect 37188 83438 37240 83444
rect 30288 76560 30340 76566
rect 30288 76502 30340 76508
rect 19246 66872 19302 66881
rect 19246 66807 19302 66816
rect 17224 59356 17276 59362
rect 17224 59298 17276 59304
rect 17868 57248 17920 57254
rect 17868 57190 17920 57196
rect 16486 50280 16542 50289
rect 16486 50215 16542 50224
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12268 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3466 16528 50215
rect 17880 3466 17908 57190
rect 19260 3466 19288 66807
rect 23386 65512 23442 65521
rect 23386 65447 23442 65456
rect 22006 59936 22062 59945
rect 22006 59871 22062 59880
rect 20626 21312 20682 21321
rect 20626 21247 20682 21256
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 15948 480 15976 3402
rect 17052 480 17080 3402
rect 18248 480 18276 3402
rect 19444 480 19472 3538
rect 20640 480 20668 21247
rect 22020 6914 22048 59871
rect 23400 6914 23428 65447
rect 27528 53168 27580 53174
rect 27528 53110 27580 53116
rect 26148 53100 26200 53106
rect 26148 53042 26200 53048
rect 24768 28280 24820 28286
rect 24768 28222 24820 28228
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3466 24808 28222
rect 26160 3466 26188 53042
rect 27540 3466 27568 53110
rect 28906 24168 28962 24177
rect 28906 24103 28962 24112
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3402
rect 26528 480 26556 3402
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27724 480 27752 3334
rect 28920 480 28948 24103
rect 30300 6914 30328 76502
rect 34428 75200 34480 75206
rect 34428 75142 34480 75148
rect 33046 57216 33102 57225
rect 33046 57151 33102 57160
rect 31666 30968 31722 30977
rect 31666 30903 31722 30912
rect 31680 6914 31708 30903
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3466 33088 57151
rect 34440 3466 34468 75142
rect 35808 64184 35860 64190
rect 35808 64126 35860 64132
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 32416 480 32444 3402
rect 33612 480 33640 3402
rect 35820 3398 35848 64126
rect 37096 22772 37148 22778
rect 37096 22714 37148 22720
rect 37108 16574 37136 22714
rect 37016 16546 37136 16574
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34808 480 34836 3334
rect 36004 480 36032 3606
rect 37016 3482 37044 16546
rect 37200 6914 37228 83438
rect 50988 77988 51040 77994
rect 50988 77930 51040 77936
rect 41328 73908 41380 73914
rect 41328 73850 41380 73856
rect 39948 54528 40000 54534
rect 39948 54470 40000 54476
rect 38568 42084 38620 42090
rect 38568 42026 38620 42032
rect 38580 6914 38608 42026
rect 39960 6914 39988 54470
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37108 3670 37136 6886
rect 37096 3664 37148 3670
rect 37096 3606 37148 3612
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3398 41368 73850
rect 47584 64252 47636 64258
rect 47584 64194 47636 64200
rect 44088 55888 44140 55894
rect 44088 55830 44140 55836
rect 42708 43444 42760 43450
rect 42708 43386 42760 43392
rect 42720 3398 42748 43386
rect 44100 3398 44128 55830
rect 45468 37936 45520 37942
rect 45468 37878 45520 37884
rect 44272 7676 44324 7682
rect 44272 7618 44324 7624
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3334
rect 43088 480 43116 3334
rect 44284 480 44312 7618
rect 45480 480 45508 37878
rect 46848 24132 46900 24138
rect 46848 24074 46900 24080
rect 46860 6914 46888 24074
rect 46676 6886 46888 6914
rect 46676 480 46704 6886
rect 47596 3602 47624 64194
rect 49608 17264 49660 17270
rect 49608 17206 49660 17212
rect 47860 11756 47912 11762
rect 47860 11698 47912 11704
rect 47584 3596 47636 3602
rect 47584 3538 47636 3544
rect 47872 480 47900 11698
rect 49620 3602 49648 17206
rect 51000 3602 51028 77930
rect 51736 6866 51764 281522
rect 54484 269136 54536 269142
rect 54484 269078 54536 269084
rect 53748 62824 53800 62830
rect 53748 62766 53800 62772
rect 53656 26920 53708 26926
rect 53656 26862 53708 26868
rect 51724 6860 51776 6866
rect 51724 6802 51776 6808
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 49608 3596 49660 3602
rect 49608 3538 49660 3544
rect 50160 3596 50212 3602
rect 50160 3538 50212 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 48976 480 49004 3538
rect 50172 480 50200 3538
rect 51368 480 51396 3674
rect 53668 3602 53696 26862
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 53656 3596 53708 3602
rect 53656 3538 53708 3544
rect 52564 480 52592 3538
rect 53760 480 53788 62766
rect 54496 49026 54524 269078
rect 57256 71738 57284 287234
rect 65524 284436 65576 284442
rect 65524 284378 65576 284384
rect 65536 164218 65564 284378
rect 68296 269074 68324 565830
rect 71044 527196 71096 527202
rect 71044 527138 71096 527144
rect 68284 269068 68336 269074
rect 68284 269010 68336 269016
rect 71056 262206 71084 527138
rect 89640 290562 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 699718 105492 703520
rect 137848 702434 137876 703520
rect 137848 702406 137968 702434
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 89628 290556 89680 290562
rect 89628 290498 89680 290504
rect 71044 262200 71096 262206
rect 71044 262142 71096 262148
rect 106200 239426 106228 699654
rect 112444 656940 112496 656946
rect 112444 656882 112496 656888
rect 112456 291922 112484 656882
rect 112444 291916 112496 291922
rect 112444 291858 112496 291864
rect 137940 254590 137968 702406
rect 154132 700126 154160 703520
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 155224 700120 155276 700126
rect 155224 700062 155276 700068
rect 155236 289134 155264 700062
rect 170324 699718 170352 703520
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 166264 632120 166316 632126
rect 166264 632062 166316 632068
rect 162124 514820 162176 514826
rect 162124 514762 162176 514768
rect 155224 289128 155276 289134
rect 155224 289070 155276 289076
rect 137928 254584 137980 254590
rect 137928 254526 137980 254532
rect 147680 254584 147732 254590
rect 147680 254526 147732 254532
rect 147692 251190 147720 254526
rect 147680 251184 147732 251190
rect 147680 251126 147732 251132
rect 162136 239902 162164 514762
rect 166276 267714 166304 632062
rect 171060 273222 171088 699654
rect 180708 697604 180760 697610
rect 180708 697546 180760 697552
rect 177304 397520 177356 397526
rect 177304 397462 177356 397468
rect 173164 284504 173216 284510
rect 173164 284446 173216 284452
rect 171048 273216 171100 273222
rect 171048 273158 171100 273164
rect 166264 267708 166316 267714
rect 166264 267650 166316 267656
rect 170404 266416 170456 266422
rect 170404 266358 170456 266364
rect 170416 240038 170444 266358
rect 170404 240032 170456 240038
rect 170404 239974 170456 239980
rect 162124 239896 162176 239902
rect 162124 239838 162176 239844
rect 106188 239420 106240 239426
rect 106188 239362 106240 239368
rect 170404 233980 170456 233986
rect 170404 233922 170456 233928
rect 170416 202842 170444 233922
rect 170404 202836 170456 202842
rect 170404 202778 170456 202784
rect 173176 189038 173204 284446
rect 177316 238610 177344 397462
rect 178040 273964 178092 273970
rect 178040 273906 178092 273912
rect 178052 269006 178080 273906
rect 178040 269000 178092 269006
rect 178040 268942 178092 268948
rect 178684 257372 178736 257378
rect 178684 257314 178736 257320
rect 177304 238604 177356 238610
rect 177304 238546 177356 238552
rect 178696 238513 178724 257314
rect 180616 252612 180668 252618
rect 180616 252554 180668 252560
rect 180064 242208 180116 242214
rect 180064 242150 180116 242156
rect 180076 238678 180104 242150
rect 180064 238672 180116 238678
rect 180064 238614 180116 238620
rect 178682 238504 178738 238513
rect 178682 238439 178738 238448
rect 178684 229900 178736 229906
rect 178684 229842 178736 229848
rect 173164 189032 173216 189038
rect 173164 188974 173216 188980
rect 130936 181076 130988 181082
rect 130936 181018 130988 181024
rect 173256 181076 173308 181082
rect 173256 181018 173308 181024
rect 128176 181008 128228 181014
rect 128176 180950 128228 180956
rect 102048 180940 102100 180946
rect 102048 180882 102100 180888
rect 99472 180872 99524 180878
rect 99472 180814 99524 180820
rect 99484 176769 99512 180814
rect 102060 177585 102088 180882
rect 123300 179716 123352 179722
rect 123300 179658 123352 179664
rect 121276 179648 121328 179654
rect 121276 179590 121328 179596
rect 110696 179580 110748 179586
rect 110696 179522 110748 179528
rect 108120 179512 108172 179518
rect 108120 179454 108172 179460
rect 102046 177576 102102 177585
rect 102046 177511 102102 177520
rect 105728 177132 105780 177138
rect 105728 177074 105780 177080
rect 105740 176769 105768 177074
rect 107016 176792 107068 176798
rect 99470 176760 99526 176769
rect 99470 176695 99526 176704
rect 105726 176760 105782 176769
rect 105726 176695 105782 176704
rect 107014 176760 107016 176769
rect 108132 176769 108160 179454
rect 109592 178152 109644 178158
rect 109592 178094 109644 178100
rect 109604 176769 109632 178094
rect 110708 176769 110736 179522
rect 114560 179444 114612 179450
rect 114560 179386 114612 179392
rect 112260 178356 112312 178362
rect 112260 178298 112312 178304
rect 112272 176769 112300 178298
rect 107068 176760 107070 176769
rect 107014 176695 107070 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 109590 176760 109646 176769
rect 109590 176695 109646 176704
rect 110694 176760 110750 176769
rect 110694 176695 110750 176704
rect 112258 176760 112314 176769
rect 112258 176695 112314 176704
rect 114466 176760 114522 176769
rect 114572 176746 114600 179386
rect 116952 178288 117004 178294
rect 116952 178230 117004 178236
rect 116964 176769 116992 178230
rect 119528 178084 119580 178090
rect 119528 178026 119580 178032
rect 119540 176769 119568 178026
rect 121288 177313 121316 179590
rect 123312 177313 123340 179658
rect 125968 178220 126020 178226
rect 125968 178162 126020 178168
rect 121274 177304 121330 177313
rect 121274 177239 121330 177248
rect 123298 177304 123354 177313
rect 123298 177239 123354 177248
rect 125980 176769 126008 178162
rect 127164 176996 127216 177002
rect 127164 176938 127216 176944
rect 127176 176769 127204 176938
rect 128188 176769 128216 180950
rect 129464 179784 129516 179790
rect 129464 179726 129516 179732
rect 129476 177313 129504 179726
rect 130948 177585 130976 181018
rect 169024 180940 169076 180946
rect 169024 180882 169076 180888
rect 168380 179784 168432 179790
rect 168380 179726 168432 179732
rect 132408 178424 132460 178430
rect 132408 178366 132460 178372
rect 165344 178424 165396 178430
rect 165344 178366 165396 178372
rect 130934 177576 130990 177585
rect 130934 177511 130990 177520
rect 129462 177304 129518 177313
rect 129462 177239 129518 177248
rect 132420 176769 132448 178366
rect 134432 177064 134484 177070
rect 134432 177006 134484 177012
rect 134444 176769 134472 177006
rect 158904 176928 158956 176934
rect 158904 176870 158956 176876
rect 148232 176860 148284 176866
rect 148232 176802 148284 176808
rect 148244 176769 148272 176802
rect 158916 176769 158944 176870
rect 114522 176718 114600 176746
rect 116950 176760 117006 176769
rect 114466 176695 114522 176704
rect 116950 176695 117006 176704
rect 119526 176760 119582 176769
rect 119526 176695 119582 176704
rect 125966 176760 126022 176769
rect 125966 176695 126022 176704
rect 127162 176760 127218 176769
rect 127162 176695 127218 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 132406 176760 132462 176769
rect 132406 176695 132462 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 136086 176760 136142 176769
rect 136086 176695 136088 176704
rect 136140 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158902 176760 158958 176769
rect 158902 176695 158958 176704
rect 136088 176666 136140 176672
rect 133144 176248 133196 176254
rect 133144 176190 133196 176196
rect 124496 176180 124548 176186
rect 124496 176122 124548 176128
rect 121920 176112 121972 176118
rect 121920 176054 121972 176060
rect 118424 176044 118476 176050
rect 118424 175986 118476 175992
rect 115756 175976 115808 175982
rect 115756 175918 115808 175924
rect 115768 175001 115796 175918
rect 118436 175545 118464 175986
rect 121932 175545 121960 176054
rect 124508 175681 124536 176122
rect 133156 175681 133184 176190
rect 124494 175672 124550 175681
rect 124494 175607 124550 175616
rect 133142 175672 133198 175681
rect 133142 175607 133198 175616
rect 118422 175536 118478 175545
rect 118422 175471 118478 175480
rect 121918 175536 121974 175545
rect 121918 175471 121974 175480
rect 115754 174992 115810 175001
rect 115754 174927 115810 174936
rect 165356 173874 165384 178366
rect 166356 178356 166408 178362
rect 166356 178298 166408 178304
rect 165436 177064 165488 177070
rect 165436 177006 165488 177012
rect 165448 175234 165476 177006
rect 165528 176248 165580 176254
rect 165528 176190 165580 176196
rect 165436 175228 165488 175234
rect 165436 175170 165488 175176
rect 165540 175166 165568 176190
rect 166262 175400 166318 175409
rect 166262 175335 166318 175344
rect 165528 175160 165580 175166
rect 165528 175102 165580 175108
rect 165344 173868 165396 173874
rect 165344 173810 165396 173816
rect 65524 164212 65576 164218
rect 65524 164154 65576 164160
rect 166276 155922 166304 175335
rect 166368 164218 166396 178298
rect 167642 177032 167698 177041
rect 167642 176967 167698 176976
rect 167736 176996 167788 177002
rect 166448 176180 166500 176186
rect 166448 176122 166500 176128
rect 166460 169726 166488 176122
rect 166448 169720 166500 169726
rect 166448 169662 166500 169668
rect 166356 164212 166408 164218
rect 166356 164154 166408 164160
rect 167656 158710 167684 176967
rect 167736 176938 167788 176944
rect 167748 171086 167776 176938
rect 168392 172514 168420 179726
rect 168380 172508 168432 172514
rect 168380 172450 168432 172456
rect 167918 171592 167974 171601
rect 167918 171527 167974 171536
rect 167932 171154 167960 171527
rect 167920 171148 167972 171154
rect 167920 171090 167972 171096
rect 167736 171080 167788 171086
rect 167736 171022 167788 171028
rect 167644 158704 167696 158710
rect 167644 158646 167696 158652
rect 169036 158642 169064 180882
rect 170402 176896 170458 176905
rect 170402 176831 170458 176840
rect 169116 176112 169168 176118
rect 169116 176054 169168 176060
rect 169128 168366 169156 176054
rect 169116 168360 169168 168366
rect 169116 168302 169168 168308
rect 170416 160070 170444 176831
rect 170496 176792 170548 176798
rect 170496 176734 170548 176740
rect 170508 161430 170536 176734
rect 173164 176044 173216 176050
rect 173164 175986 173216 175992
rect 171782 175536 171838 175545
rect 171782 175471 171838 175480
rect 171796 165578 171824 175471
rect 173176 167006 173204 175986
rect 173268 173806 173296 181018
rect 175924 179716 175976 179722
rect 175924 179658 175976 179664
rect 174544 178288 174596 178294
rect 174544 178230 174596 178236
rect 173256 173800 173308 173806
rect 173256 173742 173308 173748
rect 173164 167000 173216 167006
rect 173164 166942 173216 166948
rect 174556 166938 174584 178230
rect 175936 169658 175964 179658
rect 177396 179648 177448 179654
rect 177396 179590 177448 179596
rect 177302 178120 177358 178129
rect 177302 178055 177358 178064
rect 175924 169652 175976 169658
rect 175924 169594 175976 169600
rect 174544 166932 174596 166938
rect 174544 166874 174596 166880
rect 171784 165572 171836 165578
rect 171784 165514 171836 165520
rect 170496 161424 170548 161430
rect 170496 161366 170548 161372
rect 170404 160064 170456 160070
rect 170404 160006 170456 160012
rect 169024 158636 169076 158642
rect 169024 158578 169076 158584
rect 166264 155916 166316 155922
rect 166264 155858 166316 155864
rect 177316 155854 177344 178055
rect 177408 168298 177436 179590
rect 177396 168292 177448 168298
rect 177396 168234 177448 168240
rect 177304 155848 177356 155854
rect 177304 155790 177356 155796
rect 166264 153264 166316 153270
rect 166264 153206 166316 153212
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 66180 128382 66208 129231
rect 59268 128376 59320 128382
rect 59268 128318 59320 128324
rect 66168 128376 66220 128382
rect 66168 128318 66220 128324
rect 59280 95033 59308 128318
rect 66074 128072 66130 128081
rect 66074 128007 66130 128016
rect 65982 122632 66038 122641
rect 65982 122567 66038 122576
rect 65996 121514 66024 122567
rect 63408 121508 63460 121514
rect 63408 121450 63460 121456
rect 65984 121508 66036 121514
rect 65984 121450 66036 121456
rect 62028 120148 62080 120154
rect 62028 120090 62080 120096
rect 59266 95024 59322 95033
rect 59266 94959 59322 94968
rect 62040 86873 62068 120090
rect 62026 86864 62082 86873
rect 62026 86799 62082 86808
rect 63420 81394 63448 121450
rect 65890 120864 65946 120873
rect 65890 120799 65946 120808
rect 65904 120154 65932 120799
rect 65892 120148 65944 120154
rect 65892 120090 65944 120096
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 63408 81388 63460 81394
rect 63408 81330 63460 81336
rect 65996 71738 66024 102303
rect 66088 93809 66116 128007
rect 67454 126304 67510 126313
rect 67454 126239 67510 126248
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 93800 66130 93809
rect 66074 93735 66130 93744
rect 66180 80034 66208 125151
rect 67468 91089 67496 126239
rect 67546 123584 67602 123593
rect 67546 123519 67602 123528
rect 67454 91080 67510 91089
rect 67454 91015 67510 91024
rect 66168 80028 66220 80034
rect 66168 79970 66220 79976
rect 67560 78674 67588 123519
rect 67638 100736 67694 100745
rect 67638 100671 67694 100680
rect 67652 82822 67680 100671
rect 164884 98048 164936 98054
rect 164884 97990 164936 97996
rect 151634 94888 151690 94897
rect 151634 94823 151690 94832
rect 109038 94752 109094 94761
rect 109038 94687 109094 94696
rect 110694 94752 110750 94761
rect 110694 94687 110750 94696
rect 115846 94752 115902 94761
rect 115846 94687 115902 94696
rect 119434 94752 119490 94761
rect 119434 94687 119490 94696
rect 109052 93974 109080 94687
rect 110708 94110 110736 94687
rect 110696 94104 110748 94110
rect 110696 94046 110748 94052
rect 109040 93968 109092 93974
rect 109040 93910 109092 93916
rect 115860 93906 115888 94687
rect 119448 94042 119476 94687
rect 151648 94178 151676 94823
rect 151636 94172 151688 94178
rect 151636 94114 151688 94120
rect 119436 94036 119488 94042
rect 119436 93978 119488 93984
rect 115848 93900 115900 93906
rect 115848 93842 115900 93848
rect 100574 93528 100630 93537
rect 100574 93463 100630 93472
rect 105542 93528 105598 93537
rect 105542 93463 105598 93472
rect 118238 93528 118294 93537
rect 118238 93463 118294 93472
rect 125414 93528 125470 93537
rect 125414 93463 125470 93472
rect 151542 93528 151598 93537
rect 151542 93463 151544 93472
rect 100588 93294 100616 93463
rect 100576 93288 100628 93294
rect 100576 93230 100628 93236
rect 105556 93226 105584 93463
rect 110142 93256 110198 93265
rect 105544 93220 105596 93226
rect 110142 93191 110198 93200
rect 113822 93256 113878 93265
rect 113822 93191 113878 93200
rect 105544 93162 105596 93168
rect 109592 92472 109644 92478
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 85854 92440 85910 92449
rect 85854 92375 85910 92384
rect 91466 92440 91522 92449
rect 91466 92375 91522 92384
rect 99010 92440 99066 92449
rect 99010 92375 99066 92384
rect 104438 92440 104494 92449
rect 104438 92375 104494 92384
rect 105726 92440 105782 92449
rect 105726 92375 105782 92384
rect 106738 92440 106794 92449
rect 106738 92375 106794 92384
rect 109590 92440 109592 92449
rect 109644 92440 109646 92449
rect 109590 92375 109646 92384
rect 74828 91118 74856 92375
rect 85026 91760 85082 91769
rect 85026 91695 85082 91704
rect 74816 91112 74868 91118
rect 74816 91054 74868 91060
rect 85040 89593 85068 91695
rect 85868 91186 85896 92375
rect 91006 91896 91062 91905
rect 91006 91831 91062 91840
rect 86774 91624 86830 91633
rect 86774 91559 86830 91568
rect 85856 91180 85908 91186
rect 85856 91122 85908 91128
rect 85026 89584 85082 89593
rect 85026 89519 85082 89528
rect 86788 89486 86816 91559
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 89166 91216 89222 91225
rect 89166 91151 89222 91160
rect 86776 89480 86828 89486
rect 86776 89422 86828 89428
rect 88076 85338 88104 91151
rect 89180 86902 89208 91151
rect 91020 89729 91048 91831
rect 91480 90982 91508 92375
rect 97354 91760 97410 91769
rect 97354 91695 97410 91704
rect 93122 91216 93178 91225
rect 93122 91151 93178 91160
rect 94410 91216 94466 91225
rect 94410 91151 94466 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96342 91216 96398 91225
rect 96342 91151 96398 91160
rect 91468 90976 91520 90982
rect 91468 90918 91520 90924
rect 91006 89720 91062 89729
rect 91006 89655 91062 89664
rect 89168 86896 89220 86902
rect 89168 86838 89220 86844
rect 93136 85542 93164 91151
rect 94424 88126 94452 91151
rect 94412 88120 94464 88126
rect 94412 88062 94464 88068
rect 93124 85536 93176 85542
rect 93124 85478 93176 85484
rect 88064 85332 88116 85338
rect 88064 85274 88116 85280
rect 95160 84114 95188 91151
rect 96356 88058 96384 91151
rect 97368 89622 97396 91695
rect 97814 91216 97870 91225
rect 97814 91151 97870 91160
rect 98734 91216 98790 91225
rect 98734 91151 98790 91160
rect 97356 89616 97408 89622
rect 97356 89558 97408 89564
rect 96344 88052 96396 88058
rect 96344 87994 96396 88000
rect 97828 85474 97856 91151
rect 97816 85468 97868 85474
rect 97816 85410 97868 85416
rect 98748 85202 98776 91151
rect 99024 90914 99052 92375
rect 101862 91760 101918 91769
rect 101862 91695 101918 91704
rect 99102 91216 99158 91225
rect 99102 91151 99158 91160
rect 100206 91216 100262 91225
rect 100206 91151 100262 91160
rect 99012 90908 99064 90914
rect 99012 90850 99064 90856
rect 98736 85196 98788 85202
rect 98736 85138 98788 85144
rect 95148 84108 95200 84114
rect 95148 84050 95200 84056
rect 67640 82816 67692 82822
rect 67640 82758 67692 82764
rect 99116 82754 99144 91151
rect 100220 86766 100248 91151
rect 101876 89690 101904 91695
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 101864 89684 101916 89690
rect 101864 89626 101916 89632
rect 100208 86760 100260 86766
rect 100208 86702 100260 86708
rect 101968 83978 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 102874 91216 102930 91225
rect 102874 91151 102930 91160
rect 102060 84182 102088 91151
rect 102888 88262 102916 91151
rect 104452 91050 104480 92375
rect 105740 92206 105768 92375
rect 105728 92200 105780 92206
rect 105728 92142 105780 92148
rect 104440 91044 104492 91050
rect 104440 90986 104492 90992
rect 106752 90846 106780 92375
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 107934 91216 107990 91225
rect 107934 91151 107990 91160
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 106740 90840 106792 90846
rect 106740 90782 106792 90788
rect 102876 88256 102928 88262
rect 102876 88198 102928 88204
rect 102048 84176 102100 84182
rect 102048 84118 102100 84124
rect 101956 83972 102008 83978
rect 101956 83914 102008 83920
rect 99104 82748 99156 82754
rect 99104 82690 99156 82696
rect 106188 82136 106240 82142
rect 106188 82078 106240 82084
rect 79324 80708 79376 80714
rect 79324 80650 79376 80656
rect 71044 79348 71096 79354
rect 71044 79290 71096 79296
rect 67548 78668 67600 78674
rect 67548 78610 67600 78616
rect 70308 72480 70360 72486
rect 70308 72422 70360 72428
rect 57244 71732 57296 71738
rect 57244 71674 57296 71680
rect 65984 71732 66036 71738
rect 65984 71674 66036 71680
rect 68928 69692 68980 69698
rect 68928 69634 68980 69640
rect 57886 61432 57942 61441
rect 57886 61367 57942 61376
rect 55128 51808 55180 51814
rect 55128 51750 55180 51756
rect 54484 49020 54536 49026
rect 54484 48962 54536 48968
rect 55140 6914 55168 51750
rect 56508 21412 56560 21418
rect 56508 21354 56560 21360
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 21354
rect 57900 3534 57928 61367
rect 65524 49020 65576 49026
rect 65524 48962 65576 48968
rect 58624 47660 58676 47666
rect 58624 47602 58676 47608
rect 58636 3670 58664 47602
rect 62028 32428 62080 32434
rect 62028 32370 62080 32376
rect 59268 14476 59320 14482
rect 59268 14418 59320 14424
rect 58624 3664 58676 3670
rect 58624 3606 58676 3612
rect 59280 3534 59308 14418
rect 60648 13116 60700 13122
rect 60648 13058 60700 13064
rect 60660 3534 60688 13058
rect 60832 6180 60884 6186
rect 60832 6122 60884 6128
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 6122
rect 62040 480 62068 32370
rect 65536 6914 65564 48962
rect 67546 43480 67602 43489
rect 67546 43415 67602 43424
rect 66168 15904 66220 15910
rect 66168 15846 66220 15852
rect 65444 6886 65564 6914
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 63224 2100 63276 2106
rect 63224 2042 63276 2048
rect 63236 480 63264 2042
rect 64340 480 64368 3470
rect 65444 2174 65472 6886
rect 66180 3534 66208 15846
rect 67560 3534 67588 43415
rect 68940 3534 68968 69634
rect 70216 46232 70268 46238
rect 70216 46174 70268 46180
rect 70228 3534 70256 46174
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 65432 2168 65484 2174
rect 65432 2110 65484 2116
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70320 480 70348 72422
rect 71056 3738 71084 79290
rect 73068 76628 73120 76634
rect 73068 76570 73120 76576
rect 71688 44872 71740 44878
rect 71688 44814 71740 44820
rect 71700 6914 71728 44814
rect 71516 6886 71728 6914
rect 71044 3732 71096 3738
rect 71044 3674 71096 3680
rect 71516 480 71544 6886
rect 73080 3534 73108 76570
rect 75828 73976 75880 73982
rect 75828 73918 75880 73924
rect 73804 4888 73856 4894
rect 73804 4830 73856 4836
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 72620 480 72648 3470
rect 73816 480 73844 4830
rect 75840 3534 75868 73918
rect 77208 66904 77260 66910
rect 77208 66846 77260 66852
rect 77220 3534 77248 66846
rect 78588 33788 78640 33794
rect 78588 33730 78640 33736
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 77392 3528 77444 3534
rect 77392 3470 77444 3476
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 3470
rect 78600 480 78628 33730
rect 79336 3602 79364 80650
rect 102048 78056 102100 78062
rect 102048 77998 102100 78004
rect 91008 75268 91060 75274
rect 91008 75210 91060 75216
rect 89628 72548 89680 72554
rect 89628 72490 89680 72496
rect 86868 71052 86920 71058
rect 86868 70994 86920 71000
rect 84108 65544 84160 65550
rect 84108 65486 84160 65492
rect 82728 35284 82780 35290
rect 82728 35226 82780 35232
rect 81348 28348 81400 28354
rect 81348 28290 81400 28296
rect 79692 10328 79744 10334
rect 79692 10270 79744 10276
rect 79324 3596 79376 3602
rect 79324 3538 79376 3544
rect 79704 480 79732 10270
rect 81360 3534 81388 28290
rect 82740 3534 82768 35226
rect 84120 3534 84148 65486
rect 86776 58676 86828 58682
rect 86776 58618 86828 58624
rect 86788 16574 86816 58618
rect 86696 16546 86816 16574
rect 85488 11824 85540 11830
rect 85488 11766 85540 11772
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 83292 480 83320 3470
rect 85500 3466 85528 11766
rect 85672 3664 85724 3670
rect 85672 3606 85724 3612
rect 84476 3460 84528 3466
rect 84476 3402 84528 3408
rect 85488 3460 85540 3466
rect 85488 3402 85540 3408
rect 84488 480 84516 3402
rect 85684 480 85712 3606
rect 86696 3482 86724 16546
rect 86880 6914 86908 70994
rect 88248 68332 88300 68338
rect 88248 68274 88300 68280
rect 88260 6914 88288 68274
rect 86788 6886 86908 6914
rect 87984 6886 88288 6914
rect 86788 3670 86816 6886
rect 86776 3664 86828 3670
rect 86776 3606 86828 3612
rect 86696 3454 86908 3482
rect 86880 480 86908 3454
rect 87984 480 88012 6886
rect 89640 3534 89668 72490
rect 91020 3534 91048 75210
rect 95148 74044 95200 74050
rect 95148 73986 95200 73992
rect 93768 61396 93820 61402
rect 93768 61338 93820 61344
rect 92388 44940 92440 44946
rect 92388 44882 92440 44888
rect 92400 3534 92428 44882
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 89180 480 89208 3470
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 93780 2922 93808 61338
rect 95160 3534 95188 73986
rect 97908 62892 97960 62898
rect 97908 62834 97960 62840
rect 96528 32496 96580 32502
rect 96528 32438 96580 32444
rect 96540 6914 96568 32438
rect 96264 6886 96568 6914
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 93768 2916 93820 2922
rect 93768 2858 93820 2864
rect 92768 480 92796 2858
rect 93964 480 93992 3470
rect 95148 3392 95200 3398
rect 95148 3334 95200 3340
rect 95160 480 95188 3334
rect 96264 480 96292 6886
rect 97920 3534 97948 62834
rect 99288 40724 99340 40730
rect 99288 40666 99340 40672
rect 99300 3534 99328 40666
rect 100668 36576 100720 36582
rect 100668 36518 100720 36524
rect 100680 3534 100708 36518
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 102060 3194 102088 77998
rect 104164 50380 104216 50386
rect 104164 50322 104216 50328
rect 103428 38004 103480 38010
rect 103428 37946 103480 37952
rect 103440 6914 103468 37946
rect 103348 6886 103468 6914
rect 102232 6248 102284 6254
rect 102232 6190 102284 6196
rect 101036 3188 101088 3194
rect 101036 3130 101088 3136
rect 102048 3188 102100 3194
rect 102048 3130 102100 3136
rect 101048 480 101076 3130
rect 102244 480 102272 6190
rect 103348 480 103376 6886
rect 104176 3602 104204 50322
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 104164 3596 104216 3602
rect 104164 3538 104216 3544
rect 104544 480 104572 8910
rect 106200 3602 106228 82078
rect 107580 77246 107608 91151
rect 107948 88330 107976 91151
rect 107936 88324 107988 88330
rect 107936 88266 107988 88272
rect 108960 81258 108988 91151
rect 110156 89418 110184 93191
rect 113270 92440 113326 92449
rect 113270 92375 113272 92384
rect 113324 92375 113326 92384
rect 113272 92346 113324 92352
rect 111338 91216 111394 91225
rect 111338 91151 111394 91160
rect 112074 91216 112130 91225
rect 112074 91151 112130 91160
rect 112718 91216 112774 91225
rect 112718 91151 112774 91160
rect 110144 89412 110196 89418
rect 110144 89354 110196 89360
rect 111352 86834 111380 91151
rect 111340 86828 111392 86834
rect 111340 86770 111392 86776
rect 112088 86698 112116 91151
rect 112732 86970 112760 91151
rect 113836 88194 113864 93191
rect 118252 93158 118280 93463
rect 125428 93362 125456 93463
rect 151596 93463 151598 93472
rect 152094 93528 152150 93537
rect 152094 93463 152150 93472
rect 151544 93434 151596 93440
rect 152108 93430 152136 93463
rect 152096 93424 152148 93430
rect 152096 93366 152148 93372
rect 125416 93356 125468 93362
rect 125416 93298 125468 93304
rect 118240 93152 118292 93158
rect 118240 93094 118292 93100
rect 115754 92440 115810 92449
rect 115754 92375 115810 92384
rect 121182 92440 121238 92449
rect 121182 92375 121238 92384
rect 123022 92440 123078 92449
rect 123022 92375 123078 92384
rect 125782 92440 125838 92449
rect 125782 92375 125838 92384
rect 136178 92440 136234 92449
rect 136178 92375 136234 92384
rect 115768 92274 115796 92375
rect 115756 92268 115808 92274
rect 115756 92210 115808 92216
rect 117134 91760 117190 91769
rect 117134 91695 117190 91704
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 115018 91216 115074 91225
rect 115018 91151 115074 91160
rect 116584 91180 116636 91186
rect 113824 88188 113876 88194
rect 113824 88130 113876 88136
rect 112720 86964 112772 86970
rect 112720 86906 112772 86912
rect 112076 86692 112128 86698
rect 112076 86634 112128 86640
rect 114480 84046 114508 91151
rect 115032 85270 115060 91151
rect 116584 91122 116636 91128
rect 115204 91112 115256 91118
rect 115204 91054 115256 91060
rect 115020 85264 115072 85270
rect 115020 85206 115072 85212
rect 114468 84040 114520 84046
rect 114468 83982 114520 83988
rect 108948 81252 109000 81258
rect 108948 81194 109000 81200
rect 113088 80776 113140 80782
rect 113088 80718 113140 80724
rect 108948 79416 109000 79422
rect 108948 79358 109000 79364
rect 107568 77240 107620 77246
rect 107568 77182 107620 77188
rect 107568 69828 107620 69834
rect 107568 69770 107620 69776
rect 107580 3602 107608 69770
rect 108960 3602 108988 79358
rect 111708 69760 111760 69766
rect 111708 69702 111760 69708
rect 111616 55956 111668 55962
rect 111616 55898 111668 55904
rect 110328 42152 110380 42158
rect 110328 42094 110380 42100
rect 110340 3602 110368 42094
rect 105728 3596 105780 3602
rect 105728 3538 105780 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 106924 3596 106976 3602
rect 106924 3538 106976 3544
rect 107568 3596 107620 3602
rect 107568 3538 107620 3544
rect 108120 3596 108172 3602
rect 108120 3538 108172 3544
rect 108948 3596 109000 3602
rect 108948 3538 109000 3544
rect 109316 3596 109368 3602
rect 109316 3538 109368 3544
rect 110328 3596 110380 3602
rect 110328 3538 110380 3544
rect 105740 480 105768 3538
rect 106936 480 106964 3538
rect 108132 480 108160 3538
rect 109328 480 109356 3538
rect 110512 3188 110564 3194
rect 110512 3130 110564 3136
rect 110524 480 110552 3130
rect 111628 480 111656 55898
rect 111720 3194 111748 69702
rect 113100 6914 113128 80718
rect 115216 75886 115244 91054
rect 115204 75880 115256 75886
rect 115204 75822 115256 75828
rect 116596 74526 116624 91122
rect 117148 89554 117176 91695
rect 119710 91216 119766 91225
rect 119710 91151 119766 91160
rect 117136 89548 117188 89554
rect 117136 89490 117188 89496
rect 119724 85406 119752 91151
rect 121196 90778 121224 92375
rect 123036 92342 123064 92375
rect 123024 92336 123076 92342
rect 123024 92278 123076 92284
rect 125796 92138 125824 92375
rect 125784 92132 125836 92138
rect 125784 92074 125836 92080
rect 126610 91624 126666 91633
rect 126610 91559 126666 91568
rect 121274 91216 121330 91225
rect 121274 91151 121330 91160
rect 121918 91216 121974 91225
rect 121918 91151 121974 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 123298 91216 123354 91225
rect 123298 91151 123354 91160
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 121184 90772 121236 90778
rect 121184 90714 121236 90720
rect 119712 85400 119764 85406
rect 119712 85342 119764 85348
rect 119986 84824 120042 84833
rect 119986 84759 120042 84768
rect 116584 74520 116636 74526
rect 116584 74462 116636 74468
rect 115848 72616 115900 72622
rect 115848 72558 115900 72564
rect 114468 29708 114520 29714
rect 114468 29650 114520 29656
rect 112824 6886 113128 6914
rect 111708 3188 111760 3194
rect 111708 3130 111760 3136
rect 112824 480 112852 6886
rect 114480 3602 114508 29650
rect 115860 3602 115888 72558
rect 117228 68400 117280 68406
rect 117228 68342 117280 68348
rect 117240 3602 117268 68342
rect 119896 58744 119948 58750
rect 119896 58686 119948 58692
rect 118608 26988 118660 26994
rect 118608 26930 118660 26936
rect 118620 3602 118648 26930
rect 119908 16574 119936 58686
rect 119816 16546 119936 16574
rect 119816 3602 119844 16546
rect 120000 6914 120028 84759
rect 121288 82618 121316 91151
rect 121932 86630 121960 91151
rect 121920 86624 121972 86630
rect 121920 86566 121972 86572
rect 122760 82686 122788 91151
rect 123312 88233 123340 91151
rect 123298 88224 123354 88233
rect 123298 88159 123354 88168
rect 124140 87990 124168 91151
rect 126624 89350 126652 91559
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 131026 91216 131082 91225
rect 131026 91151 131082 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 133786 91216 133842 91225
rect 133786 91151 133842 91160
rect 135166 91216 135222 91225
rect 135166 91151 135222 91160
rect 126612 89344 126664 89350
rect 126612 89286 126664 89292
rect 124128 87984 124180 87990
rect 124128 87926 124180 87932
rect 122748 82680 122800 82686
rect 122748 82622 122800 82628
rect 121276 82612 121328 82618
rect 121276 82554 121328 82560
rect 124128 79484 124180 79490
rect 124128 79426 124180 79432
rect 122748 71120 122800 71126
rect 122748 71062 122800 71068
rect 119908 6886 120028 6914
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 117596 3596 117648 3602
rect 117596 3538 117648 3544
rect 118608 3596 118660 3602
rect 118608 3538 118660 3544
rect 118792 3596 118844 3602
rect 118792 3538 118844 3544
rect 119804 3596 119856 3602
rect 119804 3538 119856 3544
rect 114020 480 114048 3538
rect 115216 480 115244 3538
rect 116412 480 116440 3538
rect 117608 480 117636 3538
rect 118804 480 118832 3538
rect 119908 480 119936 6886
rect 122760 3602 122788 71062
rect 124140 3602 124168 79426
rect 126900 78538 126928 91151
rect 128280 79966 128308 91151
rect 129660 81326 129688 91151
rect 129648 81320 129700 81326
rect 129648 81262 129700 81268
rect 128268 79960 128320 79966
rect 128268 79902 128320 79908
rect 126888 78532 126940 78538
rect 126888 78474 126940 78480
rect 131040 77178 131068 91151
rect 132420 83910 132448 91151
rect 132408 83904 132460 83910
rect 132408 83846 132460 83852
rect 131028 77172 131080 77178
rect 131028 77114 131080 77120
rect 125508 76696 125560 76702
rect 125508 76638 125560 76644
rect 125520 3602 125548 76638
rect 133800 75818 133828 91151
rect 135180 78606 135208 91151
rect 136192 90710 136220 92375
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 136180 90704 136232 90710
rect 136180 90646 136232 90652
rect 151740 82550 151768 91151
rect 164896 89486 164924 97990
rect 166276 94178 166304 153206
rect 170404 151836 170456 151842
rect 170404 151778 170456 151784
rect 166356 147688 166408 147694
rect 166356 147630 166408 147636
rect 166264 94172 166316 94178
rect 166264 94114 166316 94120
rect 166368 90710 166396 147630
rect 169024 136672 169076 136678
rect 169024 136614 169076 136620
rect 167736 131164 167788 131170
rect 167736 131106 167788 131112
rect 167644 125656 167696 125662
rect 167644 125598 167696 125604
rect 166448 109064 166500 109070
rect 166448 109006 166500 109012
rect 166356 90704 166408 90710
rect 166356 90646 166408 90652
rect 164884 89480 164936 89486
rect 164884 89422 164936 89428
rect 166460 88058 166488 109006
rect 166540 99408 166592 99414
rect 166540 99350 166592 99356
rect 166448 88052 166500 88058
rect 166448 87994 166500 88000
rect 166552 85338 166580 99350
rect 167656 89350 167684 125598
rect 167748 93945 167776 131106
rect 167828 111784 167880 111790
rect 167826 111752 167828 111761
rect 167880 111752 167882 111761
rect 167826 111687 167882 111696
rect 167828 110424 167880 110430
rect 167828 110366 167880 110372
rect 167840 110129 167868 110366
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 167828 108996 167880 109002
rect 167828 108938 167880 108944
rect 167840 108769 167868 108938
rect 167826 108760 167882 108769
rect 167826 108695 167882 108704
rect 167828 107704 167880 107710
rect 167828 107646 167880 107652
rect 167734 93936 167790 93945
rect 167734 93871 167790 93880
rect 167644 89344 167696 89350
rect 167644 89286 167696 89292
rect 167840 88126 167868 107646
rect 169036 93673 169064 136614
rect 169116 111852 169168 111858
rect 169116 111794 169168 111800
rect 169022 93664 169078 93673
rect 169022 93599 169078 93608
rect 169128 93294 169156 111794
rect 169208 106956 169260 106962
rect 169208 106898 169260 106904
rect 169116 93288 169168 93294
rect 169116 93230 169168 93236
rect 169220 92206 169248 106898
rect 169300 99476 169352 99482
rect 169300 99418 169352 99424
rect 169208 92200 169260 92206
rect 169208 92142 169260 92148
rect 167828 88120 167880 88126
rect 167828 88062 167880 88068
rect 169312 86902 169340 99418
rect 170416 93498 170444 151778
rect 177396 140820 177448 140826
rect 177396 140762 177448 140768
rect 177304 138712 177356 138718
rect 177304 138654 177356 138660
rect 173348 133952 173400 133958
rect 173348 133894 173400 133900
rect 173256 132524 173308 132530
rect 173256 132466 173308 132472
rect 170496 128376 170548 128382
rect 170496 128318 170548 128324
rect 170404 93492 170456 93498
rect 170404 93434 170456 93440
rect 169300 86896 169352 86902
rect 169300 86838 169352 86844
rect 166540 85332 166592 85338
rect 166540 85274 166592 85280
rect 170508 83978 170536 128318
rect 171784 122868 171836 122874
rect 171784 122810 171836 122816
rect 170588 103556 170640 103562
rect 170588 103498 170640 103504
rect 170496 83972 170548 83978
rect 170496 83914 170548 83920
rect 151728 82544 151780 82550
rect 151728 82486 151780 82492
rect 170600 80034 170628 103498
rect 171796 90778 171824 122810
rect 171876 117360 171928 117366
rect 171876 117302 171928 117308
rect 171784 90772 171836 90778
rect 171784 90714 171836 90720
rect 171888 89418 171916 117302
rect 173164 96688 173216 96694
rect 173164 96630 173216 96636
rect 171876 89412 171928 89418
rect 171876 89354 171928 89360
rect 170588 80028 170640 80034
rect 170588 79970 170640 79976
rect 135168 78600 135220 78606
rect 135168 78542 135220 78548
rect 133788 75812 133840 75818
rect 133788 75754 133840 75760
rect 173176 4826 173204 96630
rect 173268 77246 173296 132466
rect 173360 94110 173388 133894
rect 175924 132592 175976 132598
rect 175924 132534 175976 132540
rect 174636 129804 174688 129810
rect 174636 129746 174688 129752
rect 174544 127016 174596 127022
rect 174544 126958 174596 126964
rect 173440 122936 173492 122942
rect 173440 122878 173492 122884
rect 173348 94104 173400 94110
rect 173348 94046 173400 94052
rect 173452 86630 173480 122878
rect 173440 86624 173492 86630
rect 173440 86566 173492 86572
rect 174556 85202 174584 126958
rect 174648 92177 174676 129746
rect 174634 92168 174690 92177
rect 174634 92103 174690 92112
rect 174544 85196 174596 85202
rect 174544 85138 174596 85144
rect 175936 81258 175964 132534
rect 176016 100768 176068 100774
rect 176016 100710 176068 100716
rect 176028 89593 176056 100710
rect 177316 92138 177344 138654
rect 177304 92132 177356 92138
rect 177304 92074 177356 92080
rect 177408 90953 177436 140762
rect 177580 114572 177632 114578
rect 177580 114514 177632 114520
rect 177488 110492 177540 110498
rect 177488 110434 177540 110440
rect 177394 90944 177450 90953
rect 177394 90879 177450 90888
rect 177304 90364 177356 90370
rect 177304 90306 177356 90312
rect 176014 89584 176070 89593
rect 176014 89519 176070 89528
rect 175924 81252 175976 81258
rect 175924 81194 175976 81200
rect 173256 77240 173308 77246
rect 173256 77182 173308 77188
rect 173164 4820 173216 4826
rect 173164 4762 173216 4768
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 124680 3596 124732 3602
rect 124680 3538 124732 3544
rect 125508 3596 125560 3602
rect 125508 3538 125560 3544
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 121090 3360 121146 3369
rect 121090 3295 121146 3304
rect 121104 480 121132 3295
rect 122300 480 122328 3538
rect 123496 480 123524 3538
rect 124692 480 124720 3538
rect 125888 480 125916 3538
rect 177316 3466 177344 90306
rect 177500 86766 177528 110434
rect 177592 93226 177620 114514
rect 177580 93220 177632 93226
rect 177580 93162 177632 93168
rect 177488 86760 177540 86766
rect 177488 86702 177540 86708
rect 178696 3602 178724 229842
rect 180628 193866 180656 252554
rect 180720 248402 180748 697546
rect 196624 670744 196676 670750
rect 196624 670686 196676 670692
rect 191748 623076 191800 623082
rect 191748 623018 191800 623024
rect 188988 456816 189040 456822
rect 188988 456758 189040 456764
rect 182088 286000 182140 286006
rect 182088 285942 182140 285948
rect 180708 248396 180760 248402
rect 180708 248338 180760 248344
rect 180616 193860 180668 193866
rect 180616 193802 180668 193808
rect 182100 189922 182128 285942
rect 183468 281648 183520 281654
rect 183468 281590 183520 281596
rect 182088 189916 182140 189922
rect 182088 189858 182140 189864
rect 183480 181694 183508 281590
rect 188896 278792 188948 278798
rect 188896 278734 188948 278740
rect 187608 274712 187660 274718
rect 187608 274654 187660 274660
rect 184848 273284 184900 273290
rect 184848 273226 184900 273232
rect 184756 263628 184808 263634
rect 184756 263570 184808 263576
rect 183468 181688 183520 181694
rect 183468 181630 183520 181636
rect 184388 181008 184440 181014
rect 184388 180950 184440 180956
rect 182824 179580 182876 179586
rect 182824 179522 182876 179528
rect 181444 179512 181496 179518
rect 181444 179454 181496 179460
rect 180064 178152 180116 178158
rect 180064 178094 180116 178100
rect 178774 177168 178830 177177
rect 178774 177103 178830 177112
rect 178788 163538 178816 177103
rect 178776 163532 178828 163538
rect 178776 163474 178828 163480
rect 180076 162858 180104 178094
rect 180064 162852 180116 162858
rect 180064 162794 180116 162800
rect 181456 161362 181484 179454
rect 182836 162790 182864 179522
rect 184296 175976 184348 175982
rect 184296 175918 184348 175924
rect 184204 171148 184256 171154
rect 184204 171090 184256 171096
rect 182824 162784 182876 162790
rect 182824 162726 182876 162732
rect 181444 161356 181496 161362
rect 181444 161298 181496 161304
rect 180064 153332 180116 153338
rect 180064 153274 180116 153280
rect 178776 124228 178828 124234
rect 178776 124170 178828 124176
rect 178788 87990 178816 124170
rect 178868 110560 178920 110566
rect 178868 110502 178920 110508
rect 178880 90914 178908 110502
rect 178868 90908 178920 90914
rect 178868 90850 178920 90856
rect 178776 87984 178828 87990
rect 178776 87926 178828 87932
rect 180076 82550 180104 153274
rect 184216 150414 184244 171090
rect 184308 165510 184336 175918
rect 184400 172446 184428 180950
rect 184768 178702 184796 263570
rect 184860 182889 184888 273226
rect 187516 270632 187568 270638
rect 187516 270574 187568 270580
rect 186228 270564 186280 270570
rect 186228 270506 186280 270512
rect 186136 253224 186188 253230
rect 186136 253166 186188 253172
rect 184846 182880 184902 182889
rect 184846 182815 184902 182824
rect 186148 178770 186176 253166
rect 186240 180033 186268 270506
rect 187424 259480 187476 259486
rect 187424 259422 187476 259428
rect 187436 181626 187464 259422
rect 187528 189689 187556 270574
rect 187620 192574 187648 274654
rect 188804 256760 188856 256766
rect 188804 256702 188856 256708
rect 188712 248464 188764 248470
rect 188712 248406 188764 248412
rect 187608 192568 187660 192574
rect 187608 192510 187660 192516
rect 187514 189680 187570 189689
rect 187514 189615 187570 189624
rect 188724 187066 188752 248406
rect 188816 211818 188844 256702
rect 188804 211812 188856 211818
rect 188804 211754 188856 211760
rect 188712 187060 188764 187066
rect 188712 187002 188764 187008
rect 187424 181620 187476 181626
rect 187424 181562 187476 181568
rect 186226 180024 186282 180033
rect 186226 179959 186282 179968
rect 186136 178764 186188 178770
rect 186136 178706 186188 178712
rect 184756 178696 184808 178702
rect 184756 178638 184808 178644
rect 186964 178220 187016 178226
rect 186964 178162 187016 178168
rect 184388 172440 184440 172446
rect 184388 172382 184440 172388
rect 186976 171018 187004 178162
rect 188908 175982 188936 278734
rect 189000 242894 189028 456758
rect 191656 276072 191708 276078
rect 191656 276014 191708 276020
rect 190368 273352 190420 273358
rect 190368 273294 190420 273300
rect 190276 248532 190328 248538
rect 190276 248474 190328 248480
rect 188988 242888 189040 242894
rect 188988 242830 189040 242836
rect 190288 181529 190316 248474
rect 190380 186969 190408 273294
rect 191564 258596 191616 258602
rect 191564 258538 191616 258544
rect 191472 254040 191524 254046
rect 191472 253982 191524 253988
rect 191484 209098 191512 253982
rect 191472 209092 191524 209098
rect 191472 209034 191524 209040
rect 190366 186960 190422 186969
rect 190366 186895 190422 186904
rect 190274 181520 190330 181529
rect 190274 181455 190330 181464
rect 191104 177132 191156 177138
rect 191104 177074 191156 177080
rect 188896 175976 188948 175982
rect 188896 175918 188948 175924
rect 186964 171012 187016 171018
rect 186964 170954 187016 170960
rect 184296 165504 184348 165510
rect 184296 165446 184348 165452
rect 191116 160002 191144 177074
rect 191576 176594 191604 258538
rect 191668 184210 191696 276014
rect 191760 244186 191788 623018
rect 195796 293276 195848 293282
rect 195796 293218 195848 293224
rect 194508 285864 194560 285870
rect 194508 285806 194560 285812
rect 194416 277772 194468 277778
rect 194416 277714 194468 277720
rect 193128 269204 193180 269210
rect 193128 269146 193180 269152
rect 193036 262268 193088 262274
rect 193036 262210 193088 262216
rect 192944 255332 192996 255338
rect 192944 255274 192996 255280
rect 191748 244180 191800 244186
rect 191748 244122 191800 244128
rect 191748 241528 191800 241534
rect 191748 241470 191800 241476
rect 191656 184204 191708 184210
rect 191656 184146 191708 184152
rect 191760 177313 191788 241470
rect 192956 189786 192984 255274
rect 192944 189780 192996 189786
rect 192944 189722 192996 189728
rect 193048 186998 193076 262210
rect 193140 187105 193168 269146
rect 194324 253020 194376 253026
rect 194324 252962 194376 252968
rect 194336 229770 194364 252962
rect 194324 229764 194376 229770
rect 194324 229706 194376 229712
rect 194428 191049 194456 277714
rect 194414 191040 194470 191049
rect 194414 190975 194470 190984
rect 193126 187096 193182 187105
rect 193126 187031 193182 187040
rect 193036 186992 193088 186998
rect 193036 186934 193088 186940
rect 191746 177304 191802 177313
rect 191746 177239 191802 177248
rect 191564 176588 191616 176594
rect 191564 176530 191616 176536
rect 194520 175098 194548 285806
rect 195612 266416 195664 266422
rect 195612 266358 195664 266364
rect 195624 232626 195652 266358
rect 195704 256828 195756 256834
rect 195704 256770 195756 256776
rect 195612 232620 195664 232626
rect 195612 232562 195664 232568
rect 195716 188426 195744 256770
rect 195808 256698 195836 293218
rect 196636 287094 196664 670686
rect 202144 660340 202196 660346
rect 202144 660282 202196 660288
rect 198648 380180 198700 380186
rect 198648 380122 198700 380128
rect 198554 295352 198610 295361
rect 198554 295287 198610 295296
rect 196624 287088 196676 287094
rect 196624 287030 196676 287036
rect 195888 286068 195940 286074
rect 195888 286010 195940 286016
rect 195796 256692 195848 256698
rect 195796 256634 195848 256640
rect 195796 247104 195848 247110
rect 195796 247046 195848 247052
rect 195704 188420 195756 188426
rect 195704 188362 195756 188368
rect 195808 178838 195836 247046
rect 195900 184249 195928 286010
rect 198568 282985 198596 295287
rect 198554 282976 198610 282985
rect 198554 282911 198610 282920
rect 197450 282432 197506 282441
rect 197450 282367 197506 282376
rect 197464 281654 197492 282367
rect 197452 281648 197504 281654
rect 197358 281616 197414 281625
rect 197452 281590 197504 281596
rect 197358 281551 197360 281560
rect 197412 281551 197414 281560
rect 197360 281522 197412 281528
rect 198660 280809 198688 380122
rect 200396 289196 200448 289202
rect 200396 289138 200448 289144
rect 200028 285796 200080 285802
rect 200028 285738 200080 285744
rect 199936 285728 199988 285734
rect 199936 285670 199988 285676
rect 198646 280800 198702 280809
rect 198646 280735 198702 280744
rect 197174 280256 197230 280265
rect 197174 280191 197230 280200
rect 196990 260944 197046 260953
rect 196990 260879 197046 260888
rect 197004 228410 197032 260879
rect 197082 250880 197138 250889
rect 197082 250815 197138 250824
rect 196992 228404 197044 228410
rect 196992 228346 197044 228352
rect 197096 184414 197124 250815
rect 197188 189854 197216 280191
rect 197358 279440 197414 279449
rect 197358 279375 197414 279384
rect 197372 278798 197400 279375
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 198002 278624 198058 278633
rect 198002 278559 198058 278568
rect 197358 278080 197414 278089
rect 197358 278015 197414 278024
rect 197372 277778 197400 278015
rect 197360 277772 197412 277778
rect 197360 277714 197412 277720
rect 197450 277264 197506 277273
rect 197450 277199 197506 277208
rect 197266 276720 197322 276729
rect 197266 276655 197322 276664
rect 197176 189848 197228 189854
rect 197176 189790 197228 189796
rect 197084 184408 197136 184414
rect 197084 184350 197136 184356
rect 195886 184240 195942 184249
rect 195886 184175 195942 184184
rect 195796 178832 195848 178838
rect 195796 178774 195848 178780
rect 197280 178673 197308 276655
rect 197464 276078 197492 277199
rect 197452 276072 197504 276078
rect 197452 276014 197504 276020
rect 197360 276004 197412 276010
rect 197360 275946 197412 275952
rect 197372 275913 197400 275946
rect 197358 275904 197414 275913
rect 197358 275839 197414 275848
rect 197358 275088 197414 275097
rect 197358 275023 197414 275032
rect 197372 274718 197400 275023
rect 197360 274712 197412 274718
rect 197360 274654 197412 274660
rect 197450 274544 197506 274553
rect 197450 274479 197506 274488
rect 197358 273728 197414 273737
rect 197358 273663 197414 273672
rect 197372 273290 197400 273663
rect 197464 273358 197492 274479
rect 197452 273352 197504 273358
rect 197452 273294 197504 273300
rect 197360 273284 197412 273290
rect 197360 273226 197412 273232
rect 197452 273216 197504 273222
rect 197452 273158 197504 273164
rect 197464 272377 197492 273158
rect 197450 272368 197506 272377
rect 197450 272303 197506 272312
rect 197450 271552 197506 271561
rect 197450 271487 197506 271496
rect 197358 271008 197414 271017
rect 197358 270943 197414 270952
rect 197372 270638 197400 270943
rect 197360 270632 197412 270638
rect 197360 270574 197412 270580
rect 197464 270570 197492 271487
rect 197452 270564 197504 270570
rect 197452 270506 197504 270512
rect 197450 270192 197506 270201
rect 197450 270127 197506 270136
rect 197358 269376 197414 269385
rect 197358 269311 197414 269320
rect 197372 269142 197400 269311
rect 197464 269210 197492 270127
rect 197452 269204 197504 269210
rect 197452 269146 197504 269152
rect 197360 269136 197412 269142
rect 197360 269078 197412 269084
rect 197452 269068 197504 269074
rect 197452 269010 197504 269016
rect 197360 269000 197412 269006
rect 197360 268942 197412 268948
rect 197372 268025 197400 268942
rect 197464 268841 197492 269010
rect 197450 268832 197506 268841
rect 197450 268767 197506 268776
rect 197358 268016 197414 268025
rect 197358 267951 197414 267960
rect 197360 267708 197412 267714
rect 197360 267650 197412 267656
rect 197372 266665 197400 267650
rect 197910 267200 197966 267209
rect 197910 267135 197966 267144
rect 197358 266656 197414 266665
rect 197358 266591 197414 266600
rect 197924 266422 197952 267135
rect 197912 266416 197964 266422
rect 197912 266358 197964 266364
rect 197450 265840 197506 265849
rect 197450 265775 197506 265784
rect 197464 264994 197492 265775
rect 197452 264988 197504 264994
rect 197452 264930 197504 264936
rect 197360 264920 197412 264926
rect 197360 264862 197412 264868
rect 197372 264489 197400 264862
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197358 263664 197414 263673
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197450 262304 197506 262313
rect 197450 262239 197452 262248
rect 197504 262239 197506 262248
rect 197452 262210 197504 262216
rect 197360 262200 197412 262206
rect 197360 262142 197412 262148
rect 197372 261497 197400 262142
rect 197358 261488 197414 261497
rect 197358 261423 197414 261432
rect 197358 260128 197414 260137
rect 197358 260063 197414 260072
rect 197372 259486 197400 260063
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197450 259312 197506 259321
rect 197450 259247 197506 259256
rect 197358 258768 197414 258777
rect 197358 258703 197414 258712
rect 197372 258126 197400 258703
rect 197464 258602 197492 259247
rect 197452 258596 197504 258602
rect 197452 258538 197504 258544
rect 197360 258120 197412 258126
rect 197360 258062 197412 258068
rect 197358 257952 197414 257961
rect 197358 257887 197414 257896
rect 197372 256766 197400 257887
rect 197542 257408 197598 257417
rect 197542 257343 197598 257352
rect 197556 256834 197584 257343
rect 197544 256828 197596 256834
rect 197544 256770 197596 256776
rect 197360 256760 197412 256766
rect 197360 256702 197412 256708
rect 197912 256692 197964 256698
rect 197912 256634 197964 256640
rect 197358 256592 197414 256601
rect 197358 256527 197414 256536
rect 197372 255338 197400 256527
rect 197924 255785 197952 256634
rect 197910 255776 197966 255785
rect 197910 255711 197966 255720
rect 197360 255332 197412 255338
rect 197360 255274 197412 255280
rect 197450 255232 197506 255241
rect 197450 255167 197506 255176
rect 197358 254416 197414 254425
rect 197358 254351 197414 254360
rect 197372 253978 197400 254351
rect 197464 254046 197492 255167
rect 197452 254040 197504 254046
rect 197452 253982 197504 253988
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197358 253600 197414 253609
rect 197358 253535 197414 253544
rect 197372 252618 197400 253535
rect 198016 253230 198044 278559
rect 198554 272912 198610 272921
rect 198554 272847 198610 272856
rect 198094 265296 198150 265305
rect 198094 265231 198150 265240
rect 198004 253224 198056 253230
rect 198004 253166 198056 253172
rect 198108 253026 198136 265231
rect 198568 259457 198596 272847
rect 198646 263120 198702 263129
rect 198646 263055 198702 263064
rect 198554 259448 198610 259457
rect 198554 259383 198610 259392
rect 198554 253056 198610 253065
rect 198096 253020 198148 253026
rect 198554 252991 198610 253000
rect 198096 252962 198148 252968
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 198370 251696 198426 251705
rect 198370 251631 198426 251640
rect 197360 251184 197412 251190
rect 197360 251126 197412 251132
rect 197372 250073 197400 251126
rect 197358 250064 197414 250073
rect 197358 249999 197414 250008
rect 197450 249520 197506 249529
rect 197450 249455 197506 249464
rect 197358 248704 197414 248713
rect 197358 248639 197414 248648
rect 197372 248538 197400 248639
rect 197360 248532 197412 248538
rect 197360 248474 197412 248480
rect 197464 248470 197492 249455
rect 197452 248464 197504 248470
rect 197452 248406 197504 248412
rect 197360 248396 197412 248402
rect 197360 248338 197412 248344
rect 197372 247353 197400 248338
rect 197634 247888 197690 247897
rect 197634 247823 197690 247832
rect 197358 247344 197414 247353
rect 197358 247279 197414 247288
rect 197648 247110 197676 247823
rect 197636 247104 197688 247110
rect 197636 247046 197688 247052
rect 197360 247036 197412 247042
rect 197360 246978 197412 246984
rect 197372 245993 197400 246978
rect 197358 245984 197414 245993
rect 197358 245919 197414 245928
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243817 197400 244190
rect 197452 244180 197504 244186
rect 197452 244122 197504 244128
rect 197358 243808 197414 243817
rect 197358 243743 197414 243752
rect 197464 243001 197492 244122
rect 197450 242992 197506 243001
rect 197450 242927 197506 242936
rect 197360 242888 197412 242894
rect 197360 242830 197412 242836
rect 197372 241641 197400 242830
rect 197450 242176 197506 242185
rect 197450 242111 197506 242120
rect 197358 241632 197414 241641
rect 197358 241567 197414 241576
rect 197464 241534 197492 242111
rect 197452 241528 197504 241534
rect 197452 241470 197504 241476
rect 198384 225593 198412 251631
rect 198462 246528 198518 246537
rect 198462 246463 198518 246472
rect 198370 225584 198426 225593
rect 198370 225519 198426 225528
rect 198476 196654 198504 246463
rect 198464 196648 198516 196654
rect 198464 196590 198516 196596
rect 198568 181393 198596 252991
rect 198554 181384 198610 181393
rect 198554 181319 198610 181328
rect 197266 178664 197322 178673
rect 197266 178599 197322 178608
rect 198660 177342 198688 263055
rect 199750 245168 199806 245177
rect 199750 245103 199806 245112
rect 199106 241496 199162 241505
rect 199106 241431 199162 241440
rect 199120 240242 199148 241431
rect 199108 240236 199160 240242
rect 199108 240178 199160 240184
rect 199764 238754 199792 245103
rect 199842 244352 199898 244361
rect 199842 244287 199898 244296
rect 199856 239562 199884 244287
rect 199844 239556 199896 239562
rect 199844 239498 199896 239504
rect 199764 238726 199884 238754
rect 199856 195362 199884 238726
rect 199844 195356 199896 195362
rect 199844 195298 199896 195304
rect 199948 184346 199976 285670
rect 199936 184340 199988 184346
rect 199936 184282 199988 184288
rect 200040 180198 200068 285738
rect 200408 284036 200436 289138
rect 201316 287224 201368 287230
rect 201316 287166 201368 287172
rect 200946 284064 201002 284073
rect 200790 284022 200946 284050
rect 201328 284036 201356 287166
rect 201684 287156 201736 287162
rect 201684 287098 201736 287104
rect 201500 284232 201552 284238
rect 201406 284200 201462 284209
rect 201462 284180 201500 284186
rect 201462 284174 201552 284180
rect 201462 284158 201540 284174
rect 201406 284135 201462 284144
rect 201696 284036 201724 287098
rect 202156 284238 202184 660282
rect 202800 294710 202828 703520
rect 215944 700324 215996 700330
rect 215944 700266 215996 700272
rect 204904 448588 204956 448594
rect 204904 448530 204956 448536
rect 202788 294704 202840 294710
rect 202788 294646 202840 294652
rect 204260 289128 204312 289134
rect 204260 289070 204312 289076
rect 202234 288552 202290 288561
rect 202234 288487 202290 288496
rect 202144 284232 202196 284238
rect 202144 284174 202196 284180
rect 202248 284036 202276 288487
rect 202788 287088 202840 287094
rect 202788 287030 202840 287036
rect 202800 284036 202828 287030
rect 203156 286068 203208 286074
rect 203156 286010 203208 286016
rect 203168 284036 203196 286010
rect 203708 285864 203760 285870
rect 203708 285806 203760 285812
rect 203720 284036 203748 285806
rect 204272 284036 204300 289070
rect 204628 286000 204680 286006
rect 204628 285942 204680 285948
rect 204640 284036 204668 285942
rect 204916 285734 204944 448530
rect 206284 404388 206336 404394
rect 206284 404330 206336 404336
rect 206296 289202 206324 404330
rect 209044 382968 209096 382974
rect 209044 382910 209096 382916
rect 206284 289196 206336 289202
rect 206284 289138 206336 289144
rect 206652 288448 206704 288454
rect 206652 288390 206704 288396
rect 206100 285932 206152 285938
rect 206100 285874 206152 285880
rect 205548 285796 205600 285802
rect 205548 285738 205600 285744
rect 204904 285728 204956 285734
rect 204904 285670 204956 285676
rect 205560 284036 205588 285738
rect 206112 284036 206140 285874
rect 206664 284036 206692 288390
rect 207570 287192 207626 287201
rect 207570 287127 207626 287136
rect 207020 285864 207072 285870
rect 207020 285806 207072 285812
rect 207032 284036 207060 285806
rect 207584 284036 207612 287127
rect 208492 286408 208544 286414
rect 208492 286350 208544 286356
rect 208124 285728 208176 285734
rect 208124 285670 208176 285676
rect 208136 284036 208164 285670
rect 208504 284036 208532 286350
rect 209056 284036 209084 382910
rect 214564 298784 214616 298790
rect 214564 298726 214616 298732
rect 209688 296744 209740 296750
rect 209688 296686 209740 296692
rect 209700 284050 209728 296686
rect 213828 294636 213880 294642
rect 213828 294578 213880 294584
rect 211068 291848 211120 291854
rect 211068 291790 211120 291796
rect 210884 286340 210936 286346
rect 210884 286282 210936 286288
rect 209964 285728 210016 285734
rect 209964 285670 210016 285676
rect 209438 284022 209728 284050
rect 209976 284036 210004 285670
rect 210896 284036 210924 286282
rect 211080 285734 211108 291790
rect 211986 285832 212042 285841
rect 211986 285767 212042 285776
rect 213460 285796 213512 285802
rect 211068 285728 211120 285734
rect 211068 285670 211120 285676
rect 212000 284036 212028 285767
rect 213460 285738 213512 285744
rect 212908 285728 212960 285734
rect 212908 285670 212960 285676
rect 212356 284572 212408 284578
rect 212356 284514 212408 284520
rect 212368 284036 212396 284514
rect 212920 284036 212948 285670
rect 213472 284036 213500 285738
rect 213840 285734 213868 294578
rect 214576 285802 214604 298726
rect 215208 290012 215260 290018
rect 215208 289954 215260 289960
rect 214564 285796 214616 285802
rect 214564 285738 214616 285744
rect 214748 285796 214800 285802
rect 214748 285738 214800 285744
rect 213828 285728 213880 285734
rect 213828 285670 213880 285676
rect 214380 285728 214432 285734
rect 214380 285670 214432 285676
rect 213828 284436 213880 284442
rect 213828 284378 213880 284384
rect 213840 284036 213868 284378
rect 214392 284036 214420 285670
rect 214760 284036 214788 285738
rect 215220 285734 215248 289954
rect 215956 289814 215984 700266
rect 218992 699825 219020 703520
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 252560 700392 252612 700398
rect 252560 700334 252612 700340
rect 238024 700324 238076 700330
rect 238024 700266 238076 700272
rect 218978 699816 219034 699825
rect 218978 699751 219034 699760
rect 222844 696244 222896 696250
rect 222844 696186 222896 696192
rect 220084 605872 220136 605878
rect 220084 605814 220136 605820
rect 219348 292732 219400 292738
rect 219348 292674 219400 292680
rect 216586 291272 216642 291281
rect 216586 291207 216642 291216
rect 216496 290080 216548 290086
rect 216496 290022 216548 290028
rect 215944 289808 215996 289814
rect 215944 289750 215996 289756
rect 215208 285728 215260 285734
rect 215208 285670 215260 285676
rect 215300 285728 215352 285734
rect 215300 285670 215352 285676
rect 215312 284036 215340 285670
rect 215852 284980 215904 284986
rect 215852 284922 215904 284928
rect 215864 284036 215892 284922
rect 216508 284050 216536 290022
rect 216600 285734 216628 291207
rect 218244 289808 218296 289814
rect 218244 289750 218296 289756
rect 216588 285728 216640 285734
rect 216588 285670 216640 285676
rect 217322 285696 217378 285705
rect 217322 285631 217378 285640
rect 217046 284064 217102 284073
rect 216246 284022 216536 284050
rect 216798 284022 217046 284050
rect 200946 283999 201002 284008
rect 217336 284036 217364 285631
rect 218256 284036 218284 289750
rect 218612 286476 218664 286482
rect 218612 286418 218664 286424
rect 218624 284036 218652 286418
rect 219360 284050 219388 292674
rect 219714 288688 219770 288697
rect 219714 288623 219770 288632
rect 219190 284022 219388 284050
rect 219728 284036 219756 288623
rect 220096 288386 220124 605814
rect 220084 288380 220136 288386
rect 220084 288322 220136 288328
rect 222108 287088 222160 287094
rect 222108 287030 222160 287036
rect 220634 286104 220690 286113
rect 220634 286039 220690 286048
rect 220082 284336 220138 284345
rect 220082 284271 220138 284280
rect 220096 284036 220124 284271
rect 220648 284036 220676 286039
rect 221186 285968 221242 285977
rect 221186 285903 221242 285912
rect 221200 285802 221228 285903
rect 221188 285796 221240 285802
rect 221188 285738 221240 285744
rect 221556 285796 221608 285802
rect 221556 285738 221608 285744
rect 221188 284708 221240 284714
rect 221188 284650 221240 284656
rect 221200 284036 221228 284650
rect 221568 284036 221596 285738
rect 222120 284036 222148 287030
rect 222856 286482 222884 696186
rect 226984 579692 227036 579698
rect 226984 579634 227036 579640
rect 224224 318844 224276 318850
rect 224224 318786 224276 318792
rect 224236 291990 224264 318786
rect 226248 300144 226300 300150
rect 226248 300086 226300 300092
rect 224224 291984 224276 291990
rect 224224 291926 224276 291932
rect 224868 291304 224920 291310
rect 224868 291246 224920 291252
rect 223394 290456 223450 290465
rect 223394 290391 223450 290400
rect 222844 286476 222896 286482
rect 222844 286418 222896 286424
rect 223408 284050 223436 290391
rect 224880 285734 224908 291246
rect 225420 288380 225472 288386
rect 225420 288322 225472 288328
rect 223580 285728 223632 285734
rect 223580 285670 223632 285676
rect 224868 285728 224920 285734
rect 224868 285670 224920 285676
rect 223054 284022 223436 284050
rect 223592 284036 223620 285670
rect 223948 284504 224000 284510
rect 223948 284446 224000 284452
rect 223960 284036 223988 284446
rect 225432 284036 225460 288322
rect 226260 284050 226288 300086
rect 226996 290601 227024 579634
rect 233884 501016 233936 501022
rect 233884 500958 233936 500964
rect 232504 345092 232556 345098
rect 232504 345034 232556 345040
rect 228364 338768 228416 338774
rect 228364 338710 228416 338716
rect 227628 294024 227680 294030
rect 227628 293966 227680 293972
rect 226982 290592 227038 290601
rect 226982 290527 227038 290536
rect 227640 285734 227668 293966
rect 227812 285864 227864 285870
rect 227812 285806 227864 285812
rect 226524 285728 226576 285734
rect 226524 285670 226576 285676
rect 227628 285728 227680 285734
rect 227628 285670 227680 285676
rect 225998 284022 226288 284050
rect 226536 284036 226564 285670
rect 227444 284368 227496 284374
rect 227444 284310 227496 284316
rect 227456 284036 227484 284310
rect 227824 284036 227852 285806
rect 228376 284036 228404 338710
rect 232516 290494 232544 345034
rect 232596 292664 232648 292670
rect 232596 292606 232648 292612
rect 232504 290488 232556 290494
rect 232504 290430 232556 290436
rect 229836 287428 229888 287434
rect 229836 287370 229888 287376
rect 228914 284472 228970 284481
rect 228914 284407 228970 284416
rect 228928 284036 228956 284407
rect 229848 284036 229876 287370
rect 230388 287292 230440 287298
rect 230388 287234 230440 287240
rect 230400 284036 230428 287234
rect 232608 286414 232636 292606
rect 232780 290556 232832 290562
rect 232780 290498 232832 290504
rect 232596 286408 232648 286414
rect 232596 286350 232648 286356
rect 231676 286068 231728 286074
rect 231676 286010 231728 286016
rect 231582 284064 231638 284073
rect 231334 284022 231582 284050
rect 217046 283999 217102 284008
rect 231688 284036 231716 286010
rect 232228 285932 232280 285938
rect 232228 285874 232280 285880
rect 232240 284036 232268 285874
rect 232792 284036 232820 290498
rect 233896 289134 233924 500958
rect 235724 295996 235776 296002
rect 235724 295938 235776 295944
rect 233884 289128 233936 289134
rect 233884 289070 233936 289076
rect 233148 287292 233200 287298
rect 233148 287234 233200 287240
rect 233160 284036 233188 287234
rect 235736 285802 235764 295938
rect 236920 292596 236972 292602
rect 236920 292538 236972 292544
rect 235816 289944 235868 289950
rect 235816 289886 235868 289892
rect 234620 285796 234672 285802
rect 234620 285738 234672 285744
rect 235724 285796 235776 285802
rect 235724 285738 235776 285744
rect 233698 284336 233754 284345
rect 233698 284271 233754 284280
rect 233712 284036 233740 284271
rect 234632 284036 234660 285738
rect 235828 284322 235856 289886
rect 236644 288652 236696 288658
rect 236644 288594 236696 288600
rect 235908 288380 235960 288386
rect 235908 288322 235960 288328
rect 235460 284294 235856 284322
rect 235460 284050 235488 284294
rect 235920 284050 235948 288322
rect 236656 286346 236684 288594
rect 236644 286340 236696 286346
rect 236644 286282 236696 286288
rect 236092 286000 236144 286006
rect 236092 285942 236144 285948
rect 235198 284022 235488 284050
rect 235566 284022 235948 284050
rect 236104 284036 236132 285942
rect 236932 284050 236960 292538
rect 237380 288516 237432 288522
rect 237380 288458 237432 288464
rect 237392 284986 237420 288458
rect 238036 288386 238064 700266
rect 249064 698964 249116 698970
rect 249064 698906 249116 698912
rect 240508 665848 240560 665854
rect 240508 665790 240560 665796
rect 240140 291984 240192 291990
rect 240140 291926 240192 291932
rect 239956 289876 240008 289882
rect 239956 289818 240008 289824
rect 238024 288380 238076 288386
rect 238024 288322 238076 288328
rect 239588 287360 239640 287366
rect 239588 287302 239640 287308
rect 238482 286104 238538 286113
rect 238482 286039 238538 286048
rect 237380 284980 237432 284986
rect 237380 284922 237432 284928
rect 237012 284640 237064 284646
rect 237012 284582 237064 284588
rect 236670 284022 236960 284050
rect 237024 284036 237052 284582
rect 238116 284504 238168 284510
rect 238116 284446 238168 284452
rect 237564 284436 237616 284442
rect 237564 284378 237616 284384
rect 237576 284036 237604 284378
rect 238128 284036 238156 284446
rect 238496 284036 238524 286039
rect 239036 285796 239088 285802
rect 239036 285738 239088 285744
rect 239048 284036 239076 285738
rect 239600 284036 239628 287302
rect 239968 285802 239996 289818
rect 239956 285796 240008 285802
rect 239956 285738 240008 285744
rect 240152 285326 240180 291926
rect 240140 285320 240192 285326
rect 240140 285262 240192 285268
rect 239956 284368 240008 284374
rect 239956 284310 240008 284316
rect 239968 284036 239996 284310
rect 240520 284036 240548 665790
rect 244924 474768 244976 474774
rect 244924 474710 244976 474716
rect 244280 294704 244332 294710
rect 244280 294646 244332 294652
rect 242716 291236 242768 291242
rect 242716 291178 242768 291184
rect 240876 288584 240928 288590
rect 240876 288526 240928 288532
rect 240888 284036 240916 288526
rect 241980 285796 242032 285802
rect 241980 285738 242032 285744
rect 241060 285320 241112 285326
rect 241060 285262 241112 285268
rect 241072 284050 241100 285262
rect 241072 284022 241454 284050
rect 241992 284036 242020 285738
rect 242728 284050 242756 291178
rect 243820 290488 243872 290494
rect 243820 290430 243872 290436
rect 242900 290148 242952 290154
rect 242900 290090 242952 290096
rect 242374 284022 242756 284050
rect 242912 284036 242940 290090
rect 243634 284064 243690 284073
rect 243478 284022 243634 284050
rect 231582 283999 231638 284008
rect 243832 284036 243860 290430
rect 244004 286068 244056 286074
rect 244004 286010 244056 286016
rect 243634 283999 243690 284008
rect 234528 283960 234580 283966
rect 204902 283928 204958 283937
rect 210698 283928 210754 283937
rect 204958 283886 205206 283914
rect 210542 283886 210698 283914
rect 204902 283863 204958 283872
rect 211710 283928 211766 283937
rect 211462 283886 211710 283914
rect 210698 283863 210754 283872
rect 211710 283863 211766 283872
rect 217598 283928 217654 283937
rect 222658 283928 222714 283937
rect 217654 283886 217718 283914
rect 222502 283886 222658 283914
rect 217598 283863 217654 283872
rect 222658 283863 222714 283872
rect 224222 283928 224278 283937
rect 225234 283928 225290 283937
rect 224278 283886 224526 283914
rect 225078 283886 225234 283914
rect 224222 283863 224278 283872
rect 225234 283863 225290 283872
rect 226614 283928 226670 283937
rect 229466 283928 229522 283937
rect 226670 283886 226918 283914
rect 229310 283886 229466 283914
rect 226614 283863 226670 283872
rect 231030 283928 231086 283937
rect 230782 283886 231030 283914
rect 229466 283863 229522 283872
rect 234278 283908 234528 283914
rect 234278 283902 234580 283908
rect 234278 283886 234568 283902
rect 231030 283863 231086 283872
rect 244016 279721 244044 286010
rect 244096 284436 244148 284442
rect 244096 284378 244148 284384
rect 244108 283626 244136 284378
rect 244096 283620 244148 283626
rect 244096 283562 244148 283568
rect 244002 279712 244058 279721
rect 244002 279647 244058 279656
rect 244292 278905 244320 294646
rect 244278 278896 244334 278905
rect 244278 278831 244334 278840
rect 244278 260944 244334 260953
rect 244278 260879 244334 260888
rect 244186 244216 244242 244225
rect 244186 244151 244242 244160
rect 244096 241528 244148 241534
rect 244096 241470 244148 241476
rect 200224 237726 200252 240244
rect 200212 237720 200264 237726
rect 200212 237662 200264 237668
rect 200592 237454 200620 240244
rect 201144 237590 201172 240244
rect 201512 237794 201540 240244
rect 201500 237788 201552 237794
rect 201500 237730 201552 237736
rect 201316 237720 201368 237726
rect 201316 237662 201368 237668
rect 201132 237584 201184 237590
rect 201132 237526 201184 237532
rect 200580 237448 200632 237454
rect 200580 237390 200632 237396
rect 201328 215966 201356 237662
rect 201408 237448 201460 237454
rect 201408 237390 201460 237396
rect 201316 215960 201368 215966
rect 201316 215902 201368 215908
rect 200028 180192 200080 180198
rect 200028 180134 200080 180140
rect 201420 180130 201448 237390
rect 202064 235958 202092 240244
rect 202052 235952 202104 235958
rect 202052 235894 202104 235900
rect 202616 181490 202644 240244
rect 202696 237788 202748 237794
rect 202696 237730 202748 237736
rect 202708 221474 202736 237730
rect 202984 237522 203012 240244
rect 202972 237516 203024 237522
rect 202972 237458 203024 237464
rect 203536 237454 203564 240244
rect 204088 238754 204116 240244
rect 204088 238726 204208 238754
rect 203892 237516 203944 237522
rect 203892 237458 203944 237464
rect 203524 237448 203576 237454
rect 203524 237390 203576 237396
rect 202696 221468 202748 221474
rect 202696 221410 202748 221416
rect 203904 188358 203932 237458
rect 203984 237448 204036 237454
rect 203984 237390 204036 237396
rect 203996 227050 204024 237390
rect 203984 227044 204036 227050
rect 203984 226986 204036 226992
rect 203892 188352 203944 188358
rect 203892 188294 203944 188300
rect 204180 187134 204208 238726
rect 204456 237425 204484 240244
rect 204718 240136 204774 240145
rect 204718 240071 204774 240080
rect 204732 238754 204760 240071
rect 204732 238726 204944 238754
rect 204442 237416 204498 237425
rect 204442 237351 204498 237360
rect 204916 200802 204944 238726
rect 205008 231130 205036 240244
rect 205376 238754 205404 240244
rect 205546 240136 205602 240145
rect 205546 240071 205602 240080
rect 205376 238726 205496 238754
rect 204996 231124 205048 231130
rect 204996 231066 205048 231072
rect 205468 203590 205496 238726
rect 205456 203584 205508 203590
rect 205456 203526 205508 203532
rect 204904 200796 204956 200802
rect 204904 200738 204956 200744
rect 204168 187128 204220 187134
rect 204168 187070 204220 187076
rect 202604 181484 202656 181490
rect 202604 181426 202656 181432
rect 203524 180872 203576 180878
rect 203524 180814 203576 180820
rect 201408 180124 201460 180130
rect 201408 180066 201460 180072
rect 200764 178084 200816 178090
rect 200764 178026 200816 178032
rect 198648 177336 198700 177342
rect 198648 177278 198700 177284
rect 198096 176860 198148 176866
rect 198096 176802 198148 176808
rect 194508 175092 194560 175098
rect 194508 175034 194560 175040
rect 191104 159996 191156 160002
rect 191104 159938 191156 159944
rect 184296 151904 184348 151910
rect 184296 151846 184348 151852
rect 184204 150408 184256 150414
rect 184204 150350 184256 150356
rect 184204 144968 184256 144974
rect 184204 144910 184256 144916
rect 182824 135924 182876 135930
rect 182824 135866 182876 135872
rect 181444 135312 181496 135318
rect 181444 135254 181496 135260
rect 180156 104916 180208 104922
rect 180156 104858 180208 104864
rect 180168 93809 180196 104858
rect 180154 93800 180210 93809
rect 180154 93735 180210 93744
rect 181456 86698 181484 135254
rect 181536 116000 181588 116006
rect 181536 115942 181588 115948
rect 181548 93974 181576 115942
rect 181536 93968 181588 93974
rect 181536 93910 181588 93916
rect 182836 92274 182864 135866
rect 182916 106344 182968 106350
rect 182916 106286 182968 106292
rect 182824 92268 182876 92274
rect 182824 92210 182876 92216
rect 182928 90982 182956 106286
rect 182916 90976 182968 90982
rect 182916 90918 182968 90924
rect 181444 86692 181496 86698
rect 181444 86634 181496 86640
rect 184216 83910 184244 144910
rect 184308 93430 184336 151846
rect 198004 150476 198056 150482
rect 198004 150418 198056 150424
rect 195244 146328 195296 146334
rect 195244 146270 195296 146276
rect 191104 145036 191156 145042
rect 191104 144978 191156 144984
rect 188344 143608 188396 143614
rect 188344 143550 188396 143556
rect 186964 142180 187016 142186
rect 186964 142122 187016 142128
rect 185584 138032 185636 138038
rect 185584 137974 185636 137980
rect 184388 104984 184440 104990
rect 184388 104926 184440 104932
rect 184296 93424 184348 93430
rect 184296 93366 184348 93372
rect 184400 89729 184428 104926
rect 185596 94042 185624 137974
rect 185676 114640 185728 114646
rect 185676 114582 185728 114588
rect 185584 94036 185636 94042
rect 185584 93978 185636 93984
rect 185688 90846 185716 114582
rect 185676 90840 185728 90846
rect 185676 90782 185728 90788
rect 184386 89720 184442 89729
rect 184386 89655 184442 89664
rect 184296 86284 184348 86290
rect 184296 86226 184348 86232
rect 184204 83904 184256 83910
rect 184204 83846 184256 83852
rect 180064 82544 180116 82550
rect 180064 82486 180116 82492
rect 184308 42158 184336 86226
rect 186976 78538 187004 142122
rect 187148 139460 187200 139466
rect 187148 139402 187200 139408
rect 187056 90432 187108 90438
rect 187056 90374 187108 90380
rect 186964 78532 187016 78538
rect 186964 78474 187016 78480
rect 184296 42152 184348 42158
rect 184296 42094 184348 42100
rect 187068 32434 187096 90374
rect 187160 82618 187188 139402
rect 187148 82612 187200 82618
rect 187148 82554 187200 82560
rect 188356 79966 188384 143550
rect 189724 140888 189776 140894
rect 189724 140830 189776 140836
rect 189736 88233 189764 140830
rect 189816 117428 189868 117434
rect 189816 117370 189868 117376
rect 189722 88224 189778 88233
rect 189722 88159 189778 88168
rect 189828 86834 189856 117370
rect 189816 86828 189868 86834
rect 189816 86770 189868 86776
rect 188344 79960 188396 79966
rect 188344 79902 188396 79908
rect 191116 77178 191144 144978
rect 193956 125724 194008 125730
rect 193956 125666 194008 125672
rect 193864 118788 193916 118794
rect 193864 118730 193916 118736
rect 192484 118720 192536 118726
rect 192484 118662 192536 118668
rect 191288 107772 191340 107778
rect 191288 107714 191340 107720
rect 191196 87644 191248 87650
rect 191196 87586 191248 87592
rect 191104 77172 191156 77178
rect 191104 77114 191156 77120
rect 191208 40730 191236 87586
rect 191300 84114 191328 107714
rect 192496 88194 192524 118662
rect 192484 88188 192536 88194
rect 192484 88130 192536 88136
rect 193876 85270 193904 118730
rect 193968 93362 193996 125666
rect 193956 93356 194008 93362
rect 193956 93298 194008 93304
rect 193864 85264 193916 85270
rect 193864 85206 193916 85212
rect 191288 84108 191340 84114
rect 191288 84050 191340 84056
rect 195256 75818 195284 146270
rect 195428 124296 195480 124302
rect 195428 124238 195480 124244
rect 195336 93220 195388 93226
rect 195336 93162 195388 93168
rect 195244 75812 195296 75818
rect 195244 75754 195296 75760
rect 191196 40724 191248 40730
rect 191196 40666 191248 40672
rect 187056 32428 187108 32434
rect 187056 32370 187108 32376
rect 195348 28354 195376 93162
rect 195440 92342 195468 124238
rect 196808 120148 196860 120154
rect 196808 120090 196860 120096
rect 196716 113212 196768 113218
rect 196716 113154 196768 113160
rect 195520 102196 195572 102202
rect 195520 102138 195572 102144
rect 195428 92336 195480 92342
rect 195428 92278 195480 92284
rect 195532 81394 195560 102138
rect 196624 96892 196676 96898
rect 196624 96834 196676 96840
rect 195520 81388 195572 81394
rect 195520 81330 195572 81336
rect 195336 28348 195388 28354
rect 195336 28290 195388 28296
rect 196636 19990 196664 96834
rect 196728 88262 196756 113154
rect 196820 93906 196848 120090
rect 198016 111790 198044 150418
rect 198108 150346 198136 176802
rect 200776 166870 200804 178026
rect 200764 166864 200816 166870
rect 200764 166806 200816 166812
rect 203536 157350 203564 180814
rect 203524 157344 203576 157350
rect 203524 157286 203576 157292
rect 200764 151088 200816 151094
rect 200764 151030 200816 151036
rect 198096 150340 198148 150346
rect 198096 150282 198148 150288
rect 198096 143676 198148 143682
rect 198096 143618 198148 143624
rect 198004 111784 198056 111790
rect 198004 111726 198056 111732
rect 196808 93900 196860 93906
rect 196808 93842 196860 93848
rect 198004 89140 198056 89146
rect 198004 89082 198056 89088
rect 196716 88256 196768 88262
rect 196716 88198 196768 88204
rect 196624 19984 196676 19990
rect 196624 19926 196676 19932
rect 198016 6254 198044 89082
rect 198108 81326 198136 143618
rect 198188 109132 198240 109138
rect 198188 109074 198240 109080
rect 198200 89622 198228 109074
rect 200776 109002 200804 151030
rect 202144 146396 202196 146402
rect 202144 146338 202196 146344
rect 200856 113280 200908 113286
rect 200856 113222 200908 113228
rect 200764 108996 200816 109002
rect 200764 108938 200816 108944
rect 199384 106412 199436 106418
rect 199384 106354 199436 106360
rect 198188 89616 198240 89622
rect 198188 89558 198240 89564
rect 199396 85542 199424 106354
rect 200764 91996 200816 92002
rect 200764 91938 200816 91944
rect 199384 85536 199436 85542
rect 199384 85478 199436 85484
rect 198096 81320 198148 81326
rect 198096 81262 198148 81268
rect 200776 43450 200804 91938
rect 200868 91050 200896 113222
rect 200856 91044 200908 91050
rect 200856 90986 200908 90992
rect 202156 78606 202184 146338
rect 204996 128444 205048 128450
rect 204996 128386 205048 128392
rect 202328 127084 202380 127090
rect 202328 127026 202380 127032
rect 202236 89004 202288 89010
rect 202236 88946 202288 88952
rect 202144 78600 202196 78606
rect 202144 78542 202196 78548
rect 200764 43444 200816 43450
rect 200764 43386 200816 43392
rect 202248 37942 202276 88946
rect 202340 85474 202368 127026
rect 203524 121508 203576 121514
rect 203524 121450 203576 121456
rect 202328 85468 202380 85474
rect 202328 85410 202380 85416
rect 203536 85406 203564 121450
rect 203616 98116 203668 98122
rect 203616 98058 203668 98064
rect 203524 85400 203576 85406
rect 203524 85342 203576 85348
rect 203628 74526 203656 98058
rect 204904 93288 204956 93294
rect 204904 93230 204956 93236
rect 203616 74520 203668 74526
rect 203616 74462 203668 74468
rect 202236 37936 202288 37942
rect 202236 37878 202288 37884
rect 204916 35222 204944 93230
rect 205008 82754 205036 128386
rect 205560 96422 205588 240071
rect 205928 237726 205956 240244
rect 206480 238270 206508 240244
rect 206468 238264 206520 238270
rect 206468 238206 206520 238212
rect 205916 237720 205968 237726
rect 205916 237662 205968 237668
rect 206744 237720 206796 237726
rect 206744 237662 206796 237668
rect 206756 185609 206784 237662
rect 206742 185600 206798 185609
rect 206742 185535 206798 185544
rect 206848 184482 206876 240244
rect 206928 238264 206980 238270
rect 206928 238206 206980 238212
rect 206836 184476 206888 184482
rect 206836 184418 206888 184424
rect 206940 178906 206968 238206
rect 207400 237726 207428 240244
rect 207952 239494 207980 240244
rect 207940 239488 207992 239494
rect 207940 239430 207992 239436
rect 207388 237720 207440 237726
rect 207388 237662 207440 237668
rect 208216 237720 208268 237726
rect 208216 237662 208268 237668
rect 208228 210458 208256 237662
rect 208216 210452 208268 210458
rect 208216 210394 208268 210400
rect 206928 178900 206980 178906
rect 206928 178842 206980 178848
rect 206282 178120 206338 178129
rect 206282 178055 206338 178064
rect 205548 96416 205600 96422
rect 205548 96358 205600 96364
rect 206296 96354 206324 178055
rect 208320 177410 208348 240244
rect 208872 238649 208900 240244
rect 209136 239556 209188 239562
rect 209136 239498 209188 239504
rect 208858 238640 208914 238649
rect 208858 238575 208914 238584
rect 209044 237584 209096 237590
rect 209044 237526 209096 237532
rect 208400 237448 208452 237454
rect 208400 237390 208452 237396
rect 208412 233918 208440 237390
rect 208400 233912 208452 233918
rect 208400 233854 208452 233860
rect 208308 177404 208360 177410
rect 208308 177346 208360 177352
rect 207664 176928 207716 176934
rect 207664 176870 207716 176876
rect 207676 149054 207704 176870
rect 209056 174554 209084 237526
rect 209148 203658 209176 239498
rect 209240 238610 209268 240244
rect 209792 239578 209820 240244
rect 209792 239550 209912 239578
rect 209780 239420 209832 239426
rect 209780 239362 209832 239368
rect 209792 238746 209820 239362
rect 209780 238740 209832 238746
rect 209780 238682 209832 238688
rect 209228 238604 209280 238610
rect 209228 238546 209280 238552
rect 209884 233918 209912 239550
rect 210344 237454 210372 240244
rect 210712 238754 210740 240244
rect 210712 238726 211108 238754
rect 210332 237448 210384 237454
rect 210332 237390 210384 237396
rect 209872 233912 209924 233918
rect 209872 233854 209924 233860
rect 209136 203652 209188 203658
rect 209136 203594 209188 203600
rect 211080 192545 211108 238726
rect 211264 238134 211292 240244
rect 211252 238128 211304 238134
rect 211252 238070 211304 238076
rect 211816 237454 211844 240244
rect 211804 237448 211856 237454
rect 211804 237390 211856 237396
rect 212184 235278 212212 240244
rect 212736 240038 212764 240244
rect 212724 240032 212776 240038
rect 212724 239974 212776 239980
rect 213104 237454 213132 240244
rect 213184 240168 213236 240174
rect 213184 240110 213236 240116
rect 212448 237448 212500 237454
rect 212448 237390 212500 237396
rect 213092 237448 213144 237454
rect 213092 237390 213144 237396
rect 212172 235272 212224 235278
rect 212172 235214 212224 235220
rect 211066 192536 211122 192545
rect 211066 192471 211122 192480
rect 212460 178974 212488 237390
rect 212448 178968 212500 178974
rect 212448 178910 212500 178916
rect 212446 178800 212502 178809
rect 212446 178735 212502 178744
rect 209044 174548 209096 174554
rect 209044 174490 209096 174496
rect 207664 149048 207716 149054
rect 207664 148990 207716 148996
rect 206376 139528 206428 139534
rect 206376 139470 206428 139476
rect 206284 96348 206336 96354
rect 206284 96290 206336 96296
rect 206284 91928 206336 91934
rect 206284 91870 206336 91876
rect 204996 82748 205048 82754
rect 204996 82690 205048 82696
rect 206296 50386 206324 91870
rect 206388 82686 206416 139470
rect 209136 135380 209188 135386
rect 209136 135322 209188 135328
rect 206468 121576 206520 121582
rect 206468 121518 206520 121524
rect 206480 93158 206508 121518
rect 207664 120216 207716 120222
rect 207664 120158 207716 120164
rect 206560 96960 206612 96966
rect 206560 96902 206612 96908
rect 206468 93152 206520 93158
rect 206468 93094 206520 93100
rect 206376 82680 206428 82686
rect 206376 82622 206428 82628
rect 206572 71738 206600 96902
rect 207676 89554 207704 120158
rect 207664 89548 207716 89554
rect 207664 89490 207716 89496
rect 209044 87780 209096 87786
rect 209044 87722 209096 87728
rect 206560 71732 206612 71738
rect 206560 71674 206612 71680
rect 206284 50380 206336 50386
rect 206284 50322 206336 50328
rect 204904 35216 204956 35222
rect 204904 35158 204956 35164
rect 209056 13122 209084 87722
rect 209148 84046 209176 135322
rect 210424 129872 210476 129878
rect 210424 129814 210476 129820
rect 209228 118856 209280 118862
rect 209228 118798 209280 118804
rect 209240 86970 209268 118798
rect 209320 96824 209372 96830
rect 209320 96766 209372 96772
rect 209228 86964 209280 86970
rect 209228 86906 209280 86912
rect 209136 84040 209188 84046
rect 209136 83982 209188 83988
rect 209332 82822 209360 96766
rect 210436 84182 210464 129814
rect 211804 111920 211856 111926
rect 211804 111862 211856 111868
rect 211816 89690 211844 111862
rect 211896 95260 211948 95266
rect 211896 95202 211948 95208
rect 211804 89684 211856 89690
rect 211804 89626 211856 89632
rect 211804 84856 211856 84862
rect 211804 84798 211856 84804
rect 210424 84176 210476 84182
rect 210424 84118 210476 84124
rect 209320 82816 209372 82822
rect 209320 82758 209372 82764
rect 211816 24138 211844 84798
rect 211908 75886 211936 95202
rect 212460 95198 212488 178735
rect 212448 95192 212500 95198
rect 212448 95134 212500 95140
rect 213196 93838 213224 240110
rect 213656 238754 213684 240244
rect 213656 238726 213868 238754
rect 213736 237448 213788 237454
rect 213736 237390 213788 237396
rect 213748 206281 213776 237390
rect 213734 206272 213790 206281
rect 213734 206207 213790 206216
rect 213840 184550 213868 238726
rect 214208 238066 214236 240244
rect 214576 238746 214604 240244
rect 215128 238754 215156 240244
rect 214564 238740 214616 238746
rect 215128 238726 215248 238754
rect 214564 238682 214616 238688
rect 214196 238060 214248 238066
rect 214196 238002 214248 238008
rect 215024 238060 215076 238066
rect 215024 238002 215076 238008
rect 214564 203652 214616 203658
rect 214564 203594 214616 203600
rect 214576 189990 214604 203594
rect 215036 202162 215064 238002
rect 215024 202156 215076 202162
rect 215024 202098 215076 202104
rect 214564 189984 214616 189990
rect 214564 189926 214616 189932
rect 213828 184544 213880 184550
rect 213828 184486 213880 184492
rect 215220 180266 215248 238726
rect 215680 237454 215708 240244
rect 216048 238610 216076 240244
rect 216036 238604 216088 238610
rect 216036 238546 216088 238552
rect 216600 238542 216628 240244
rect 216588 238536 216640 238542
rect 216588 238478 216640 238484
rect 215668 237448 215720 237454
rect 215668 237390 215720 237396
rect 216588 237448 216640 237454
rect 216588 237390 216640 237396
rect 216600 209001 216628 237390
rect 217152 236706 217180 240244
rect 217520 238754 217548 240244
rect 217520 238726 217916 238754
rect 217140 236700 217192 236706
rect 217140 236642 217192 236648
rect 216586 208992 216642 209001
rect 216586 208927 216642 208936
rect 217888 195294 217916 238726
rect 218072 237522 218100 240244
rect 218060 237516 218112 237522
rect 218060 237458 218112 237464
rect 218440 237454 218468 240244
rect 218428 237448 218480 237454
rect 218428 237390 218480 237396
rect 218992 229838 219020 240244
rect 219346 240136 219402 240145
rect 219346 240071 219402 240080
rect 219256 237448 219308 237454
rect 219256 237390 219308 237396
rect 218980 229832 219032 229838
rect 218980 229774 219032 229780
rect 219268 204950 219296 237390
rect 219256 204944 219308 204950
rect 219256 204886 219308 204892
rect 217876 195288 217928 195294
rect 217876 195230 217928 195236
rect 215208 180260 215260 180266
rect 215208 180202 215260 180208
rect 214564 179444 214616 179450
rect 214564 179386 214616 179392
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173641 213960 173810
rect 214012 173800 214064 173806
rect 214012 173742 214064 173748
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173742
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 214012 172440 214064 172446
rect 214012 172382 214064 172388
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214024 171601 214052 172382
rect 214010 171592 214066 171601
rect 214010 171527 214066 171536
rect 213920 171080 213972 171086
rect 213918 171048 213920 171057
rect 213972 171048 213974 171057
rect 213918 170983 213974 170992
rect 214012 171012 214064 171018
rect 214012 170954 214064 170960
rect 214024 170377 214052 170954
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 213920 169720 213972 169726
rect 213918 169688 213920 169697
rect 213972 169688 213974 169697
rect 213918 169623 213974 169632
rect 214012 169652 214064 169658
rect 214012 169594 214064 169600
rect 214024 169017 214052 169594
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 214024 167657 214052 168234
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 214104 167000 214156 167006
rect 213918 166968 213974 166977
rect 214104 166942 214156 166948
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 213932 166870 213960 166903
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 214024 165753 214052 166874
rect 214116 166433 214144 166942
rect 214102 166424 214158 166433
rect 214102 166359 214158 166368
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 214012 165572 214064 165578
rect 214012 165514 214064 165520
rect 213920 165504 213972 165510
rect 213920 165446 213972 165452
rect 213932 165073 213960 165446
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165514
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163033 213960 164154
rect 214576 163713 214604 179386
rect 219360 177478 219388 240071
rect 219544 237386 219572 240244
rect 219912 237454 219940 240244
rect 220084 238128 220136 238134
rect 220084 238070 220136 238076
rect 219900 237448 219952 237454
rect 219900 237390 219952 237396
rect 219532 237380 219584 237386
rect 219532 237322 219584 237328
rect 220096 192506 220124 238070
rect 220464 238066 220492 240244
rect 220452 238060 220504 238066
rect 220452 238002 220504 238008
rect 220176 237516 220228 237522
rect 220176 237458 220228 237464
rect 220188 199442 220216 237458
rect 221016 237454 221044 240244
rect 220728 237448 220780 237454
rect 220728 237390 220780 237396
rect 221004 237448 221056 237454
rect 221004 237390 221056 237396
rect 220740 224262 220768 237390
rect 221384 237386 221412 240244
rect 221936 238474 221964 240244
rect 221924 238468 221976 238474
rect 221924 238410 221976 238416
rect 222016 237448 222068 237454
rect 222016 237390 222068 237396
rect 221372 237380 221424 237386
rect 221372 237322 221424 237328
rect 222028 227118 222056 237390
rect 222304 231198 222332 240244
rect 222856 237998 222884 240244
rect 222844 237992 222896 237998
rect 222844 237934 222896 237940
rect 222292 231192 222344 231198
rect 222292 231134 222344 231140
rect 222016 227112 222068 227118
rect 222016 227054 222068 227060
rect 220728 224256 220780 224262
rect 220728 224198 220780 224204
rect 220176 199436 220228 199442
rect 220176 199378 220228 199384
rect 220084 192500 220136 192506
rect 220084 192442 220136 192448
rect 223408 178022 223436 240244
rect 223776 238338 223804 240244
rect 224328 238754 224356 240244
rect 224328 238726 224724 238754
rect 223764 238332 223816 238338
rect 223764 238274 223816 238280
rect 223488 237992 223540 237998
rect 223488 237934 223540 237940
rect 223396 178016 223448 178022
rect 223396 177958 223448 177964
rect 219348 177472 219400 177478
rect 219348 177414 219400 177420
rect 223500 176050 223528 237934
rect 224696 218754 224724 238726
rect 224776 238332 224828 238338
rect 224776 238274 224828 238280
rect 224684 218748 224736 218754
rect 224684 218690 224736 218696
rect 224788 179042 224816 238274
rect 224776 179036 224828 179042
rect 224776 178978 224828 178984
rect 224880 176118 224908 240244
rect 225248 240106 225276 240244
rect 225236 240100 225288 240106
rect 225236 240042 225288 240048
rect 225800 237454 225828 240244
rect 225788 237448 225840 237454
rect 225788 237390 225840 237396
rect 226168 225622 226196 240244
rect 226720 237454 226748 240244
rect 226248 237448 226300 237454
rect 226248 237390 226300 237396
rect 226708 237448 226760 237454
rect 226708 237390 226760 237396
rect 226156 225616 226208 225622
rect 226156 225558 226208 225564
rect 226260 185638 226288 237390
rect 227272 234054 227300 240244
rect 227640 238474 227668 240244
rect 228192 238649 228220 240244
rect 228744 238754 228772 240244
rect 228744 238726 229048 238754
rect 228178 238640 228234 238649
rect 228178 238575 228234 238584
rect 227628 238468 227680 238474
rect 227628 238410 227680 238416
rect 227628 237448 227680 237454
rect 227628 237390 227680 237396
rect 227260 234048 227312 234054
rect 227260 233990 227312 233996
rect 227640 198014 227668 237390
rect 227628 198008 227680 198014
rect 227628 197950 227680 197956
rect 228364 189916 228416 189922
rect 228364 189858 228416 189864
rect 226248 185632 226300 185638
rect 226248 185574 226300 185580
rect 227626 180160 227682 180169
rect 227626 180095 227682 180104
rect 224868 176112 224920 176118
rect 224868 176054 224920 176060
rect 223488 176044 223540 176050
rect 223488 175986 223540 175992
rect 220910 175944 220966 175953
rect 220910 175879 220966 175888
rect 220924 175846 220952 175879
rect 220912 175840 220964 175846
rect 224224 175840 224276 175846
rect 220912 175782 220964 175788
rect 224222 175808 224224 175817
rect 227640 175817 227668 180095
rect 228376 176089 228404 189858
rect 229020 184278 229048 238726
rect 229112 235346 229140 240244
rect 229100 235340 229152 235346
rect 229100 235282 229152 235288
rect 229664 232558 229692 240244
rect 229742 240136 229798 240145
rect 229742 240071 229798 240080
rect 229652 232552 229704 232558
rect 229652 232494 229704 232500
rect 229008 184272 229060 184278
rect 229008 184214 229060 184220
rect 229468 178968 229520 178974
rect 229468 178910 229520 178916
rect 229192 178764 229244 178770
rect 229192 178706 229244 178712
rect 229098 177984 229154 177993
rect 229098 177919 229154 177928
rect 228362 176080 228418 176089
rect 228362 176015 228418 176024
rect 224276 175808 224278 175817
rect 224222 175743 224278 175752
rect 227626 175808 227682 175817
rect 227626 175743 227682 175752
rect 229008 175160 229060 175166
rect 229008 175102 229060 175108
rect 229020 174010 229048 175102
rect 229008 174004 229060 174010
rect 229008 173946 229060 173952
rect 229112 173369 229140 177919
rect 229204 173777 229232 178706
rect 229376 178016 229428 178022
rect 229376 177958 229428 177964
rect 229284 175228 229336 175234
rect 229284 175170 229336 175176
rect 229190 173768 229246 173777
rect 229190 173703 229246 173712
rect 229192 173664 229244 173670
rect 229192 173606 229244 173612
rect 229098 173360 229154 173369
rect 229098 173295 229154 173304
rect 229100 173256 229152 173262
rect 229100 173198 229152 173204
rect 214562 163704 214618 163713
rect 214562 163639 214618 163648
rect 214932 163532 214984 163538
rect 214932 163474 214984 163480
rect 213918 163024 213974 163033
rect 213918 162959 213974 162968
rect 214012 162852 214064 162858
rect 214012 162794 214064 162800
rect 213920 162784 213972 162790
rect 213920 162726 213972 162732
rect 213932 162353 213960 162726
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162794
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161129 213960 161298
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161366
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 214012 160064 214064 160070
rect 214012 160006 214064 160012
rect 213920 159996 213972 160002
rect 213920 159938 213972 159944
rect 213932 159769 213960 159938
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 160006
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 158409 213960 158646
rect 214012 158636 214064 158642
rect 214012 158578 214064 158584
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214024 157729 214052 158578
rect 214010 157720 214066 157729
rect 214010 157655 214066 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 156505 213960 157286
rect 214944 157185 214972 163474
rect 214930 157176 214986 157185
rect 214930 157111 214986 157120
rect 213918 156496 213974 156505
rect 213918 156431 213974 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 214012 155848 214064 155854
rect 213918 155816 213974 155825
rect 214012 155790 214064 155796
rect 213918 155751 213974 155760
rect 214024 155145 214052 155790
rect 229112 155281 229140 173198
rect 229204 155825 229232 173606
rect 229296 158137 229324 175170
rect 229388 173670 229416 177958
rect 229376 173664 229428 173670
rect 229376 173606 229428 173612
rect 229480 173262 229508 178910
rect 229756 176769 229784 240071
rect 230216 235414 230244 240244
rect 230584 237862 230612 240244
rect 230572 237856 230624 237862
rect 230572 237798 230624 237804
rect 230204 235408 230256 235414
rect 230204 235350 230256 235356
rect 231136 233238 231164 240244
rect 231504 238678 231532 240244
rect 231492 238672 231544 238678
rect 231492 238614 231544 238620
rect 231768 237856 231820 237862
rect 231768 237798 231820 237804
rect 231124 233232 231176 233238
rect 231124 233174 231176 233180
rect 230756 199436 230808 199442
rect 230756 199378 230808 199384
rect 230572 188420 230624 188426
rect 230572 188362 230624 188368
rect 229742 176760 229798 176769
rect 229742 176695 229798 176704
rect 230480 175024 230532 175030
rect 230478 174992 230480 175001
rect 230532 174992 230534 175001
rect 230478 174927 230534 174936
rect 229468 173256 229520 173262
rect 229468 173198 229520 173204
rect 230480 165912 230532 165918
rect 230480 165854 230532 165860
rect 230492 165753 230520 165854
rect 230478 165744 230534 165753
rect 230478 165679 230534 165688
rect 230478 161664 230534 161673
rect 230478 161599 230534 161608
rect 229836 160812 229888 160818
rect 229836 160754 229888 160760
rect 229282 158128 229338 158137
rect 229282 158063 229338 158072
rect 229190 155816 229246 155825
rect 229190 155751 229246 155760
rect 229098 155272 229154 155281
rect 229098 155207 229154 155216
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 214010 153096 214066 153105
rect 214010 153031 214066 153040
rect 213918 152552 213974 152561
rect 213918 152487 213974 152496
rect 213932 151910 213960 152487
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 153031
rect 229744 152584 229796 152590
rect 229744 152526 229796 152532
rect 214470 151872 214526 151881
rect 214012 151836 214064 151842
rect 214470 151807 214526 151816
rect 214012 151778 214064 151784
rect 214484 151094 214512 151807
rect 215206 151192 215262 151201
rect 215206 151127 215262 151136
rect 214472 151088 214524 151094
rect 214472 151030 214524 151036
rect 213918 150512 213974 150521
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149841 213960 150282
rect 213918 149832 213974 149841
rect 213918 149767 213974 149776
rect 214024 149161 214052 150350
rect 214010 149152 214066 149161
rect 215220 149138 215248 151127
rect 215220 149110 215340 149138
rect 214010 149087 214066 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146334 213960 146503
rect 214024 146402 214052 147183
rect 214012 146396 214064 146402
rect 214012 146338 214064 146344
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 145042 213960 145143
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 214024 144974 214052 145823
rect 214012 144968 214064 144974
rect 214012 144910 214064 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 214024 143682 214052 144463
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142186 213960 143239
rect 214930 142624 214986 142633
rect 214930 142559 214986 142568
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141944 214066 141953
rect 214010 141879 214066 141888
rect 213918 141264 213974 141273
rect 213918 141199 213974 141208
rect 213932 140894 213960 141199
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141879
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 214010 140584 214066 140593
rect 214010 140519 214066 140528
rect 213918 139904 213974 139913
rect 213918 139839 213974 139848
rect 213932 139466 213960 139839
rect 214024 139534 214052 140519
rect 214012 139528 214064 139534
rect 214012 139470 214064 139476
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214010 139224 214066 139233
rect 214010 139159 214066 139168
rect 214024 138038 214052 139159
rect 214944 138718 214972 142559
rect 214932 138712 214984 138718
rect 214562 138680 214618 138689
rect 214932 138654 214984 138660
rect 214562 138615 214618 138624
rect 214012 138032 214064 138038
rect 213918 138000 213974 138009
rect 214012 137974 214064 137980
rect 213918 137935 213974 137944
rect 213932 136678 213960 137935
rect 214102 137320 214158 137329
rect 214102 137255 214158 137264
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136640 214066 136649
rect 214010 136575 214066 136584
rect 214024 135386 214052 136575
rect 214116 135930 214144 137255
rect 214104 135924 214156 135930
rect 214104 135866 214156 135872
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213918 135280 213920 135289
rect 213972 135280 213974 135289
rect 213918 135215 213974 135224
rect 213918 134600 213974 134609
rect 213918 134535 213974 134544
rect 213932 133958 213960 134535
rect 213920 133952 213972 133958
rect 213366 133920 213422 133929
rect 213920 133894 213972 133900
rect 213366 133855 213422 133864
rect 213184 93832 213236 93838
rect 213184 93774 213236 93780
rect 213276 93356 213328 93362
rect 213276 93298 213328 93304
rect 211896 75880 211948 75886
rect 211896 75822 211948 75828
rect 213288 29714 213316 93298
rect 213380 92478 213408 133855
rect 214010 133376 214066 133385
rect 214010 133311 214066 133320
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132530 213960 132631
rect 214024 132598 214052 133311
rect 214012 132592 214064 132598
rect 214012 132534 214064 132540
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 131336 213974 131345
rect 213918 131271 213974 131280
rect 213932 131170 213960 131271
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 214010 129976 214066 129985
rect 214010 129911 214066 129920
rect 214024 129878 214052 129911
rect 214012 129872 214064 129878
rect 214012 129814 214064 129820
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 214010 129296 214066 129305
rect 214010 129231 214066 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128450 213960 128687
rect 213920 128444 213972 128450
rect 213920 128386 213972 128392
rect 214024 128382 214052 129231
rect 214012 128376 214064 128382
rect 214012 128318 214064 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125730 213960 125967
rect 213920 125724 213972 125730
rect 213920 125666 213972 125672
rect 214024 125662 214052 126647
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124302 213960 124607
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 125287
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122874 213960 123383
rect 214024 122942 214052 124063
rect 214012 122936 214064 122942
rect 214012 122878 214064 122884
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121582 213960 122023
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122703
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 214024 120222 214052 121343
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214102 120048 214158 120057
rect 214102 119983 214158 119992
rect 214010 119504 214066 119513
rect 214010 119439 214066 119448
rect 213920 118856 213972 118862
rect 213918 118824 213920 118833
rect 213972 118824 213974 118833
rect 213918 118759 213974 118768
rect 214024 118726 214052 119439
rect 214116 118794 214144 119983
rect 214104 118788 214156 118794
rect 214104 118730 214156 118736
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 213918 116784 213974 116793
rect 213918 116719 213974 116728
rect 213932 116006 213960 116719
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113218 213960 113455
rect 214024 113286 214052 114135
rect 214012 113280 214064 113286
rect 214012 113222 214064 113228
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106350 213960 106791
rect 214024 106418 214052 107471
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 214024 104990 214052 106111
rect 214012 104984 214064 104990
rect 213918 104952 213974 104961
rect 214012 104926 214064 104932
rect 213918 104887 213920 104896
rect 213972 104887 213974 104896
rect 213920 104858 213972 104864
rect 213918 103592 213974 103601
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 213920 103498 213972 103504
rect 213458 102912 213514 102921
rect 213458 102847 213514 102856
rect 213368 92472 213420 92478
rect 213368 92414 213420 92420
rect 213472 78674 213500 102847
rect 214576 102785 214604 138615
rect 214654 132016 214710 132025
rect 214654 131951 214710 131960
rect 214668 106962 214696 131951
rect 215312 110430 215340 149110
rect 229756 136921 229784 152526
rect 229848 146305 229876 160754
rect 230492 158681 230520 161599
rect 230478 158672 230534 158681
rect 230478 158607 230534 158616
rect 230584 157729 230612 188362
rect 230664 180192 230716 180198
rect 230664 180134 230716 180140
rect 230676 174321 230704 180134
rect 230662 174312 230718 174321
rect 230662 174247 230718 174256
rect 230570 157720 230626 157729
rect 230570 157655 230626 157664
rect 229928 152516 229980 152522
rect 229928 152458 229980 152464
rect 229834 146296 229890 146305
rect 229834 146231 229890 146240
rect 229742 136912 229798 136921
rect 229742 136847 229798 136856
rect 216034 135960 216090 135969
rect 216034 135895 216090 135904
rect 215300 110424 215352 110430
rect 215300 110366 215352 110372
rect 214656 106956 214708 106962
rect 214656 106898 214708 106904
rect 215022 105632 215078 105641
rect 215022 105567 215078 105576
rect 214838 104272 214894 104281
rect 214838 104207 214894 104216
rect 214562 102776 214618 102785
rect 214562 102711 214618 102720
rect 213918 102232 213974 102241
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 214746 101552 214802 101561
rect 214746 101487 214802 101496
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 214024 99482 214052 100263
rect 214012 99476 214064 99482
rect 214012 99418 214064 99424
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98122 213960 98223
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 214024 98054 214052 98903
rect 214012 98048 214064 98054
rect 214012 97990 214064 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96966 213960 97543
rect 213920 96960 213972 96966
rect 213920 96902 213972 96908
rect 214010 96928 214066 96937
rect 214010 96863 214066 96872
rect 214024 96830 214052 96863
rect 214012 96824 214064 96830
rect 214012 96766 214064 96772
rect 214656 96756 214708 96762
rect 214656 96698 214708 96704
rect 214102 96384 214158 96393
rect 214102 96319 214158 96328
rect 214116 95266 214144 96319
rect 214104 95260 214156 95266
rect 214104 95202 214156 95208
rect 214562 89040 214618 89049
rect 214562 88975 214618 88984
rect 213460 78668 213512 78674
rect 213460 78610 213512 78616
rect 213276 29708 213328 29714
rect 213276 29650 213328 29656
rect 211804 24132 211856 24138
rect 211804 24074 211856 24080
rect 209044 13116 209096 13122
rect 209044 13058 209096 13064
rect 198004 6248 198056 6254
rect 198004 6190 198056 6196
rect 214576 6186 214604 88975
rect 214668 39370 214696 96698
rect 214760 86873 214788 101487
rect 214852 91089 214880 104207
rect 215036 95033 215064 105567
rect 215944 96824 215996 96830
rect 215944 96766 215996 96772
rect 215022 95024 215078 95033
rect 215022 94959 215078 94968
rect 214838 91080 214894 91089
rect 214838 91015 214894 91024
rect 214746 86864 214802 86873
rect 214746 86799 214802 86808
rect 214656 39364 214708 39370
rect 214656 39306 214708 39312
rect 215956 25566 215984 96766
rect 216048 92410 216076 135895
rect 229744 135516 229796 135522
rect 229744 135458 229796 135464
rect 216218 116104 216274 116113
rect 216218 116039 216274 116048
rect 216036 92404 216088 92410
rect 216036 92346 216088 92352
rect 216128 91860 216180 91866
rect 216128 91802 216180 91808
rect 216140 55962 216168 91802
rect 216232 88330 216260 116039
rect 229192 97300 229244 97306
rect 229192 97242 229244 97248
rect 229204 97209 229232 97242
rect 229190 97200 229246 97209
rect 229190 97135 229246 97144
rect 229098 97064 229154 97073
rect 229098 96999 229154 97008
rect 220176 95260 220228 95266
rect 220176 95202 220228 95208
rect 218704 91792 218756 91798
rect 218704 91734 218756 91740
rect 217324 89072 217376 89078
rect 217324 89014 217376 89020
rect 216220 88324 216272 88330
rect 216220 88266 216272 88272
rect 216128 55956 216180 55962
rect 216128 55898 216180 55904
rect 217336 32502 217364 89014
rect 218716 46238 218744 91734
rect 220084 90500 220136 90506
rect 220084 90442 220136 90448
rect 218704 46232 218756 46238
rect 218704 46174 218756 46180
rect 217324 32496 217376 32502
rect 217324 32438 217376 32444
rect 220096 26994 220124 90442
rect 220188 51746 220216 95202
rect 229112 95198 229140 96999
rect 229192 96892 229244 96898
rect 229192 96834 229244 96840
rect 229204 96665 229232 96834
rect 229190 96656 229246 96665
rect 229190 96591 229246 96600
rect 229100 95192 229152 95198
rect 229100 95134 229152 95140
rect 225604 94784 225656 94790
rect 225604 94726 225656 94732
rect 221556 94716 221608 94722
rect 221556 94658 221608 94664
rect 221464 87712 221516 87718
rect 221464 87654 221516 87660
rect 221476 58682 221504 87654
rect 221568 79354 221596 94658
rect 224316 94580 224368 94586
rect 224316 94522 224368 94528
rect 222844 94512 222896 94518
rect 222844 94454 222896 94460
rect 221556 79348 221608 79354
rect 221556 79290 221608 79296
rect 221464 58676 221516 58682
rect 221464 58618 221516 58624
rect 220176 51740 220228 51746
rect 220176 51682 220228 51688
rect 220084 26988 220136 26994
rect 220084 26930 220136 26936
rect 215944 25560 215996 25566
rect 215944 25502 215996 25508
rect 214564 6180 214616 6186
rect 214564 6122 214616 6128
rect 178684 3596 178736 3602
rect 178684 3538 178736 3544
rect 222856 3534 222884 94454
rect 224222 93936 224278 93945
rect 224222 93871 224278 93880
rect 222934 91760 222990 91769
rect 222934 91695 222990 91704
rect 222948 64258 222976 91695
rect 222936 64252 222988 64258
rect 222936 64194 222988 64200
rect 224236 29646 224264 93871
rect 224328 53174 224356 94522
rect 224316 53168 224368 53174
rect 224316 53110 224368 53116
rect 225616 44878 225644 94726
rect 228364 94648 228416 94654
rect 228364 94590 228416 94596
rect 226984 93152 227036 93158
rect 226984 93094 227036 93100
rect 226996 58750 227024 93094
rect 226984 58744 227036 58750
rect 226984 58686 227036 58692
rect 228376 44946 228404 94590
rect 229756 61402 229784 135458
rect 229836 122868 229888 122874
rect 229836 122810 229888 122816
rect 229848 82142 229876 122810
rect 229940 113257 229968 152458
rect 230768 149705 230796 199378
rect 231780 185745 231808 237798
rect 232056 237454 232084 240244
rect 232608 239834 232636 240244
rect 232596 239828 232648 239834
rect 232596 239770 232648 239776
rect 232976 238513 233004 240244
rect 232962 238504 233018 238513
rect 232962 238439 233018 238448
rect 233528 238406 233556 240244
rect 233516 238400 233568 238406
rect 233516 238342 233568 238348
rect 234080 238338 234108 240244
rect 234068 238332 234120 238338
rect 234068 238274 234120 238280
rect 232044 237448 232096 237454
rect 232044 237390 232096 237396
rect 233148 237448 233200 237454
rect 233148 237390 233200 237396
rect 232136 236700 232188 236706
rect 232136 236642 232188 236648
rect 231766 185736 231822 185745
rect 231766 185671 231822 185680
rect 231952 179036 232004 179042
rect 231952 178978 232004 178984
rect 231860 176112 231912 176118
rect 231860 176054 231912 176060
rect 230940 175976 230992 175982
rect 230940 175918 230992 175924
rect 230952 164801 230980 175918
rect 231766 175264 231822 175273
rect 231124 175228 231176 175234
rect 231766 175199 231822 175208
rect 231124 175170 231176 175176
rect 231136 174729 231164 175170
rect 231780 175166 231808 175199
rect 231768 175160 231820 175166
rect 231768 175102 231820 175108
rect 231122 174720 231178 174729
rect 231122 174655 231178 174664
rect 231584 173868 231636 173874
rect 231584 173810 231636 173816
rect 231596 172825 231624 173810
rect 231582 172816 231638 172825
rect 231582 172751 231638 172760
rect 231676 172508 231728 172514
rect 231676 172450 231728 172456
rect 231492 172236 231544 172242
rect 231492 172178 231544 172184
rect 231504 171465 231532 172178
rect 231688 171873 231716 172450
rect 231768 172440 231820 172446
rect 231766 172408 231768 172417
rect 231820 172408 231822 172417
rect 231766 172343 231822 172352
rect 231674 171864 231730 171873
rect 231674 171799 231730 171808
rect 231490 171456 231546 171465
rect 231490 171391 231546 171400
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231492 171012 231544 171018
rect 231492 170954 231544 170960
rect 231216 170808 231268 170814
rect 231216 170750 231268 170756
rect 231228 170513 231256 170750
rect 231214 170504 231270 170513
rect 231214 170439 231270 170448
rect 231504 169969 231532 170954
rect 231780 170921 231808 171022
rect 231766 170912 231822 170921
rect 231766 170847 231822 170856
rect 231490 169960 231546 169969
rect 231490 169895 231546 169904
rect 231124 169720 231176 169726
rect 231872 169674 231900 176054
rect 231124 169662 231176 169668
rect 231136 168609 231164 169662
rect 231688 169646 231900 169674
rect 231688 169561 231716 169646
rect 231768 169584 231820 169590
rect 231674 169552 231730 169561
rect 231768 169526 231820 169532
rect 231674 169487 231730 169496
rect 231780 169017 231808 169526
rect 231766 169008 231822 169017
rect 231766 168943 231822 168952
rect 231122 168600 231178 168609
rect 231122 168535 231178 168544
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231400 168292 231452 168298
rect 231400 168234 231452 168240
rect 231412 167657 231440 168234
rect 231676 168088 231728 168094
rect 231674 168056 231676 168065
rect 231728 168056 231730 168065
rect 231674 167991 231730 168000
rect 231398 167648 231454 167657
rect 231398 167583 231454 167592
rect 231780 167113 231808 168302
rect 231766 167104 231822 167113
rect 231766 167039 231822 167048
rect 231032 166728 231084 166734
rect 231030 166696 231032 166705
rect 231084 166696 231086 166705
rect 231030 166631 231086 166640
rect 231308 166592 231360 166598
rect 231308 166534 231360 166540
rect 231124 166320 231176 166326
rect 231124 166262 231176 166268
rect 230938 164792 230994 164801
rect 230938 164727 230994 164736
rect 231136 162897 231164 166262
rect 231320 166161 231348 166534
rect 231306 166152 231362 166161
rect 231306 166087 231362 166096
rect 231400 165572 231452 165578
rect 231400 165514 231452 165520
rect 231412 165209 231440 165514
rect 231398 165200 231454 165209
rect 231308 165164 231360 165170
rect 231398 165135 231454 165144
rect 231308 165106 231360 165112
rect 231320 164393 231348 165106
rect 231306 164384 231362 164393
rect 231306 164319 231362 164328
rect 231400 164212 231452 164218
rect 231400 164154 231452 164160
rect 231412 163849 231440 164154
rect 231398 163840 231454 163849
rect 231398 163775 231454 163784
rect 231122 162888 231178 162897
rect 231122 162823 231178 162832
rect 231400 162852 231452 162858
rect 231400 162794 231452 162800
rect 230940 162784 230992 162790
rect 230940 162726 230992 162732
rect 230952 161945 230980 162726
rect 231412 162489 231440 162794
rect 231398 162480 231454 162489
rect 231398 162415 231454 162424
rect 230938 161936 230994 161945
rect 230938 161871 230994 161880
rect 231400 161900 231452 161906
rect 231400 161842 231452 161848
rect 231412 161537 231440 161842
rect 231398 161528 231454 161537
rect 231398 161463 231454 161472
rect 230940 161424 230992 161430
rect 230940 161366 230992 161372
rect 230952 160585 230980 161366
rect 231400 161220 231452 161226
rect 231400 161162 231452 161168
rect 231412 160993 231440 161162
rect 231398 160984 231454 160993
rect 231398 160919 231454 160928
rect 230938 160576 230994 160585
rect 230938 160511 230994 160520
rect 231400 160064 231452 160070
rect 231398 160032 231400 160041
rect 231452 160032 231454 160041
rect 230940 159996 230992 160002
rect 231398 159967 231454 159976
rect 230940 159938 230992 159944
rect 230952 159089 230980 159938
rect 230938 159080 230994 159089
rect 230938 159015 230994 159024
rect 231216 158024 231268 158030
rect 231216 157966 231268 157972
rect 231124 157276 231176 157282
rect 231124 157218 231176 157224
rect 231136 156777 231164 157218
rect 231122 156768 231178 156777
rect 231122 156703 231178 156712
rect 230940 155916 230992 155922
rect 230940 155858 230992 155864
rect 230952 154873 230980 155858
rect 230938 154864 230994 154873
rect 230938 154799 230994 154808
rect 231228 151814 231256 157966
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231780 157185 231808 157286
rect 231766 157176 231822 157185
rect 231766 157111 231822 157120
rect 231768 154556 231820 154562
rect 231768 154498 231820 154504
rect 231780 154329 231808 154498
rect 231766 154320 231822 154329
rect 231766 154255 231822 154264
rect 231492 154012 231544 154018
rect 231492 153954 231544 153960
rect 231504 153377 231532 153954
rect 231674 153776 231730 153785
rect 231674 153711 231730 153720
rect 231490 153368 231546 153377
rect 231490 153303 231546 153312
rect 231400 153196 231452 153202
rect 231400 153138 231452 153144
rect 231412 152017 231440 153138
rect 231688 152969 231716 153711
rect 231768 153128 231820 153134
rect 231768 153070 231820 153076
rect 231674 152960 231730 152969
rect 231674 152895 231730 152904
rect 231780 152561 231808 153070
rect 231766 152552 231822 152561
rect 231766 152487 231822 152496
rect 231398 152008 231454 152017
rect 231398 151943 231454 151952
rect 231964 151814 231992 178978
rect 232044 176044 232096 176050
rect 232044 175986 232096 175992
rect 231044 151786 231256 151814
rect 231872 151786 231992 151814
rect 230940 150408 230992 150414
rect 230940 150350 230992 150356
rect 230848 150340 230900 150346
rect 230848 150282 230900 150288
rect 230754 149696 230810 149705
rect 230754 149631 230810 149640
rect 230860 149161 230888 150282
rect 230952 150113 230980 150350
rect 230938 150104 230994 150113
rect 230938 150039 230994 150048
rect 230846 149152 230902 149161
rect 230846 149087 230902 149096
rect 230938 145616 230994 145625
rect 230938 145551 230994 145560
rect 230952 143041 230980 145551
rect 230938 143032 230994 143041
rect 230938 142967 230994 142976
rect 231044 134065 231072 151786
rect 231216 151632 231268 151638
rect 231214 151600 231216 151609
rect 231268 151600 231270 151609
rect 231214 151535 231270 151544
rect 231216 151088 231268 151094
rect 231216 151030 231268 151036
rect 231124 148368 231176 148374
rect 231124 148310 231176 148316
rect 231136 148209 231164 148310
rect 231122 148200 231178 148209
rect 231122 148135 231178 148144
rect 231228 135969 231256 151030
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148753 231808 148990
rect 231766 148744 231822 148753
rect 231766 148679 231822 148688
rect 231400 148300 231452 148306
rect 231400 148242 231452 148248
rect 231308 144900 231360 144906
rect 231308 144842 231360 144848
rect 231320 144401 231348 144842
rect 231306 144392 231362 144401
rect 231306 144327 231362 144336
rect 231308 143404 231360 143410
rect 231308 143346 231360 143352
rect 231320 142497 231348 143346
rect 231306 142488 231362 142497
rect 231306 142423 231362 142432
rect 231308 138712 231360 138718
rect 231308 138654 231360 138660
rect 231214 135960 231270 135969
rect 231124 135924 231176 135930
rect 231214 135895 231270 135904
rect 231124 135866 231176 135872
rect 231030 134056 231086 134065
rect 231030 133991 231086 134000
rect 231136 133113 231164 135866
rect 231216 133612 231268 133618
rect 231216 133554 231268 133560
rect 231122 133104 231178 133113
rect 231122 133039 231178 133048
rect 231124 129124 231176 129130
rect 231124 129066 231176 129072
rect 230848 128308 230900 128314
rect 230848 128250 230900 128256
rect 230860 127945 230888 128250
rect 230846 127936 230902 127945
rect 230846 127871 230902 127880
rect 231032 127628 231084 127634
rect 231032 127570 231084 127576
rect 230940 124636 230992 124642
rect 230940 124578 230992 124584
rect 230756 124160 230808 124166
rect 230754 124128 230756 124137
rect 230808 124128 230810 124137
rect 230754 124063 230810 124072
rect 230756 123616 230808 123622
rect 230952 123593 230980 124578
rect 230756 123558 230808 123564
rect 230938 123584 230994 123593
rect 230768 121689 230796 123558
rect 230938 123519 230994 123528
rect 231044 122834 231072 127570
rect 231136 126041 231164 129066
rect 231122 126032 231178 126041
rect 231122 125967 231178 125976
rect 231044 122806 231164 122834
rect 230754 121680 230810 121689
rect 230754 121615 230810 121624
rect 230756 120760 230808 120766
rect 230756 120702 230808 120708
rect 230768 118969 230796 120702
rect 230940 120080 230992 120086
rect 230940 120022 230992 120028
rect 230952 119785 230980 120022
rect 230938 119776 230994 119785
rect 230938 119711 230994 119720
rect 230754 118960 230810 118969
rect 230754 118895 230810 118904
rect 230664 117020 230716 117026
rect 230664 116962 230716 116968
rect 230676 116113 230704 116962
rect 230662 116104 230718 116113
rect 230662 116039 230718 116048
rect 230020 115252 230072 115258
rect 230020 115194 230072 115200
rect 229926 113248 229982 113257
rect 229926 113183 229982 113192
rect 230032 93362 230060 115194
rect 230848 113824 230900 113830
rect 230848 113766 230900 113772
rect 230572 111716 230624 111722
rect 230572 111658 230624 111664
rect 230584 110809 230612 111658
rect 230570 110800 230626 110809
rect 230570 110735 230626 110744
rect 230572 110356 230624 110362
rect 230572 110298 230624 110304
rect 230584 109449 230612 110298
rect 230570 109440 230626 109449
rect 230570 109375 230626 109384
rect 230860 107953 230888 113766
rect 230846 107944 230902 107953
rect 230846 107879 230902 107888
rect 230572 106140 230624 106146
rect 230572 106082 230624 106088
rect 230584 105233 230612 106082
rect 230570 105224 230626 105233
rect 230570 105159 230626 105168
rect 230848 104780 230900 104786
rect 230848 104722 230900 104728
rect 230860 104281 230888 104722
rect 230846 104272 230902 104281
rect 230756 104236 230808 104242
rect 230846 104207 230902 104216
rect 230756 104178 230808 104184
rect 230768 100473 230796 104178
rect 231136 101833 231164 122806
rect 231228 116521 231256 133554
rect 231320 131209 231348 138654
rect 231412 135425 231440 148242
rect 231766 146840 231822 146849
rect 231872 146826 231900 151786
rect 232056 150657 232084 175986
rect 232148 165918 232176 236642
rect 233160 213246 233188 237390
rect 233332 233232 233384 233238
rect 233332 233174 233384 233180
rect 233148 213240 233200 213246
rect 233148 213182 233200 213188
rect 232136 165912 232188 165918
rect 232136 165854 232188 165860
rect 232504 155236 232556 155242
rect 232504 155178 232556 155184
rect 232042 150648 232098 150657
rect 232042 150583 232098 150592
rect 231822 146798 231900 146826
rect 231766 146775 231822 146784
rect 231768 146260 231820 146266
rect 231768 146202 231820 146208
rect 231780 145897 231808 146202
rect 231766 145888 231822 145897
rect 231766 145823 231822 145832
rect 231676 145444 231728 145450
rect 231676 145386 231728 145392
rect 231688 144945 231716 145386
rect 231674 144936 231730 144945
rect 231674 144871 231730 144880
rect 231492 144832 231544 144838
rect 231492 144774 231544 144780
rect 231504 143993 231532 144774
rect 231490 143984 231546 143993
rect 231490 143919 231546 143928
rect 231768 142112 231820 142118
rect 231768 142054 231820 142060
rect 231780 141137 231808 142054
rect 231766 141128 231822 141137
rect 231766 141063 231822 141072
rect 231676 140752 231728 140758
rect 231676 140694 231728 140700
rect 231766 140720 231822 140729
rect 231688 140185 231716 140694
rect 231766 140655 231768 140664
rect 231820 140655 231822 140664
rect 231768 140626 231820 140632
rect 231674 140176 231730 140185
rect 231674 140111 231730 140120
rect 231768 139392 231820 139398
rect 231768 139334 231820 139340
rect 231780 138281 231808 139334
rect 231766 138272 231822 138281
rect 231766 138207 231822 138216
rect 231676 137896 231728 137902
rect 231674 137864 231676 137873
rect 231728 137864 231730 137873
rect 231674 137799 231730 137808
rect 231398 135416 231454 135425
rect 231398 135351 231454 135360
rect 231768 135244 231820 135250
rect 231768 135186 231820 135192
rect 231676 135176 231728 135182
rect 231676 135118 231728 135124
rect 231688 134473 231716 135118
rect 231780 135017 231808 135186
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231676 133884 231728 133890
rect 231676 133826 231728 133832
rect 231688 132569 231716 133826
rect 231768 133816 231820 133822
rect 231768 133758 231820 133764
rect 231780 133521 231808 133758
rect 231766 133512 231822 133521
rect 231766 133447 231822 133456
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231676 132388 231728 132394
rect 231676 132330 231728 132336
rect 231688 131617 231716 132330
rect 231780 132161 231808 132398
rect 231766 132152 231822 132161
rect 231766 132087 231822 132096
rect 231674 131608 231730 131617
rect 231674 131543 231730 131552
rect 231306 131200 231362 131209
rect 231306 131135 231362 131144
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231676 131028 231728 131034
rect 231676 130970 231728 130976
rect 231584 130960 231636 130966
rect 231584 130902 231636 130908
rect 231596 129849 231624 130902
rect 231688 130257 231716 130970
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231674 130248 231730 130257
rect 231674 130183 231730 130192
rect 231582 129840 231638 129849
rect 231582 129775 231638 129784
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231676 129668 231728 129674
rect 231676 129610 231728 129616
rect 231584 129056 231636 129062
rect 231584 128998 231636 129004
rect 231492 125588 231544 125594
rect 231492 125530 231544 125536
rect 231504 124545 231532 125530
rect 231490 124536 231546 124545
rect 231490 124471 231546 124480
rect 231596 123185 231624 128998
rect 231688 128897 231716 129610
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231674 128888 231730 128897
rect 231674 128823 231730 128832
rect 231766 128344 231822 128353
rect 231766 128279 231822 128288
rect 231780 128246 231808 128279
rect 231768 128240 231820 128246
rect 231768 128182 231820 128188
rect 231766 126984 231822 126993
rect 231766 126919 231768 126928
rect 231820 126919 231822 126928
rect 231768 126890 231820 126896
rect 231676 126880 231728 126886
rect 231676 126822 231728 126828
rect 231688 126449 231716 126822
rect 231674 126440 231730 126449
rect 231674 126375 231730 126384
rect 231768 125520 231820 125526
rect 231766 125488 231768 125497
rect 231820 125488 231822 125497
rect 231766 125423 231822 125432
rect 231768 125112 231820 125118
rect 231766 125080 231768 125089
rect 231820 125080 231822 125089
rect 231766 125015 231822 125024
rect 232516 124166 232544 155178
rect 232780 153264 232832 153270
rect 232780 153206 232832 153212
rect 232596 146328 232648 146334
rect 232596 146270 232648 146276
rect 232504 124160 232556 124166
rect 232504 124102 232556 124108
rect 231582 123176 231638 123185
rect 231582 123111 231638 123120
rect 231676 122800 231728 122806
rect 231676 122742 231728 122748
rect 231688 122233 231716 122742
rect 231768 122732 231820 122738
rect 231768 122674 231820 122680
rect 231780 122641 231808 122674
rect 231766 122632 231822 122641
rect 231766 122567 231822 122576
rect 231674 122224 231730 122233
rect 231674 122159 231730 122168
rect 231676 122120 231728 122126
rect 231676 122062 231728 122068
rect 231584 121304 231636 121310
rect 231584 121246 231636 121252
rect 231596 120737 231624 121246
rect 231582 120728 231638 120737
rect 231582 120663 231638 120672
rect 231688 120329 231716 122062
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 121281 231808 121382
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231674 120320 231730 120329
rect 231674 120255 231730 120264
rect 232504 120148 232556 120154
rect 232504 120090 232556 120096
rect 231400 120012 231452 120018
rect 231400 119954 231452 119960
rect 231412 119377 231440 119954
rect 231398 119368 231454 119377
rect 231398 119303 231454 119312
rect 231308 118720 231360 118726
rect 231308 118662 231360 118668
rect 231214 116512 231270 116521
rect 231214 116447 231270 116456
rect 231320 111761 231348 118662
rect 231492 118652 231544 118658
rect 231492 118594 231544 118600
rect 231504 117473 231532 118594
rect 231768 118584 231820 118590
rect 231768 118526 231820 118532
rect 231676 118448 231728 118454
rect 231674 118416 231676 118425
rect 231728 118416 231730 118425
rect 231674 118351 231730 118360
rect 231780 118017 231808 118526
rect 231766 118008 231822 118017
rect 231766 117943 231822 117952
rect 231490 117464 231546 117473
rect 231490 117399 231546 117408
rect 231768 117292 231820 117298
rect 231768 117234 231820 117240
rect 231780 117065 231808 117234
rect 231766 117056 231822 117065
rect 231766 116991 231822 117000
rect 231768 115932 231820 115938
rect 231768 115874 231820 115880
rect 231676 115864 231728 115870
rect 231676 115806 231728 115812
rect 231688 114617 231716 115806
rect 231780 115569 231808 115874
rect 231766 115560 231822 115569
rect 231766 115495 231822 115504
rect 231768 115320 231820 115326
rect 231768 115262 231820 115268
rect 231674 114608 231730 114617
rect 231674 114543 231730 114552
rect 231492 114504 231544 114510
rect 231492 114446 231544 114452
rect 231504 113665 231532 114446
rect 231780 114209 231808 115262
rect 231766 114200 231822 114209
rect 231766 114135 231822 114144
rect 231490 113656 231546 113665
rect 231490 113591 231546 113600
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231676 113076 231728 113082
rect 231676 113018 231728 113024
rect 231688 112305 231716 113018
rect 231780 112713 231808 113086
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 231674 112296 231730 112305
rect 231674 112231 231730 112240
rect 231768 111784 231820 111790
rect 231306 111752 231362 111761
rect 231768 111726 231820 111732
rect 231306 111687 231362 111696
rect 231780 111353 231808 111726
rect 231766 111344 231822 111353
rect 231766 111279 231822 111288
rect 231308 111104 231360 111110
rect 231308 111046 231360 111052
rect 231320 107137 231348 111046
rect 231676 110424 231728 110430
rect 231676 110366 231728 110372
rect 231766 110392 231822 110401
rect 231688 109857 231716 110366
rect 231766 110327 231822 110336
rect 231780 110294 231808 110327
rect 231768 110288 231820 110294
rect 231768 110230 231820 110236
rect 231674 109848 231730 109857
rect 231674 109783 231730 109792
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231780 108905 231808 108938
rect 231766 108896 231822 108905
rect 231766 108831 231822 108840
rect 231492 108656 231544 108662
rect 231492 108598 231544 108604
rect 231504 108497 231532 108598
rect 231490 108488 231546 108497
rect 231490 108423 231546 108432
rect 231400 108316 231452 108322
rect 231400 108258 231452 108264
rect 231306 107128 231362 107137
rect 231306 107063 231362 107072
rect 231216 106956 231268 106962
rect 231216 106898 231268 106904
rect 231122 101824 231178 101833
rect 231122 101759 231178 101768
rect 231124 100632 231176 100638
rect 231124 100574 231176 100580
rect 230754 100464 230810 100473
rect 230754 100399 230810 100408
rect 230664 100020 230716 100026
rect 230664 99962 230716 99968
rect 230676 98569 230704 99962
rect 231136 99929 231164 100574
rect 231122 99920 231178 99929
rect 231122 99855 231178 99864
rect 231124 99340 231176 99346
rect 231124 99282 231176 99288
rect 230662 98560 230718 98569
rect 230662 98495 230718 98504
rect 231136 98025 231164 99282
rect 231228 98977 231256 106898
rect 231412 103514 231440 108258
rect 231492 107636 231544 107642
rect 231492 107578 231544 107584
rect 231504 106593 231532 107578
rect 231768 107568 231820 107574
rect 231766 107536 231768 107545
rect 231820 107536 231822 107545
rect 231766 107471 231822 107480
rect 231490 106584 231546 106593
rect 231490 106519 231546 106528
rect 231676 106276 231728 106282
rect 231676 106218 231728 106224
rect 231688 105641 231716 106218
rect 231768 106208 231820 106214
rect 231766 106176 231768 106185
rect 231820 106176 231822 106185
rect 231766 106111 231822 106120
rect 231674 105632 231730 105641
rect 231674 105567 231730 105576
rect 231768 104712 231820 104718
rect 231766 104680 231768 104689
rect 231820 104680 231822 104689
rect 231766 104615 231822 104624
rect 231492 103896 231544 103902
rect 231492 103838 231544 103844
rect 231504 103737 231532 103838
rect 231490 103728 231546 103737
rect 231490 103663 231546 103672
rect 231320 103486 231440 103514
rect 231768 103488 231820 103494
rect 231320 100881 231348 103486
rect 231768 103430 231820 103436
rect 231676 103420 231728 103426
rect 231676 103362 231728 103368
rect 231584 103352 231636 103358
rect 231584 103294 231636 103300
rect 231596 102377 231624 103294
rect 231688 102785 231716 103362
rect 231780 103329 231808 103430
rect 231766 103320 231822 103329
rect 231766 103255 231822 103264
rect 231674 102776 231730 102785
rect 231674 102711 231730 102720
rect 231582 102368 231638 102377
rect 231582 102303 231638 102312
rect 231768 102128 231820 102134
rect 231768 102070 231820 102076
rect 231676 101448 231728 101454
rect 231780 101425 231808 102070
rect 231676 101390 231728 101396
rect 231766 101416 231822 101425
rect 231306 100872 231362 100881
rect 231306 100807 231362 100816
rect 231584 100700 231636 100706
rect 231584 100642 231636 100648
rect 231596 99521 231624 100642
rect 231582 99512 231638 99521
rect 231582 99447 231638 99456
rect 231214 98968 231270 98977
rect 231214 98903 231270 98912
rect 231216 98048 231268 98054
rect 231122 98016 231178 98025
rect 231216 97990 231268 97996
rect 231122 97951 231178 97960
rect 231122 96248 231178 96257
rect 231122 96183 231178 96192
rect 231136 95878 231164 96183
rect 231124 95872 231176 95878
rect 231124 95814 231176 95820
rect 230664 95192 230716 95198
rect 230664 95134 230716 95140
rect 230676 93770 230704 95134
rect 231228 93854 231256 97990
rect 231688 97617 231716 101390
rect 231766 101351 231822 101360
rect 231674 97608 231730 97617
rect 231674 97543 231730 97552
rect 231136 93826 231256 93854
rect 230664 93764 230716 93770
rect 230664 93706 230716 93712
rect 230020 93356 230072 93362
rect 230020 93298 230072 93304
rect 230676 92614 230704 93706
rect 230664 92608 230716 92614
rect 230664 92550 230716 92556
rect 229836 82136 229888 82142
rect 229836 82078 229888 82084
rect 229744 61396 229796 61402
rect 229744 61338 229796 61344
rect 231136 49026 231164 93826
rect 231216 92608 231268 92614
rect 231216 92550 231268 92556
rect 231124 49020 231176 49026
rect 231124 48962 231176 48968
rect 231228 47666 231256 92550
rect 231216 47660 231268 47666
rect 231216 47602 231268 47608
rect 228364 44940 228416 44946
rect 228364 44882 228416 44888
rect 225604 44872 225656 44878
rect 225604 44814 225656 44820
rect 224224 29640 224276 29646
rect 224224 29582 224276 29588
rect 232516 4894 232544 120090
rect 232608 104786 232636 146270
rect 232688 122936 232740 122942
rect 232688 122878 232740 122884
rect 232596 104780 232648 104786
rect 232596 104722 232648 104728
rect 232700 89146 232728 122878
rect 232792 118726 232820 153206
rect 233344 151638 233372 233174
rect 233884 201884 233936 201890
rect 233884 201826 233936 201832
rect 233422 177440 233478 177449
rect 233422 177375 233478 177384
rect 233436 169726 233464 177375
rect 233424 169720 233476 169726
rect 233424 169662 233476 169668
rect 233896 166734 233924 201826
rect 233884 166728 233936 166734
rect 233884 166670 233936 166676
rect 234448 161430 234476 240244
rect 235000 239970 235028 240244
rect 234988 239964 235040 239970
rect 234988 239906 235040 239912
rect 234528 238332 234580 238338
rect 234528 238274 234580 238280
rect 234540 181558 234568 238274
rect 235264 236836 235316 236842
rect 235264 236778 235316 236784
rect 234618 236056 234674 236065
rect 234618 235991 234674 236000
rect 234528 181552 234580 181558
rect 234528 181494 234580 181500
rect 234436 161424 234488 161430
rect 234436 161366 234488 161372
rect 234160 160744 234212 160750
rect 234160 160686 234212 160692
rect 234068 155984 234120 155990
rect 234068 155926 234120 155932
rect 233332 151632 233384 151638
rect 233332 151574 233384 151580
rect 233884 140820 233936 140826
rect 233884 140762 233936 140768
rect 232780 118720 232832 118726
rect 232780 118662 232832 118668
rect 233896 99346 233924 140762
rect 233976 136672 234028 136678
rect 233976 136614 234028 136620
rect 233884 99340 233936 99346
rect 233884 99282 233936 99288
rect 233884 95872 233936 95878
rect 233884 95814 233936 95820
rect 232688 89140 232740 89146
rect 232688 89082 232740 89088
rect 232504 4888 232556 4894
rect 232504 4830 232556 4836
rect 222844 3528 222896 3534
rect 222844 3470 222896 3476
rect 177304 3460 177356 3466
rect 177304 3402 177356 3408
rect 233896 3058 233924 95814
rect 233988 69834 234016 136614
rect 234080 117026 234108 155926
rect 234172 121310 234200 160686
rect 234252 149796 234304 149802
rect 234252 149738 234304 149744
rect 234264 137902 234292 149738
rect 234632 148374 234660 235991
rect 234804 177472 234856 177478
rect 234804 177414 234856 177420
rect 234710 175944 234766 175953
rect 234710 175879 234766 175888
rect 234724 155922 234752 175879
rect 234816 168094 234844 177414
rect 235276 172242 235304 236778
rect 235368 236706 235396 240244
rect 235920 240106 235948 240244
rect 235908 240100 235960 240106
rect 235908 240042 235960 240048
rect 236472 238678 236500 240244
rect 236460 238672 236512 238678
rect 236460 238614 236512 238620
rect 236840 237454 236868 240244
rect 237392 237454 237420 240244
rect 236828 237448 236880 237454
rect 236828 237390 236880 237396
rect 237288 237448 237340 237454
rect 237288 237390 237340 237396
rect 237380 237448 237432 237454
rect 237380 237390 237432 237396
rect 235356 236700 235408 236706
rect 235356 236642 235408 236648
rect 236000 184476 236052 184482
rect 236000 184418 236052 184424
rect 235264 172236 235316 172242
rect 235264 172178 235316 172184
rect 234804 168088 234856 168094
rect 234804 168030 234856 168036
rect 235540 163124 235592 163130
rect 235540 163066 235592 163072
rect 234712 155916 234764 155922
rect 234712 155858 234764 155864
rect 235448 149116 235500 149122
rect 235448 149058 235500 149064
rect 234620 148368 234672 148374
rect 234620 148310 234672 148316
rect 235356 144968 235408 144974
rect 235356 144910 235408 144916
rect 234252 137896 234304 137902
rect 234252 137838 234304 137844
rect 235264 124228 235316 124234
rect 235264 124170 235316 124176
rect 234160 121304 234212 121310
rect 234160 121246 234212 121252
rect 234068 117020 234120 117026
rect 234068 116962 234120 116968
rect 234160 116612 234212 116618
rect 234160 116554 234212 116560
rect 234066 114472 234122 114481
rect 234066 114407 234122 114416
rect 234080 96898 234108 114407
rect 234068 96892 234120 96898
rect 234068 96834 234120 96840
rect 234080 93702 234108 96834
rect 234172 94790 234200 116554
rect 234160 94784 234212 94790
rect 234160 94726 234212 94732
rect 234068 93696 234120 93702
rect 234068 93638 234120 93644
rect 233976 69828 234028 69834
rect 233976 69770 234028 69776
rect 235276 68406 235304 124170
rect 235368 103902 235396 144910
rect 235460 108662 235488 149058
rect 235552 124642 235580 163066
rect 236012 145450 236040 184418
rect 237300 180198 237328 237390
rect 237944 201890 237972 240244
rect 238312 237425 238340 240244
rect 238864 240038 238892 240244
rect 238852 240032 238904 240038
rect 238852 239974 238904 239980
rect 239232 238746 239260 240244
rect 239784 240145 239812 240244
rect 239770 240136 239826 240145
rect 239770 240071 239826 240080
rect 239220 238740 239272 238746
rect 239220 238682 239272 238688
rect 238760 238060 238812 238066
rect 238760 238002 238812 238008
rect 238668 237448 238720 237454
rect 238298 237416 238354 237425
rect 238668 237390 238720 237396
rect 238298 237351 238354 237360
rect 237932 201884 237984 201890
rect 237932 201826 237984 201832
rect 237564 180260 237616 180266
rect 237564 180202 237616 180208
rect 237288 180192 237340 180198
rect 237288 180134 237340 180140
rect 237472 178900 237524 178906
rect 237472 178842 237524 178848
rect 236092 178832 236144 178838
rect 236092 178774 236144 178780
rect 236104 170814 236132 178774
rect 236184 178696 236236 178702
rect 236184 178638 236236 178644
rect 236092 170808 236144 170814
rect 236092 170750 236144 170756
rect 236196 166598 236224 178638
rect 236276 173936 236328 173942
rect 236276 173878 236328 173884
rect 236184 166592 236236 166598
rect 236184 166534 236236 166540
rect 236288 161226 236316 173878
rect 236828 164280 236880 164286
rect 236828 164222 236880 164228
rect 236276 161220 236328 161226
rect 236276 161162 236328 161168
rect 236736 158772 236788 158778
rect 236736 158714 236788 158720
rect 236000 145444 236052 145450
rect 236000 145386 236052 145392
rect 236644 136740 236696 136746
rect 236644 136682 236696 136688
rect 235540 124636 235592 124642
rect 235540 124578 235592 124584
rect 235448 108656 235500 108662
rect 235448 108598 235500 108604
rect 235448 104168 235500 104174
rect 235448 104110 235500 104116
rect 235356 103896 235408 103902
rect 235356 103838 235408 103844
rect 235460 92002 235488 104110
rect 235448 91996 235500 92002
rect 235448 91938 235500 91944
rect 235264 68400 235316 68406
rect 235264 68342 235316 68348
rect 236656 36582 236684 136682
rect 236748 118454 236776 158714
rect 236840 125118 236868 164222
rect 237484 161906 237512 178842
rect 237576 165170 237604 180202
rect 238680 178702 238708 237390
rect 238668 178696 238720 178702
rect 238668 178638 238720 178644
rect 237656 174548 237708 174554
rect 237656 174490 237708 174496
rect 237564 165164 237616 165170
rect 237564 165106 237616 165112
rect 237472 161900 237524 161906
rect 237472 161842 237524 161848
rect 237668 154018 237696 174490
rect 238772 169590 238800 238002
rect 240336 237454 240364 240244
rect 240508 240168 240560 240174
rect 240600 240168 240652 240174
rect 240508 240110 240560 240116
rect 240598 240136 240600 240145
rect 240652 240136 240654 240145
rect 240324 237448 240376 237454
rect 240324 237390 240376 237396
rect 240520 236162 240548 240110
rect 240704 240122 240732 240244
rect 240968 240168 241020 240174
rect 240704 240116 240968 240122
rect 240704 240110 241020 240116
rect 240704 240094 241008 240110
rect 241152 240100 241204 240106
rect 240598 240071 240654 240080
rect 241152 240042 241204 240048
rect 241164 239986 241192 240042
rect 240980 239970 241192 239986
rect 240968 239964 241192 239970
rect 241020 239958 241192 239964
rect 240968 239906 241020 239912
rect 240508 236156 240560 236162
rect 240508 236098 240560 236104
rect 240968 236156 241020 236162
rect 240968 236098 241020 236104
rect 239404 233572 239456 233578
rect 239404 233514 239456 233520
rect 238850 183016 238906 183025
rect 238850 182951 238906 182960
rect 238760 169584 238812 169590
rect 238760 169526 238812 169532
rect 238864 164218 238892 182951
rect 238852 164212 238904 164218
rect 238852 164154 238904 164160
rect 238024 161492 238076 161498
rect 238024 161434 238076 161440
rect 237656 154012 237708 154018
rect 237656 153954 237708 153960
rect 237380 144220 237432 144226
rect 237380 144162 237432 144168
rect 237392 143410 237420 144162
rect 237380 143404 237432 143410
rect 237380 143346 237432 143352
rect 236920 125656 236972 125662
rect 236920 125598 236972 125604
rect 236828 125112 236880 125118
rect 236828 125054 236880 125060
rect 236736 118448 236788 118454
rect 236736 118390 236788 118396
rect 236736 110492 236788 110498
rect 236736 110434 236788 110440
rect 236748 72622 236776 110434
rect 236932 93294 236960 125598
rect 238036 123622 238064 161434
rect 238300 157412 238352 157418
rect 238300 157354 238352 157360
rect 238208 142180 238260 142186
rect 238208 142122 238260 142128
rect 238116 133952 238168 133958
rect 238116 133894 238168 133900
rect 238024 123616 238076 123622
rect 238024 123558 238076 123564
rect 238024 109064 238076 109070
rect 238024 109006 238076 109012
rect 236920 93288 236972 93294
rect 236920 93230 236972 93236
rect 236736 72616 236788 72622
rect 236736 72558 236788 72564
rect 236644 36576 236696 36582
rect 236644 36518 236696 36524
rect 238036 8974 238064 109006
rect 238128 35290 238156 133894
rect 238220 100638 238248 142122
rect 238312 133618 238340 157354
rect 239416 144838 239444 233514
rect 240980 219434 241008 236098
rect 241256 234614 241284 240244
rect 241428 237448 241480 237454
rect 241428 237390 241480 237396
rect 241256 234586 241376 234614
rect 241348 228478 241376 234586
rect 241336 228472 241388 228478
rect 241336 228414 241388 228420
rect 240796 219406 241008 219434
rect 240416 189984 240468 189990
rect 240416 189926 240468 189932
rect 240428 184414 240456 189926
rect 240140 184408 240192 184414
rect 240140 184350 240192 184356
rect 240416 184408 240468 184414
rect 240416 184350 240468 184356
rect 239496 169788 239548 169794
rect 239496 169730 239548 169736
rect 239404 144832 239456 144838
rect 239404 144774 239456 144780
rect 239508 138718 239536 169730
rect 240152 160818 240180 184350
rect 240230 178664 240286 178673
rect 240230 178599 240286 178608
rect 240244 171018 240272 178599
rect 240232 171012 240284 171018
rect 240232 170954 240284 170960
rect 240140 160812 240192 160818
rect 240140 160754 240192 160760
rect 239680 154624 239732 154630
rect 239680 154566 239732 154572
rect 239588 143608 239640 143614
rect 239588 143550 239640 143556
rect 239496 138712 239548 138718
rect 239496 138654 239548 138660
rect 239404 138032 239456 138038
rect 239404 137974 239456 137980
rect 238300 133612 238352 133618
rect 238300 133554 238352 133560
rect 238300 120216 238352 120222
rect 238300 120158 238352 120164
rect 238208 100632 238260 100638
rect 238208 100574 238260 100580
rect 238312 93226 238340 120158
rect 238300 93220 238352 93226
rect 238300 93162 238352 93168
rect 239416 69766 239444 137974
rect 239496 134020 239548 134026
rect 239496 133962 239548 133968
rect 239508 73982 239536 133962
rect 239600 127634 239628 143550
rect 239588 127628 239640 127634
rect 239588 127570 239640 127576
rect 239588 124296 239640 124302
rect 239588 124238 239640 124244
rect 239600 80782 239628 124238
rect 239692 115326 239720 154566
rect 240796 150346 240824 219406
rect 241440 178770 241468 237390
rect 241612 181688 241664 181694
rect 241612 181630 241664 181636
rect 241428 178764 241480 178770
rect 241428 178706 241480 178712
rect 241520 176588 241572 176594
rect 241520 176530 241572 176536
rect 241532 176497 241560 176530
rect 241518 176488 241574 176497
rect 241518 176423 241574 176432
rect 240968 172712 241020 172718
rect 240968 172654 241020 172660
rect 240876 160132 240928 160138
rect 240876 160074 240928 160080
rect 240784 150340 240836 150346
rect 240784 150282 240836 150288
rect 240784 136808 240836 136814
rect 240784 136750 240836 136756
rect 239680 115320 239732 115326
rect 239680 115262 239732 115268
rect 239588 80776 239640 80782
rect 239588 80718 239640 80724
rect 239496 73976 239548 73982
rect 239496 73918 239548 73924
rect 239404 69760 239456 69766
rect 239404 69702 239456 69708
rect 240796 38010 240824 136750
rect 240888 120018 240916 160074
rect 240980 158030 241008 172654
rect 241152 167068 241204 167074
rect 241152 167010 241204 167016
rect 240968 158024 241020 158030
rect 240968 157966 241020 157972
rect 241060 142248 241112 142254
rect 241060 142190 241112 142196
rect 240968 140888 241020 140894
rect 240968 140830 241020 140836
rect 240876 120012 240928 120018
rect 240876 119954 240928 119960
rect 240876 102400 240928 102406
rect 240876 102342 240928 102348
rect 240784 38004 240836 38010
rect 240784 37946 240836 37952
rect 238116 35284 238168 35290
rect 238116 35226 238168 35232
rect 238024 8968 238076 8974
rect 238024 8910 238076 8916
rect 240888 7682 240916 102342
rect 240980 100026 241008 140830
rect 241072 108322 241100 142190
rect 241164 141409 241192 167010
rect 241624 162790 241652 181630
rect 241612 162784 241664 162790
rect 241612 162726 241664 162732
rect 241244 156052 241296 156058
rect 241244 155994 241296 156000
rect 241150 141400 241206 141409
rect 241150 141335 241206 141344
rect 241256 137329 241284 155994
rect 241808 144226 241836 240244
rect 242176 233578 242204 240244
rect 242728 239902 242756 240244
rect 242716 239896 242768 239902
rect 242716 239838 242768 239844
rect 243280 236842 243308 240244
rect 243268 236836 243320 236842
rect 243268 236778 243320 236784
rect 243648 234122 243676 240244
rect 244108 238746 244136 241470
rect 244096 238740 244148 238746
rect 244096 238682 244148 238688
rect 244200 234705 244228 244151
rect 244186 234696 244242 234705
rect 244186 234631 244242 234640
rect 243636 234116 243688 234122
rect 243636 234058 243688 234064
rect 242164 233572 242216 233578
rect 242164 233514 242216 233520
rect 242900 192568 242952 192574
rect 242900 192510 242952 192516
rect 242440 165640 242492 165646
rect 242440 165582 242492 165588
rect 242348 162988 242400 162994
rect 242348 162930 242400 162936
rect 242164 145036 242216 145042
rect 242164 144978 242216 144984
rect 241796 144220 241848 144226
rect 241796 144162 241848 144168
rect 241242 137320 241298 137329
rect 241242 137255 241298 137264
rect 241060 108316 241112 108322
rect 241060 108258 241112 108264
rect 241152 107908 241204 107914
rect 241152 107850 241204 107856
rect 240968 100020 241020 100026
rect 240968 99962 241020 99968
rect 241164 75274 241192 107850
rect 242176 103426 242204 144978
rect 242256 143676 242308 143682
rect 242256 143618 242308 143624
rect 242164 103420 242216 103426
rect 242164 103362 242216 103368
rect 242268 103358 242296 143618
rect 242360 122738 242388 162930
rect 242452 129130 242480 165582
rect 242912 140690 242940 192510
rect 242992 184544 243044 184550
rect 242992 184486 243044 184492
rect 243004 154562 243032 184486
rect 243728 160200 243780 160206
rect 243728 160142 243780 160148
rect 242992 154556 243044 154562
rect 242992 154498 243044 154504
rect 242900 140684 242952 140690
rect 242900 140626 242952 140632
rect 243544 139460 243596 139466
rect 243544 139402 243596 139408
rect 242440 129124 242492 129130
rect 242440 129066 242492 129072
rect 242348 122732 242400 122738
rect 242348 122674 242400 122680
rect 242532 120284 242584 120290
rect 242532 120226 242584 120232
rect 242348 106480 242400 106486
rect 242348 106422 242400 106428
rect 242256 103352 242308 103358
rect 242256 103294 242308 103300
rect 242164 99408 242216 99414
rect 242164 99350 242216 99356
rect 241152 75268 241204 75274
rect 241152 75210 241204 75216
rect 240876 7676 240928 7682
rect 240876 7618 240928 7624
rect 242176 7614 242204 99350
rect 242360 66910 242388 106422
rect 242440 102264 242492 102270
rect 242440 102206 242492 102212
rect 242452 73914 242480 102206
rect 242544 91934 242572 120226
rect 242532 91928 242584 91934
rect 242532 91870 242584 91876
rect 243556 76702 243584 139402
rect 243740 122126 243768 160142
rect 244292 144906 244320 260879
rect 244936 260778 244964 474710
rect 246304 356720 246356 356726
rect 246304 356662 246356 356668
rect 245660 291916 245712 291922
rect 245660 291858 245712 291864
rect 245672 283801 245700 291858
rect 245750 290592 245806 290601
rect 245750 290527 245806 290536
rect 245658 283792 245714 283801
rect 245658 283727 245714 283736
rect 245764 263945 245792 290527
rect 245844 289128 245896 289134
rect 245844 289070 245896 289076
rect 245856 267594 245884 289070
rect 246028 282872 246080 282878
rect 246028 282814 246080 282820
rect 245934 282432 245990 282441
rect 245934 282367 245990 282376
rect 245948 281586 245976 282367
rect 246040 281625 246068 282814
rect 246026 281616 246082 281625
rect 245936 281580 245988 281586
rect 246026 281551 246082 281560
rect 245936 281522 245988 281528
rect 246026 281072 246082 281081
rect 246026 281007 246082 281016
rect 246040 280294 246068 281007
rect 246028 280288 246080 280294
rect 245934 280256 245990 280265
rect 246028 280230 246080 280236
rect 245934 280191 245936 280200
rect 245988 280191 245990 280200
rect 245936 280162 245988 280168
rect 245934 279440 245990 279449
rect 245934 279375 245990 279384
rect 245948 278798 245976 279375
rect 245936 278792 245988 278798
rect 245936 278734 245988 278740
rect 245936 278180 245988 278186
rect 245936 278122 245988 278128
rect 245948 278089 245976 278122
rect 245934 278080 245990 278089
rect 245934 278015 245990 278024
rect 245934 277536 245990 277545
rect 245934 277471 245990 277480
rect 245948 277438 245976 277471
rect 245936 277432 245988 277438
rect 245936 277374 245988 277380
rect 246026 276720 246082 276729
rect 246026 276655 246082 276664
rect 246040 276078 246068 276655
rect 246028 276072 246080 276078
rect 246028 276014 246080 276020
rect 245936 276004 245988 276010
rect 245936 275946 245988 275952
rect 245948 275913 245976 275946
rect 245934 275904 245990 275913
rect 245934 275839 245990 275848
rect 245936 275392 245988 275398
rect 245934 275360 245936 275369
rect 245988 275360 245990 275369
rect 245934 275295 245990 275304
rect 246026 274544 246082 274553
rect 246026 274479 246082 274488
rect 245934 273728 245990 273737
rect 245934 273663 245990 273672
rect 245948 273358 245976 273663
rect 245936 273352 245988 273358
rect 245936 273294 245988 273300
rect 246040 273290 246068 274479
rect 246028 273284 246080 273290
rect 246028 273226 246080 273232
rect 246026 273184 246082 273193
rect 246026 273119 246082 273128
rect 245934 272368 245990 272377
rect 245934 272303 245990 272312
rect 245948 271930 245976 272303
rect 246040 271998 246068 273119
rect 246028 271992 246080 271998
rect 246028 271934 246080 271940
rect 245936 271924 245988 271930
rect 245936 271866 245988 271872
rect 246026 271552 246082 271561
rect 246026 271487 246082 271496
rect 245934 271008 245990 271017
rect 245934 270943 245990 270952
rect 245948 270570 245976 270943
rect 246040 270638 246068 271487
rect 246028 270632 246080 270638
rect 246028 270574 246080 270580
rect 245936 270564 245988 270570
rect 245936 270506 245988 270512
rect 245934 269648 245990 269657
rect 245934 269583 245990 269592
rect 245948 269142 245976 269583
rect 245936 269136 245988 269142
rect 245936 269078 245988 269084
rect 246026 268832 246082 268841
rect 246026 268767 246082 268776
rect 245934 268016 245990 268025
rect 245934 267951 245990 267960
rect 245948 267782 245976 267951
rect 246040 267850 246068 268767
rect 246028 267844 246080 267850
rect 246028 267786 246080 267792
rect 245936 267776 245988 267782
rect 245936 267718 245988 267724
rect 245856 267566 246160 267594
rect 246026 267472 246082 267481
rect 246026 267407 246082 267416
rect 246040 266422 246068 267407
rect 246028 266416 246080 266422
rect 246028 266358 246080 266364
rect 245936 266348 245988 266354
rect 245936 266290 245988 266296
rect 245842 265840 245898 265849
rect 245842 265775 245898 265784
rect 245856 264994 245884 265775
rect 245948 265305 245976 266290
rect 245934 265296 245990 265305
rect 245934 265231 245990 265240
rect 245844 264988 245896 264994
rect 245844 264930 245896 264936
rect 245934 264480 245990 264489
rect 245934 264415 245990 264424
rect 245750 263936 245806 263945
rect 245750 263871 245806 263880
rect 245948 263634 245976 264415
rect 245936 263628 245988 263634
rect 245936 263570 245988 263576
rect 245658 263120 245714 263129
rect 245658 263055 245714 263064
rect 244924 260772 244976 260778
rect 244924 260714 244976 260720
rect 244370 250880 244426 250889
rect 244370 250815 244426 250824
rect 244384 157282 244412 250815
rect 245672 229906 245700 263055
rect 245934 262304 245990 262313
rect 245934 262239 245936 262248
rect 245988 262239 245990 262248
rect 245936 262210 245988 262216
rect 245842 261760 245898 261769
rect 245842 261695 245898 261704
rect 245856 260914 245884 261695
rect 245844 260908 245896 260914
rect 245844 260850 245896 260856
rect 245844 260772 245896 260778
rect 245844 260714 245896 260720
rect 245752 256692 245804 256698
rect 245752 256634 245804 256640
rect 245764 256057 245792 256634
rect 245750 256048 245806 256057
rect 245750 255983 245806 255992
rect 245856 254425 245884 260714
rect 246132 260137 246160 267566
rect 246118 260128 246174 260137
rect 246118 260063 246174 260072
rect 245934 259584 245990 259593
rect 245934 259519 245990 259528
rect 245948 259486 245976 259519
rect 245936 259480 245988 259486
rect 245936 259422 245988 259428
rect 246026 258768 246082 258777
rect 246026 258703 246082 258712
rect 245934 258224 245990 258233
rect 246040 258194 246068 258703
rect 245934 258159 245990 258168
rect 246028 258188 246080 258194
rect 245948 258126 245976 258159
rect 246028 258130 246080 258136
rect 245936 258120 245988 258126
rect 245936 258062 245988 258068
rect 245934 257408 245990 257417
rect 245934 257343 245990 257352
rect 245948 256766 245976 257343
rect 245936 256760 245988 256766
rect 245936 256702 245988 256708
rect 245934 255232 245990 255241
rect 245934 255167 245990 255176
rect 245842 254416 245898 254425
rect 245842 254351 245898 254360
rect 245948 253978 245976 255167
rect 245936 253972 245988 253978
rect 245936 253914 245988 253920
rect 245934 253872 245990 253881
rect 245934 253807 245990 253816
rect 245842 253056 245898 253065
rect 245842 252991 245898 253000
rect 245856 252618 245884 252991
rect 245948 252686 245976 253807
rect 245936 252680 245988 252686
rect 245936 252622 245988 252628
rect 245844 252612 245896 252618
rect 245844 252554 245896 252560
rect 245936 252544 245988 252550
rect 245936 252486 245988 252492
rect 245948 252249 245976 252486
rect 245934 252240 245990 252249
rect 245934 252175 245990 252184
rect 245934 251696 245990 251705
rect 245934 251631 245990 251640
rect 245948 251258 245976 251631
rect 245936 251252 245988 251258
rect 245936 251194 245988 251200
rect 245842 250336 245898 250345
rect 245842 250271 245898 250280
rect 245856 249830 245884 250271
rect 245844 249824 245896 249830
rect 245844 249766 245896 249772
rect 245936 249756 245988 249762
rect 245936 249698 245988 249704
rect 245948 249529 245976 249698
rect 245934 249520 245990 249529
rect 245934 249455 245990 249464
rect 245844 248396 245896 248402
rect 245844 248338 245896 248344
rect 245856 248169 245884 248338
rect 245936 248328 245988 248334
rect 245936 248270 245988 248276
rect 245842 248160 245898 248169
rect 245842 248095 245898 248104
rect 245948 247353 245976 248270
rect 245934 247344 245990 247353
rect 245934 247279 245990 247288
rect 245934 245984 245990 245993
rect 245934 245919 245990 245928
rect 245948 245682 245976 245919
rect 245936 245676 245988 245682
rect 245936 245618 245988 245624
rect 246026 245168 246082 245177
rect 246026 245103 246082 245112
rect 245934 244624 245990 244633
rect 245934 244559 245990 244568
rect 245948 244322 245976 244559
rect 245936 244316 245988 244322
rect 245936 244258 245988 244264
rect 245842 243808 245898 243817
rect 245842 243743 245898 243752
rect 245856 242962 245884 243743
rect 245844 242956 245896 242962
rect 245844 242898 245896 242904
rect 245842 242448 245898 242457
rect 245842 242383 245898 242392
rect 245750 241632 245806 241641
rect 245856 241602 245884 242383
rect 245750 241567 245806 241576
rect 245844 241596 245896 241602
rect 245764 233986 245792 241567
rect 245844 241538 245896 241544
rect 245934 240816 245990 240825
rect 245934 240751 245990 240760
rect 245948 240378 245976 240751
rect 246040 240446 246068 245103
rect 246316 243001 246344 356662
rect 247040 291304 247092 291310
rect 247040 291246 247092 291252
rect 246394 266656 246450 266665
rect 246394 266591 246450 266600
rect 246408 257378 246436 266591
rect 246396 257372 246448 257378
rect 246396 257314 246448 257320
rect 246394 256592 246450 256601
rect 246394 256527 246450 256536
rect 246302 242992 246358 243001
rect 246302 242927 246358 242936
rect 246028 240440 246080 240446
rect 246028 240382 246080 240388
rect 245936 240372 245988 240378
rect 245936 240314 245988 240320
rect 245752 233980 245804 233986
rect 245752 233922 245804 233928
rect 245660 229900 245712 229906
rect 245660 229842 245712 229848
rect 245660 195356 245712 195362
rect 245660 195298 245712 195304
rect 244464 187128 244516 187134
rect 244464 187070 244516 187076
rect 244372 157276 244424 157282
rect 244372 157218 244424 157224
rect 244476 149054 244504 187070
rect 244924 168428 244976 168434
rect 244924 168370 244976 168376
rect 244464 149048 244516 149054
rect 244464 148990 244516 148996
rect 244280 144900 244332 144906
rect 244280 144842 244332 144848
rect 244936 129674 244964 168370
rect 245108 151836 245160 151842
rect 245108 151778 245160 151784
rect 245016 135380 245068 135386
rect 245016 135322 245068 135328
rect 244924 129668 244976 129674
rect 244924 129610 244976 129616
rect 243728 122120 243780 122126
rect 243728 122062 243780 122068
rect 243636 121508 243688 121514
rect 243636 121450 243688 121456
rect 243544 76696 243596 76702
rect 243544 76638 243596 76644
rect 242440 73908 242492 73914
rect 242440 73850 242492 73856
rect 243648 68338 243676 121450
rect 244924 111852 244976 111858
rect 244924 111794 244976 111800
rect 243728 107772 243780 107778
rect 243728 107714 243780 107720
rect 243740 74050 243768 107714
rect 243728 74044 243780 74050
rect 243728 73986 243780 73992
rect 243636 68332 243688 68338
rect 243636 68274 243688 68280
rect 242348 66904 242400 66910
rect 242348 66846 242400 66852
rect 244936 18630 244964 111794
rect 245028 72554 245056 135322
rect 245120 110294 245148 151778
rect 245200 146396 245252 146402
rect 245200 146338 245252 146344
rect 245108 110288 245160 110294
rect 245108 110230 245160 110236
rect 245212 106146 245240 146338
rect 245672 139398 245700 195298
rect 245752 184340 245804 184346
rect 245752 184282 245804 184288
rect 245764 153134 245792 184282
rect 246408 182850 246436 256527
rect 246488 254584 246540 254590
rect 246488 254526 246540 254532
rect 246500 246537 246528 254526
rect 246486 246528 246542 246537
rect 246486 246463 246542 246472
rect 246396 182844 246448 182850
rect 246396 182786 246448 182792
rect 246396 175296 246448 175302
rect 246396 175238 246448 175244
rect 246304 163056 246356 163062
rect 246304 162998 246356 163004
rect 245752 153128 245804 153134
rect 245752 153070 245804 153076
rect 245660 139392 245712 139398
rect 245660 139334 245712 139340
rect 246316 129062 246344 162998
rect 246304 129056 246356 129062
rect 246304 128998 246356 129004
rect 246304 121576 246356 121582
rect 246304 121518 246356 121524
rect 245200 106140 245252 106146
rect 245200 106082 245252 106088
rect 245108 98116 245160 98122
rect 245108 98058 245160 98064
rect 245016 72548 245068 72554
rect 245016 72490 245068 72496
rect 245120 53106 245148 98058
rect 245108 53100 245160 53106
rect 245108 53042 245160 53048
rect 244924 18624 244976 18630
rect 244924 18566 244976 18572
rect 246316 11830 246344 121518
rect 246408 106962 246436 175238
rect 247052 168298 247080 291246
rect 249076 275398 249104 698906
rect 249984 305040 250036 305046
rect 249984 304982 250036 304988
rect 249800 288652 249852 288658
rect 249800 288594 249852 288600
rect 249156 284572 249208 284578
rect 249156 284514 249208 284520
rect 249064 275392 249116 275398
rect 249064 275334 249116 275340
rect 247130 270192 247186 270201
rect 247130 270127 247186 270136
rect 247144 173874 247172 270127
rect 248420 263628 248472 263634
rect 248420 263570 248472 263576
rect 247224 181620 247276 181626
rect 247224 181562 247276 181568
rect 247132 173868 247184 173874
rect 247132 173810 247184 173816
rect 247040 168292 247092 168298
rect 247040 168234 247092 168240
rect 246580 149728 246632 149734
rect 246580 149670 246632 149676
rect 246488 128376 246540 128382
rect 246488 128318 246540 128324
rect 246396 106956 246448 106962
rect 246396 106898 246448 106904
rect 246500 83502 246528 128318
rect 246592 111722 246620 149670
rect 247236 146266 247264 181562
rect 247960 173188 248012 173194
rect 247960 173130 248012 173136
rect 247868 161560 247920 161566
rect 247868 161502 247920 161508
rect 247224 146260 247276 146266
rect 247224 146202 247276 146208
rect 247776 145104 247828 145110
rect 247776 145046 247828 145052
rect 247684 134088 247736 134094
rect 247684 134030 247736 134036
rect 246580 111716 246632 111722
rect 246580 111658 246632 111664
rect 246580 107840 246632 107846
rect 246580 107782 246632 107788
rect 246488 83496 246540 83502
rect 246488 83438 246540 83444
rect 246592 65550 246620 107782
rect 246580 65544 246632 65550
rect 246580 65486 246632 65492
rect 247696 33794 247724 134030
rect 247788 103494 247816 145046
rect 247880 121446 247908 161502
rect 247972 135182 248000 173130
rect 248432 172446 248460 263570
rect 249168 259418 249196 284514
rect 249156 259412 249208 259418
rect 249156 259354 249208 259360
rect 248512 187060 248564 187066
rect 248512 187002 248564 187008
rect 248420 172440 248472 172446
rect 248420 172382 248472 172388
rect 248524 152590 248552 187002
rect 249156 171148 249208 171154
rect 249156 171090 249208 171096
rect 248512 152584 248564 152590
rect 248512 152526 248564 152532
rect 249064 150476 249116 150482
rect 249064 150418 249116 150424
rect 247960 135176 248012 135182
rect 247960 135118 248012 135124
rect 247868 121440 247920 121446
rect 247868 121382 247920 121388
rect 247868 117360 247920 117366
rect 247868 117302 247920 117308
rect 247776 103488 247828 103494
rect 247776 103430 247828 103436
rect 247880 87786 247908 117302
rect 249076 109002 249104 150418
rect 249168 132394 249196 171090
rect 249340 154692 249392 154698
rect 249340 154634 249392 154640
rect 249248 144220 249300 144226
rect 249248 144162 249300 144168
rect 249156 132388 249208 132394
rect 249156 132330 249208 132336
rect 249156 114572 249208 114578
rect 249156 114514 249208 114520
rect 249064 108996 249116 109002
rect 249064 108938 249116 108944
rect 249064 106412 249116 106418
rect 249064 106354 249116 106360
rect 247868 87780 247920 87786
rect 247868 87722 247920 87728
rect 247684 33788 247736 33794
rect 247684 33730 247736 33736
rect 246304 11824 246356 11830
rect 246304 11766 246356 11772
rect 249076 10334 249104 106354
rect 249168 64190 249196 114514
rect 249260 104718 249288 144162
rect 249352 115870 249380 154634
rect 249812 149802 249840 288594
rect 249892 284640 249944 284646
rect 249892 284582 249944 284588
rect 249904 165578 249932 284582
rect 249996 278186 250024 304982
rect 251180 292732 251232 292738
rect 251180 292674 251232 292680
rect 249984 278180 250036 278186
rect 249984 278122 250036 278128
rect 250444 171216 250496 171222
rect 250444 171158 250496 171164
rect 249892 165572 249944 165578
rect 249892 165514 249944 165520
rect 249800 149796 249852 149802
rect 249800 149738 249852 149744
rect 250456 132462 250484 171158
rect 251192 171086 251220 292674
rect 251272 264988 251324 264994
rect 251272 264930 251324 264936
rect 251180 171080 251232 171086
rect 251180 171022 251232 171028
rect 250720 164892 250772 164898
rect 250720 164834 250772 164840
rect 250628 151156 250680 151162
rect 250628 151098 250680 151104
rect 250536 147688 250588 147694
rect 250536 147630 250588 147636
rect 250444 132456 250496 132462
rect 250444 132398 250496 132404
rect 249340 115864 249392 115870
rect 249340 115806 249392 115812
rect 250548 106214 250576 147630
rect 250640 113082 250668 151098
rect 250732 126886 250760 164834
rect 251284 153202 251312 264930
rect 252572 249762 252600 700334
rect 267660 697678 267688 703520
rect 283852 700398 283880 703520
rect 269764 700392 269816 700398
rect 269764 700334 269816 700340
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 266360 697672 266412 697678
rect 266360 697614 266412 697620
rect 267648 697672 267700 697678
rect 267648 697614 267700 697620
rect 258080 463004 258132 463010
rect 258080 462946 258132 462952
rect 253940 290080 253992 290086
rect 253940 290022 253992 290028
rect 253204 286000 253256 286006
rect 253204 285942 253256 285948
rect 252652 253972 252704 253978
rect 252652 253914 252704 253920
rect 252560 249756 252612 249762
rect 252560 249698 252612 249704
rect 251364 244316 251416 244322
rect 251364 244258 251416 244264
rect 251376 168366 251404 244258
rect 252100 173936 252152 173942
rect 252100 173878 252152 173884
rect 251364 168360 251416 168366
rect 251364 168302 251416 168308
rect 251824 166388 251876 166394
rect 251824 166330 251876 166336
rect 251272 153196 251324 153202
rect 251272 153138 251324 153144
rect 250812 131776 250864 131782
rect 250812 131718 250864 131724
rect 250720 126880 250772 126886
rect 250720 126822 250772 126828
rect 250720 123004 250772 123010
rect 250720 122946 250772 122952
rect 250628 113076 250680 113082
rect 250628 113018 250680 113024
rect 250536 106208 250588 106214
rect 250536 106150 250588 106156
rect 250444 104916 250496 104922
rect 250444 104858 250496 104864
rect 249248 104712 249300 104718
rect 249248 104654 249300 104660
rect 249340 103556 249392 103562
rect 249340 103498 249392 103504
rect 249248 100768 249300 100774
rect 249248 100710 249300 100716
rect 249260 76566 249288 100710
rect 249352 94722 249380 103498
rect 249340 94716 249392 94722
rect 249340 94658 249392 94664
rect 249248 76560 249300 76566
rect 249248 76502 249300 76508
rect 249156 64184 249208 64190
rect 249156 64126 249208 64132
rect 250456 15910 250484 104858
rect 250536 99476 250588 99482
rect 250536 99418 250588 99424
rect 250548 57254 250576 99418
rect 250732 87650 250760 122946
rect 250824 106282 250852 131718
rect 251836 126954 251864 166330
rect 252008 153332 252060 153338
rect 252008 153274 252060 153280
rect 251916 151904 251968 151910
rect 251916 151846 251968 151852
rect 251824 126948 251876 126954
rect 251824 126890 251876 126896
rect 251824 111920 251876 111926
rect 251824 111862 251876 111868
rect 250812 106276 250864 106282
rect 250812 106218 250864 106224
rect 250720 87644 250772 87650
rect 250720 87586 250772 87592
rect 251836 71126 251864 111862
rect 251928 111790 251956 151846
rect 252020 113150 252048 153274
rect 252112 151094 252140 173878
rect 252664 166326 252692 253914
rect 253216 181626 253244 285942
rect 253204 181620 253256 181626
rect 253204 181562 253256 181568
rect 253480 168496 253532 168502
rect 253480 168438 253532 168444
rect 252652 166320 252704 166326
rect 252652 166262 252704 166268
rect 253296 165708 253348 165714
rect 253296 165650 253348 165656
rect 252100 151088 252152 151094
rect 252100 151030 252152 151036
rect 253204 149184 253256 149190
rect 253204 149126 253256 149132
rect 252100 140956 252152 140962
rect 252100 140898 252152 140904
rect 252008 113144 252060 113150
rect 252008 113086 252060 113092
rect 251916 111784 251968 111790
rect 251916 111726 251968 111732
rect 252112 101454 252140 140898
rect 252192 124364 252244 124370
rect 252192 124306 252244 124312
rect 252100 101448 252152 101454
rect 252100 101390 252152 101396
rect 252204 86290 252232 124306
rect 253216 107574 253244 149126
rect 253308 125526 253336 165650
rect 253388 153876 253440 153882
rect 253388 153818 253440 153824
rect 253296 125520 253348 125526
rect 253296 125462 253348 125468
rect 253400 114510 253428 153818
rect 253492 129742 253520 168438
rect 253952 150414 253980 290022
rect 255964 288584 256016 288590
rect 255964 288526 256016 288532
rect 255320 287428 255372 287434
rect 255320 287370 255372 287376
rect 254032 281580 254084 281586
rect 254032 281522 254084 281528
rect 254044 160002 254072 281522
rect 254768 168564 254820 168570
rect 254768 168506 254820 168512
rect 254032 159996 254084 160002
rect 254032 159938 254084 159944
rect 253940 150408 253992 150414
rect 253940 150350 253992 150356
rect 254676 138100 254728 138106
rect 254676 138042 254728 138048
rect 254584 129804 254636 129810
rect 254584 129746 254636 129752
rect 253480 129736 253532 129742
rect 253480 129678 253532 129684
rect 253572 127628 253624 127634
rect 253572 127570 253624 127576
rect 253480 116204 253532 116210
rect 253480 116146 253532 116152
rect 253388 114504 253440 114510
rect 253388 114446 253440 114452
rect 253296 109132 253348 109138
rect 253296 109074 253348 109080
rect 253204 107568 253256 107574
rect 253204 107510 253256 107516
rect 253204 103624 253256 103630
rect 253204 103566 253256 103572
rect 252192 86284 252244 86290
rect 252192 86226 252244 86232
rect 251824 71120 251876 71126
rect 251824 71062 251876 71068
rect 250536 57248 250588 57254
rect 250536 57190 250588 57196
rect 250444 15904 250496 15910
rect 250444 15846 250496 15852
rect 253216 14482 253244 103566
rect 253308 78062 253336 109074
rect 253492 89010 253520 116146
rect 253584 102134 253612 127570
rect 253572 102128 253624 102134
rect 253572 102070 253624 102076
rect 253480 89004 253532 89010
rect 253480 88946 253532 88952
rect 253296 78056 253348 78062
rect 253296 77998 253348 78004
rect 254596 55894 254624 129746
rect 254688 90506 254716 138042
rect 254780 130966 254808 168506
rect 254860 157480 254912 157486
rect 254860 157422 254912 157428
rect 254768 130960 254820 130966
rect 254768 130902 254820 130908
rect 254768 125724 254820 125730
rect 254768 125666 254820 125672
rect 254676 90500 254728 90506
rect 254676 90442 254728 90448
rect 254780 79490 254808 125666
rect 254872 117298 254900 157422
rect 255332 157350 255360 287370
rect 255412 271992 255464 271998
rect 255412 271934 255464 271940
rect 255424 160070 255452 271934
rect 255976 250510 256004 288526
rect 256700 273352 256752 273358
rect 256700 273294 256752 273300
rect 255964 250504 256016 250510
rect 255964 250446 256016 250452
rect 255504 240372 255556 240378
rect 255504 240314 255556 240320
rect 255516 175166 255544 240314
rect 256712 175234 256740 273294
rect 258092 252550 258120 462946
rect 266372 302258 266400 697614
rect 260196 302252 260248 302258
rect 260196 302194 260248 302200
rect 266360 302252 266412 302258
rect 266360 302194 266412 302200
rect 260104 289944 260156 289950
rect 260104 289886 260156 289892
rect 258172 270632 258224 270638
rect 258172 270574 258224 270580
rect 258080 252544 258132 252550
rect 258080 252486 258132 252492
rect 256700 175228 256752 175234
rect 256700 175170 256752 175176
rect 255504 175160 255556 175166
rect 255504 175102 255556 175108
rect 257436 174072 257488 174078
rect 257436 174014 257488 174020
rect 256148 174004 256200 174010
rect 256148 173946 256200 173952
rect 255412 160064 255464 160070
rect 255412 160006 255464 160012
rect 255320 157344 255372 157350
rect 255320 157286 255372 157292
rect 255964 156120 256016 156126
rect 255964 156062 256016 156068
rect 254860 117292 254912 117298
rect 254860 117234 254912 117240
rect 255976 115938 256004 156062
rect 256056 146940 256108 146946
rect 256056 146882 256108 146888
rect 255964 115932 256016 115938
rect 255964 115874 256016 115880
rect 256068 107642 256096 146882
rect 256160 135250 256188 173946
rect 257344 169856 257396 169862
rect 257344 169798 257396 169804
rect 256240 142316 256292 142322
rect 256240 142258 256292 142264
rect 256148 135244 256200 135250
rect 256148 135186 256200 135192
rect 256148 110560 256200 110566
rect 256148 110502 256200 110508
rect 256056 107636 256108 107642
rect 256056 107578 256108 107584
rect 256056 103692 256108 103698
rect 256056 103634 256108 103640
rect 255964 102332 256016 102338
rect 255964 102274 256016 102280
rect 254768 79484 254820 79490
rect 254768 79426 254820 79432
rect 254584 55888 254636 55894
rect 254584 55830 254636 55836
rect 255976 22778 256004 102274
rect 256068 51814 256096 103634
rect 256160 79422 256188 110502
rect 256252 104242 256280 142258
rect 257356 131034 257384 169798
rect 257448 148374 257476 174014
rect 257620 158840 257672 158846
rect 257620 158782 257672 158788
rect 257436 148368 257488 148374
rect 257436 148310 257488 148316
rect 257436 135448 257488 135454
rect 257436 135390 257488 135396
rect 257344 131028 257396 131034
rect 257344 130970 257396 130976
rect 257344 128444 257396 128450
rect 257344 128386 257396 128392
rect 256332 121644 256384 121650
rect 256332 121586 256384 121592
rect 256240 104236 256292 104242
rect 256240 104178 256292 104184
rect 256344 94654 256372 121586
rect 256332 94648 256384 94654
rect 256332 94590 256384 94596
rect 256148 79416 256200 79422
rect 256148 79358 256200 79364
rect 257356 54534 257384 128386
rect 257448 89078 257476 135390
rect 257528 125792 257580 125798
rect 257528 125734 257580 125740
rect 257436 89072 257488 89078
rect 257436 89014 257488 89020
rect 257540 84833 257568 125734
rect 257632 120766 257660 158782
rect 258184 142118 258212 270574
rect 259460 262268 259512 262274
rect 259460 262210 259512 262216
rect 258264 260908 258316 260914
rect 258264 260850 258316 260856
rect 258276 162858 258304 260850
rect 259472 172514 259500 262210
rect 260116 180266 260144 289886
rect 260208 238474 260236 302194
rect 264244 296744 264296 296750
rect 264244 296686 264296 296692
rect 260840 290012 260892 290018
rect 260840 289954 260892 289960
rect 260196 238468 260248 238474
rect 260196 238410 260248 238416
rect 260104 180260 260156 180266
rect 260104 180202 260156 180208
rect 260380 172576 260432 172582
rect 260380 172518 260432 172524
rect 259460 172508 259512 172514
rect 259460 172450 259512 172456
rect 258816 169924 258868 169930
rect 258816 169866 258868 169872
rect 258264 162852 258316 162858
rect 258264 162794 258316 162800
rect 258724 158908 258776 158914
rect 258724 158850 258776 158856
rect 258172 142112 258224 142118
rect 258172 142054 258224 142060
rect 257620 120760 257672 120766
rect 257620 120702 257672 120708
rect 258736 118590 258764 158850
rect 258828 131102 258856 169866
rect 260288 168632 260340 168638
rect 260288 168574 260340 168580
rect 260104 160268 260156 160274
rect 260104 160210 260156 160216
rect 258908 157548 258960 157554
rect 258908 157490 258960 157496
rect 258816 131096 258868 131102
rect 258816 131038 258868 131044
rect 258816 118720 258868 118726
rect 258816 118662 258868 118668
rect 258724 118584 258776 118590
rect 258724 118526 258776 118532
rect 258724 116068 258776 116074
rect 258724 116010 258776 116016
rect 257526 84824 257582 84833
rect 257526 84759 257582 84768
rect 257344 54528 257396 54534
rect 257344 54470 257396 54476
rect 256056 51808 256108 51814
rect 256056 51750 256108 51756
rect 258736 42090 258764 116010
rect 258828 72486 258856 118662
rect 258920 118658 258948 157490
rect 260116 120086 260144 160210
rect 260196 132864 260248 132870
rect 260196 132806 260248 132812
rect 260104 120080 260156 120086
rect 260104 120022 260156 120028
rect 258908 118652 258960 118658
rect 258908 118594 258960 118600
rect 260104 116136 260156 116142
rect 260104 116078 260156 116084
rect 258908 111988 258960 111994
rect 258908 111930 258960 111936
rect 258920 93158 258948 111930
rect 259000 105052 259052 105058
rect 259000 104994 259052 105000
rect 258908 93152 258960 93158
rect 258908 93094 258960 93100
rect 259012 90438 259040 104994
rect 259000 90432 259052 90438
rect 259000 90374 259052 90380
rect 258816 72480 258868 72486
rect 258816 72422 258868 72428
rect 258724 42084 258776 42090
rect 258724 42026 258776 42032
rect 255964 22772 256016 22778
rect 255964 22714 256016 22720
rect 260116 17270 260144 116078
rect 260208 69698 260236 132806
rect 260300 128246 260328 168574
rect 260392 133822 260420 172518
rect 260472 147824 260524 147830
rect 260472 147766 260524 147772
rect 260380 133816 260432 133822
rect 260380 133758 260432 133764
rect 260288 128240 260340 128246
rect 260288 128182 260340 128188
rect 260484 111110 260512 147766
rect 260852 140758 260880 289954
rect 262864 285932 262916 285938
rect 262864 285874 262916 285880
rect 261484 284504 261536 284510
rect 261484 284446 261536 284452
rect 261496 185706 261524 284446
rect 261484 185700 261536 185706
rect 261484 185642 261536 185648
rect 262876 181762 262904 285874
rect 264256 182889 264284 296686
rect 265624 288516 265676 288522
rect 265624 288458 265676 288464
rect 264336 284708 264388 284714
rect 264336 284650 264388 284656
rect 264242 182880 264298 182889
rect 264242 182815 264298 182824
rect 262864 181756 262916 181762
rect 262864 181698 262916 181704
rect 264348 177313 264376 284650
rect 265636 178673 265664 288458
rect 267004 287360 267056 287366
rect 267004 287302 267056 287308
rect 267016 181694 267044 287302
rect 268384 280288 268436 280294
rect 268384 280230 268436 280236
rect 267096 271924 267148 271930
rect 267096 271866 267148 271872
rect 267004 181688 267056 181694
rect 267004 181630 267056 181636
rect 267108 178838 267136 271866
rect 268396 178974 268424 280230
rect 268476 267844 268528 267850
rect 268476 267786 268528 267792
rect 268384 178968 268436 178974
rect 268384 178910 268436 178916
rect 267096 178832 267148 178838
rect 267096 178774 267148 178780
rect 265622 178664 265678 178673
rect 265622 178599 265678 178608
rect 264334 177304 264390 177313
rect 264334 177239 264390 177248
rect 268488 175982 268516 267786
rect 269776 240310 269804 700334
rect 299492 623082 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 660346 331260 702986
rect 348804 696250 348832 703520
rect 364996 699718 365024 703520
rect 395344 700392 395396 700398
rect 395344 700334 395396 700340
rect 363604 699712 363656 699718
rect 363604 699654 363656 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 348792 696244 348844 696250
rect 348792 696186 348844 696192
rect 331220 660340 331272 660346
rect 331220 660282 331272 660288
rect 299480 623076 299532 623082
rect 299480 623018 299532 623024
rect 309784 430636 309836 430642
rect 309784 430578 309836 430584
rect 305644 364404 305696 364410
rect 305644 364346 305696 364352
rect 273904 294024 273956 294030
rect 273904 293966 273956 293972
rect 271144 291236 271196 291242
rect 271144 291178 271196 291184
rect 269856 266416 269908 266422
rect 269856 266358 269908 266364
rect 269764 240304 269816 240310
rect 269764 240246 269816 240252
rect 269868 177478 269896 266358
rect 269948 241596 270000 241602
rect 269948 241538 270000 241544
rect 269960 179042 269988 241538
rect 269948 179036 270000 179042
rect 269948 178978 270000 178984
rect 269856 177472 269908 177478
rect 271156 177449 271184 291178
rect 271236 280220 271288 280226
rect 271236 280162 271288 280168
rect 271248 178906 271276 280162
rect 272524 256760 272576 256766
rect 272524 256702 272576 256708
rect 271328 193860 271380 193866
rect 271328 193802 271380 193808
rect 271236 178900 271288 178906
rect 271236 178842 271288 178848
rect 271340 177614 271368 193802
rect 272536 182918 272564 256702
rect 272524 182912 272576 182918
rect 272524 182854 272576 182860
rect 273916 180334 273944 293966
rect 305000 292664 305052 292670
rect 305000 292606 305052 292612
rect 302884 287292 302936 287298
rect 302884 287234 302936 287240
rect 302240 287088 302292 287094
rect 302240 287030 302292 287036
rect 276664 285864 276716 285870
rect 276664 285806 276716 285812
rect 298098 285832 298154 285841
rect 273996 242956 274048 242962
rect 273996 242898 274048 242904
rect 273904 180328 273956 180334
rect 273904 180270 273956 180276
rect 271328 177608 271380 177614
rect 271328 177550 271380 177556
rect 269856 177414 269908 177420
rect 271142 177440 271198 177449
rect 271142 177375 271198 177384
rect 274008 176050 274036 242898
rect 276676 176118 276704 285806
rect 291200 285796 291252 285802
rect 298098 285767 298154 285776
rect 291200 285738 291252 285744
rect 284300 283892 284352 283898
rect 284300 283834 284352 283840
rect 282920 283620 282972 283626
rect 282920 283562 282972 283568
rect 280804 276072 280856 276078
rect 280804 276014 280856 276020
rect 276756 270564 276808 270570
rect 276756 270506 276808 270512
rect 276768 176186 276796 270506
rect 278044 231192 278096 231198
rect 278044 231134 278096 231140
rect 276848 228404 276900 228410
rect 276848 228346 276900 228352
rect 276860 176662 276888 228346
rect 276848 176656 276900 176662
rect 276848 176598 276900 176604
rect 278056 176526 278084 231134
rect 280160 210452 280212 210458
rect 280160 210394 280212 210400
rect 279056 196648 279108 196654
rect 279056 196590 279108 196596
rect 278780 189848 278832 189854
rect 278780 189790 278832 189796
rect 278136 184408 278188 184414
rect 278136 184350 278188 184356
rect 278148 177546 278176 184350
rect 278136 177540 278188 177546
rect 278136 177482 278188 177488
rect 278044 176520 278096 176526
rect 278044 176462 278096 176468
rect 276756 176180 276808 176186
rect 276756 176122 276808 176128
rect 276664 176112 276716 176118
rect 278792 176089 278820 189790
rect 276664 176054 276716 176060
rect 278778 176080 278834 176089
rect 273996 176044 274048 176050
rect 278778 176015 278834 176024
rect 273996 175986 274048 175992
rect 268476 175976 268528 175982
rect 268476 175918 268528 175924
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175302 265020 175607
rect 264980 175296 265032 175302
rect 264980 175238 265032 175244
rect 265254 175264 265310 175273
rect 265254 175199 265310 175208
rect 264978 174856 265034 174865
rect 264978 174791 265034 174800
rect 264992 174078 265020 174791
rect 265070 174448 265126 174457
rect 265070 174383 265126 174392
rect 264980 174072 265032 174078
rect 264980 174014 265032 174020
rect 265084 174010 265112 174383
rect 265162 174040 265218 174049
rect 265072 174004 265124 174010
rect 265162 173975 265218 173984
rect 265072 173946 265124 173952
rect 264978 173632 265034 173641
rect 264978 173567 265034 173576
rect 264992 172718 265020 173567
rect 265176 173194 265204 173975
rect 265268 173942 265296 175199
rect 265256 173936 265308 173942
rect 265256 173878 265308 173884
rect 265164 173188 265216 173194
rect 265164 173130 265216 173136
rect 265070 173088 265126 173097
rect 265070 173023 265126 173032
rect 264980 172712 265032 172718
rect 264518 172680 264574 172689
rect 264980 172654 265032 172660
rect 264518 172615 264574 172624
rect 262956 171556 263008 171562
rect 262956 171498 263008 171504
rect 261760 167136 261812 167142
rect 261760 167078 261812 167084
rect 261484 164348 261536 164354
rect 261484 164290 261536 164296
rect 260840 140752 260892 140758
rect 260840 140694 260892 140700
rect 261496 125594 261524 164290
rect 261668 129872 261720 129878
rect 261668 129814 261720 129820
rect 261576 127016 261628 127022
rect 261576 126958 261628 126964
rect 261484 125588 261536 125594
rect 261484 125530 261536 125536
rect 261484 117428 261536 117434
rect 261484 117370 261536 117376
rect 260472 111104 260524 111110
rect 260472 111046 260524 111052
rect 260380 110628 260432 110634
rect 260380 110570 260432 110576
rect 260288 109200 260340 109206
rect 260288 109142 260340 109148
rect 260196 69692 260248 69698
rect 260196 69634 260248 69640
rect 260300 62898 260328 109142
rect 260392 91866 260420 110570
rect 261300 100904 261352 100910
rect 261300 100846 261352 100852
rect 261312 94586 261340 100846
rect 261300 94580 261352 94586
rect 261300 94522 261352 94528
rect 260380 91860 260432 91866
rect 260380 91802 260432 91808
rect 260288 62892 260340 62898
rect 260288 62834 260340 62840
rect 261496 26926 261524 117370
rect 261588 73846 261616 126958
rect 261680 84862 261708 129814
rect 261772 128314 261800 167078
rect 262864 147892 262916 147898
rect 262864 147834 262916 147840
rect 261852 132796 261904 132802
rect 261852 132738 261904 132744
rect 261760 128308 261812 128314
rect 261760 128250 261812 128256
rect 261864 116618 261892 132738
rect 261852 116612 261904 116618
rect 261852 116554 261904 116560
rect 262876 110362 262904 147834
rect 262968 133890 262996 171498
rect 264242 162888 264298 162897
rect 264242 162823 264298 162832
rect 263048 149252 263100 149258
rect 263048 149194 263100 149200
rect 262956 133884 263008 133890
rect 262956 133826 263008 133832
rect 262956 116000 263008 116006
rect 262956 115942 263008 115948
rect 262864 110356 262916 110362
rect 262864 110298 262916 110304
rect 262968 104174 262996 115942
rect 263060 113830 263088 149194
rect 263140 132660 263192 132666
rect 263140 132602 263192 132608
rect 263048 113824 263100 113830
rect 263048 113766 263100 113772
rect 263048 104984 263100 104990
rect 263048 104926 263100 104932
rect 262956 104168 263008 104174
rect 262956 104110 263008 104116
rect 262864 102196 262916 102202
rect 262864 102138 262916 102144
rect 261668 84856 261720 84862
rect 261668 84798 261720 84804
rect 261576 73840 261628 73846
rect 261576 73782 261628 73788
rect 261484 26920 261536 26926
rect 261484 26862 261536 26868
rect 260104 17264 260156 17270
rect 260104 17206 260156 17212
rect 253204 14476 253256 14482
rect 253204 14418 253256 14424
rect 262876 11762 262904 102138
rect 262956 100836 263008 100842
rect 262956 100778 263008 100784
rect 262968 75206 262996 100778
rect 263060 91798 263088 104926
rect 263152 100706 263180 132602
rect 264256 122806 264284 162823
rect 264428 147756 264480 147762
rect 264428 147698 264480 147704
rect 264334 135280 264390 135289
rect 264334 135215 264390 135224
rect 264244 122800 264296 122806
rect 264244 122742 264296 122748
rect 264242 118960 264298 118969
rect 264242 118895 264298 118904
rect 263140 100700 263192 100706
rect 263140 100642 263192 100648
rect 263048 91792 263100 91798
rect 263048 91734 263100 91740
rect 262956 75200 263008 75206
rect 262956 75142 263008 75148
rect 262864 11756 262916 11762
rect 262864 11698 262916 11704
rect 249064 10328 249116 10334
rect 249064 10270 249116 10276
rect 242164 7608 242216 7614
rect 242164 7550 242216 7556
rect 233884 3052 233936 3058
rect 233884 2994 233936 3000
rect 235816 3052 235868 3058
rect 235816 2994 235868 3000
rect 235828 480 235856 2994
rect 264256 2106 264284 118895
rect 264348 71058 264376 135215
rect 264440 110430 264468 147698
rect 264532 135930 264560 172615
rect 265084 172582 265112 173023
rect 265072 172576 265124 172582
rect 265072 172518 265124 172524
rect 264978 172272 265034 172281
rect 264978 172207 265034 172216
rect 264992 171562 265020 172207
rect 265070 171864 265126 171873
rect 265070 171799 265126 171808
rect 264980 171556 265032 171562
rect 264980 171498 265032 171504
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171154 265020 171391
rect 265084 171222 265112 171799
rect 265072 171216 265124 171222
rect 265072 171158 265124 171164
rect 264980 171148 265032 171154
rect 264980 171090 265032 171096
rect 265070 171048 265126 171057
rect 265070 170983 265126 170992
rect 264978 170096 265034 170105
rect 264978 170031 265034 170040
rect 264992 169862 265020 170031
rect 264980 169856 265032 169862
rect 264980 169798 265032 169804
rect 265084 169794 265112 170983
rect 265162 170504 265218 170513
rect 265162 170439 265218 170448
rect 265176 169930 265204 170439
rect 265164 169924 265216 169930
rect 265164 169866 265216 169872
rect 265072 169788 265124 169794
rect 265072 169730 265124 169736
rect 265070 169688 265126 169697
rect 265070 169623 265126 169632
rect 264978 169280 265034 169289
rect 264978 169215 265034 169224
rect 264992 168502 265020 169215
rect 265084 168570 265112 169623
rect 265162 168872 265218 168881
rect 265162 168807 265218 168816
rect 265072 168564 265124 168570
rect 265072 168506 265124 168512
rect 264980 168496 265032 168502
rect 264980 168438 265032 168444
rect 265176 168434 265204 168807
rect 265256 168632 265308 168638
rect 265256 168574 265308 168580
rect 265268 168473 265296 168574
rect 265254 168464 265310 168473
rect 265164 168428 265216 168434
rect 265254 168399 265310 168408
rect 265164 168370 265216 168376
rect 265162 167920 265218 167929
rect 265162 167855 265218 167864
rect 264978 167512 265034 167521
rect 264978 167447 265034 167456
rect 264992 167074 265020 167447
rect 265176 167142 265204 167855
rect 265164 167136 265216 167142
rect 265070 167104 265126 167113
rect 264980 167068 265032 167074
rect 265164 167078 265216 167084
rect 265070 167039 265126 167048
rect 264980 167010 265032 167016
rect 265084 166394 265112 167039
rect 265162 166696 265218 166705
rect 265162 166631 265218 166640
rect 265072 166388 265124 166394
rect 265072 166330 265124 166336
rect 265070 166288 265126 166297
rect 265070 166223 265126 166232
rect 264978 165880 265034 165889
rect 264978 165815 265034 165824
rect 264992 165714 265020 165815
rect 264980 165708 265032 165714
rect 264980 165650 265032 165656
rect 265084 165646 265112 166223
rect 265072 165640 265124 165646
rect 265072 165582 265124 165588
rect 264978 165336 265034 165345
rect 264978 165271 265034 165280
rect 264992 164286 265020 165271
rect 265070 164928 265126 164937
rect 265176 164898 265204 166631
rect 265070 164863 265126 164872
rect 265164 164892 265216 164898
rect 265084 164354 265112 164863
rect 265164 164834 265216 164840
rect 265622 164520 265678 164529
rect 265622 164455 265678 164464
rect 265072 164348 265124 164354
rect 265072 164290 265124 164296
rect 264980 164280 265032 164286
rect 264980 164222 265032 164228
rect 265162 164112 265218 164121
rect 265162 164047 265218 164056
rect 265070 163704 265126 163713
rect 265070 163639 265126 163648
rect 264978 163296 265034 163305
rect 264978 163231 265034 163240
rect 264992 162994 265020 163231
rect 265084 163062 265112 163639
rect 265176 163130 265204 164047
rect 265164 163124 265216 163130
rect 265164 163066 265216 163072
rect 265072 163056 265124 163062
rect 265072 162998 265124 163004
rect 264980 162988 265032 162994
rect 264980 162930 265032 162936
rect 265162 162344 265218 162353
rect 265162 162279 265218 162288
rect 264978 161936 265034 161945
rect 264978 161871 265034 161880
rect 264992 161566 265020 161871
rect 264980 161560 265032 161566
rect 264980 161502 265032 161508
rect 265070 161528 265126 161537
rect 264992 161472 265070 161474
rect 265176 161498 265204 162279
rect 264992 161463 265126 161472
rect 265164 161492 265216 161498
rect 264992 161446 265112 161463
rect 264992 160750 265020 161446
rect 265164 161434 265216 161440
rect 265070 161120 265126 161129
rect 265070 161055 265126 161064
rect 264980 160744 265032 160750
rect 264980 160686 265032 160692
rect 264978 160304 265034 160313
rect 264978 160239 265034 160248
rect 264992 160138 265020 160239
rect 265084 160206 265112 161055
rect 265162 160712 265218 160721
rect 265162 160647 265218 160656
rect 265176 160274 265204 160647
rect 265164 160268 265216 160274
rect 265164 160210 265216 160216
rect 265072 160200 265124 160206
rect 265072 160142 265124 160148
rect 264980 160132 265032 160138
rect 264980 160074 265032 160080
rect 265070 159760 265126 159769
rect 265070 159695 265126 159704
rect 264978 159352 265034 159361
rect 264978 159287 265034 159296
rect 264992 158778 265020 159287
rect 265084 158846 265112 159695
rect 265162 158944 265218 158953
rect 265162 158879 265164 158888
rect 265216 158879 265218 158888
rect 265164 158850 265216 158856
rect 265072 158840 265124 158846
rect 265072 158782 265124 158788
rect 264980 158772 265032 158778
rect 264980 158714 265032 158720
rect 265162 158536 265218 158545
rect 265162 158471 265218 158480
rect 265070 158128 265126 158137
rect 265070 158063 265126 158072
rect 264978 157720 265034 157729
rect 264978 157655 265034 157664
rect 264992 157418 265020 157655
rect 265084 157486 265112 158063
rect 265176 157554 265204 158471
rect 265164 157548 265216 157554
rect 265164 157490 265216 157496
rect 265072 157480 265124 157486
rect 265072 157422 265124 157428
rect 264980 157412 265032 157418
rect 264980 157354 265032 157360
rect 265162 157176 265218 157185
rect 265162 157111 265218 157120
rect 265070 156768 265126 156777
rect 265070 156703 265126 156712
rect 264978 156360 265034 156369
rect 264978 156295 265034 156304
rect 264992 156058 265020 156295
rect 265084 156126 265112 156703
rect 265072 156120 265124 156126
rect 265072 156062 265124 156068
rect 264980 156052 265032 156058
rect 264980 155994 265032 156000
rect 265176 155990 265204 157111
rect 265164 155984 265216 155990
rect 265070 155952 265126 155961
rect 265164 155926 265216 155932
rect 265070 155887 265126 155896
rect 264978 155544 265034 155553
rect 264978 155479 265034 155488
rect 264992 154630 265020 155479
rect 265084 154698 265112 155887
rect 265636 155242 265664 164455
rect 279068 155258 279096 196590
rect 279240 178764 279292 178770
rect 279240 178706 279292 178712
rect 279148 177404 279200 177410
rect 279148 177346 279200 177352
rect 279160 161474 279188 177346
rect 279252 171134 279280 178706
rect 279332 176180 279384 176186
rect 279332 176122 279384 176128
rect 279344 175273 279372 176122
rect 279330 175264 279386 175273
rect 279330 175199 279386 175208
rect 279252 171106 279372 171134
rect 279344 162217 279372 171106
rect 279330 162208 279386 162217
rect 279330 162143 279386 162152
rect 279160 161446 279464 161474
rect 279330 155272 279386 155281
rect 265624 155236 265676 155242
rect 279068 155230 279330 155258
rect 279330 155207 279386 155216
rect 265624 155178 265676 155184
rect 265162 155136 265218 155145
rect 265162 155071 265218 155080
rect 265072 154692 265124 154698
rect 265072 154634 265124 154640
rect 264980 154624 265032 154630
rect 264980 154566 265032 154572
rect 265070 154184 265126 154193
rect 265070 154119 265126 154128
rect 264978 153368 265034 153377
rect 265084 153338 265112 154119
rect 265176 153882 265204 155071
rect 265346 154592 265402 154601
rect 265346 154527 265402 154536
rect 265164 153876 265216 153882
rect 265164 153818 265216 153824
rect 265162 153776 265218 153785
rect 265162 153711 265218 153720
rect 264978 153303 265034 153312
rect 265072 153332 265124 153338
rect 264992 153270 265020 153303
rect 265072 153274 265124 153280
rect 264980 153264 265032 153270
rect 264980 153206 265032 153212
rect 265070 152960 265126 152969
rect 265070 152895 265126 152904
rect 264978 152008 265034 152017
rect 264978 151943 265034 151952
rect 264992 151842 265020 151943
rect 265084 151910 265112 152895
rect 265072 151904 265124 151910
rect 265072 151846 265124 151852
rect 264980 151836 265032 151842
rect 264980 151778 265032 151784
rect 265176 151162 265204 153711
rect 265254 152552 265310 152561
rect 265360 152522 265388 154527
rect 279436 153785 279464 161446
rect 279422 153776 279478 153785
rect 279422 153711 279478 153720
rect 265254 152487 265310 152496
rect 265348 152516 265400 152522
rect 265164 151156 265216 151162
rect 265164 151098 265216 151104
rect 264978 150784 265034 150793
rect 264978 150719 265034 150728
rect 264992 150482 265020 150719
rect 264980 150476 265032 150482
rect 264980 150418 265032 150424
rect 265070 150376 265126 150385
rect 265070 150311 265126 150320
rect 264978 149560 265034 149569
rect 264978 149495 265034 149504
rect 264992 149190 265020 149495
rect 264980 149184 265032 149190
rect 264980 149126 265032 149132
rect 265084 149122 265112 150311
rect 265268 149734 265296 152487
rect 265348 152458 265400 152464
rect 266082 151600 266138 151609
rect 266082 151535 266138 151544
rect 265346 151192 265402 151201
rect 265346 151127 265402 151136
rect 265256 149728 265308 149734
rect 265256 149670 265308 149676
rect 265072 149116 265124 149122
rect 265072 149058 265124 149064
rect 265070 149016 265126 149025
rect 265070 148951 265126 148960
rect 264978 148200 265034 148209
rect 264978 148135 265034 148144
rect 264992 147694 265020 148135
rect 265084 147830 265112 148951
rect 265162 148608 265218 148617
rect 265162 148543 265218 148552
rect 265072 147824 265124 147830
rect 265072 147766 265124 147772
rect 264980 147688 265032 147694
rect 264980 147630 265032 147636
rect 265070 147384 265126 147393
rect 265070 147319 265126 147328
rect 264978 146432 265034 146441
rect 265084 146402 265112 147319
rect 265176 146946 265204 148543
rect 265360 147898 265388 151127
rect 265438 149968 265494 149977
rect 265438 149903 265494 149912
rect 265452 149258 265480 149903
rect 265440 149252 265492 149258
rect 265440 149194 265492 149200
rect 265348 147892 265400 147898
rect 265348 147834 265400 147840
rect 265806 147792 265862 147801
rect 266096 147762 266124 151535
rect 265806 147727 265862 147736
rect 266084 147756 266136 147762
rect 265254 146976 265310 146985
rect 265164 146940 265216 146946
rect 265254 146911 265310 146920
rect 265164 146882 265216 146888
rect 264978 146367 265034 146376
rect 265072 146396 265124 146402
rect 264992 146334 265020 146367
rect 265072 146338 265124 146344
rect 264980 146328 265032 146334
rect 264980 146270 265032 146276
rect 265162 146024 265218 146033
rect 265162 145959 265218 145968
rect 265070 145616 265126 145625
rect 265070 145551 265126 145560
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 145042 265020 145143
rect 265084 145110 265112 145551
rect 265072 145104 265124 145110
rect 265072 145046 265124 145052
rect 264980 145036 265032 145042
rect 264980 144978 265032 144984
rect 265176 144974 265204 145959
rect 265164 144968 265216 144974
rect 265164 144910 265216 144916
rect 265070 144800 265126 144809
rect 265070 144735 265126 144744
rect 264978 144392 265034 144401
rect 264978 144327 265034 144336
rect 264992 143614 265020 144327
rect 265084 143682 265112 144735
rect 265268 144226 265296 146911
rect 265256 144220 265308 144226
rect 265256 144162 265308 144168
rect 265714 143848 265770 143857
rect 265714 143783 265770 143792
rect 265072 143676 265124 143682
rect 265072 143618 265124 143624
rect 264980 143608 265032 143614
rect 264980 143550 265032 143556
rect 265162 143440 265218 143449
rect 265162 143375 265218 143384
rect 264978 143032 265034 143041
rect 264978 142967 265034 142976
rect 264992 142322 265020 142967
rect 265070 142624 265126 142633
rect 265070 142559 265126 142568
rect 264980 142316 265032 142322
rect 264980 142258 265032 142264
rect 265084 142186 265112 142559
rect 265176 142254 265204 143375
rect 265164 142248 265216 142254
rect 265164 142190 265216 142196
rect 265072 142180 265124 142186
rect 265072 142122 265124 142128
rect 265070 141808 265126 141817
rect 265070 141743 265126 141752
rect 264980 140956 265032 140962
rect 264980 140898 265032 140904
rect 264992 140865 265020 140898
rect 265084 140894 265112 141743
rect 265162 141264 265218 141273
rect 265162 141199 265218 141208
rect 265072 140888 265124 140894
rect 264978 140856 265034 140865
rect 265072 140830 265124 140836
rect 265176 140826 265204 141199
rect 264978 140791 265034 140800
rect 265164 140820 265216 140826
rect 265164 140762 265216 140768
rect 264978 140040 265034 140049
rect 264978 139975 265034 139984
rect 264992 139466 265020 139975
rect 264980 139460 265032 139466
rect 264980 139402 265032 139408
rect 265070 139224 265126 139233
rect 265070 139159 265126 139168
rect 264978 138272 265034 138281
rect 264978 138207 265034 138216
rect 264992 138038 265020 138207
rect 265084 138106 265112 139159
rect 265072 138100 265124 138106
rect 265072 138042 265124 138048
rect 264980 138032 265032 138038
rect 264980 137974 265032 137980
rect 265254 137864 265310 137873
rect 265254 137799 265310 137808
rect 265070 137456 265126 137465
rect 265070 137391 265126 137400
rect 264978 137048 265034 137057
rect 264978 136983 265034 136992
rect 264992 136746 265020 136983
rect 265084 136814 265112 137391
rect 265072 136808 265124 136814
rect 265072 136750 265124 136756
rect 264980 136740 265032 136746
rect 264980 136682 265032 136688
rect 265268 136678 265296 137799
rect 265256 136672 265308 136678
rect 265162 136640 265218 136649
rect 265256 136614 265308 136620
rect 265162 136575 265218 136584
rect 265070 136232 265126 136241
rect 265070 136167 265126 136176
rect 264520 135924 264572 135930
rect 264520 135866 264572 135872
rect 264978 135688 265034 135697
rect 264978 135623 265034 135632
rect 264992 135386 265020 135623
rect 265084 135522 265112 136167
rect 265072 135516 265124 135522
rect 265072 135458 265124 135464
rect 265176 135454 265204 136575
rect 265164 135448 265216 135454
rect 265164 135390 265216 135396
rect 264980 135380 265032 135386
rect 264980 135322 265032 135328
rect 265162 134872 265218 134881
rect 265162 134807 265218 134816
rect 265070 134464 265126 134473
rect 265070 134399 265126 134408
rect 265084 134094 265112 134399
rect 265072 134088 265124 134094
rect 264978 134056 265034 134065
rect 265072 134030 265124 134036
rect 264978 133991 264980 134000
rect 265032 133991 265034 134000
rect 264980 133962 265032 133968
rect 265176 133958 265204 134807
rect 265164 133952 265216 133958
rect 265164 133894 265216 133900
rect 264978 133648 265034 133657
rect 264978 133583 265034 133592
rect 264992 132802 265020 133583
rect 265070 133104 265126 133113
rect 265070 133039 265126 133048
rect 265084 132870 265112 133039
rect 265072 132864 265124 132870
rect 265072 132806 265124 132812
rect 264980 132796 265032 132802
rect 264980 132738 265032 132744
rect 265622 132696 265678 132705
rect 265622 132631 265678 132640
rect 265070 130520 265126 130529
rect 265070 130455 265126 130464
rect 264978 130112 265034 130121
rect 264978 130047 265034 130056
rect 264992 129810 265020 130047
rect 265084 129878 265112 130455
rect 265072 129872 265124 129878
rect 265072 129814 265124 129820
rect 264980 129804 265032 129810
rect 264980 129746 265032 129752
rect 265070 129704 265126 129713
rect 265070 129639 265126 129648
rect 264978 129296 265034 129305
rect 264978 129231 265034 129240
rect 264992 128382 265020 129231
rect 265084 128450 265112 129639
rect 265072 128444 265124 128450
rect 265072 128386 265124 128392
rect 264980 128376 265032 128382
rect 264980 128318 265032 128324
rect 264978 127120 265034 127129
rect 264978 127055 265034 127064
rect 264992 127022 265020 127055
rect 264980 127016 265032 127022
rect 264980 126958 265032 126964
rect 265162 126712 265218 126721
rect 265162 126647 265218 126656
rect 265070 126304 265126 126313
rect 265070 126239 265126 126248
rect 264978 125896 265034 125905
rect 264978 125831 265034 125840
rect 264992 125798 265020 125831
rect 264980 125792 265032 125798
rect 264980 125734 265032 125740
rect 265084 125730 265112 126239
rect 265072 125724 265124 125730
rect 265072 125666 265124 125672
rect 265176 125662 265204 126647
rect 265164 125656 265216 125662
rect 265164 125598 265216 125604
rect 265162 125352 265218 125361
rect 265162 125287 265218 125296
rect 265070 124944 265126 124953
rect 265070 124879 265126 124888
rect 264978 124536 265034 124545
rect 264978 124471 265034 124480
rect 264992 124370 265020 124471
rect 264980 124364 265032 124370
rect 264980 124306 265032 124312
rect 265084 124302 265112 124879
rect 265072 124296 265124 124302
rect 265072 124238 265124 124244
rect 265176 124234 265204 125287
rect 265164 124228 265216 124234
rect 265164 124170 265216 124176
rect 265162 124128 265218 124137
rect 265162 124063 265218 124072
rect 265070 123720 265126 123729
rect 265070 123655 265126 123664
rect 264978 123312 265034 123321
rect 264978 123247 265034 123256
rect 264992 123010 265020 123247
rect 264980 123004 265032 123010
rect 264980 122946 265032 122952
rect 265084 122942 265112 123655
rect 265072 122936 265124 122942
rect 265072 122878 265124 122884
rect 265176 122874 265204 124063
rect 265164 122868 265216 122874
rect 265164 122810 265216 122816
rect 265070 122360 265126 122369
rect 265070 122295 265126 122304
rect 265084 121650 265112 122295
rect 265162 121952 265218 121961
rect 265162 121887 265218 121896
rect 265072 121644 265124 121650
rect 265072 121586 265124 121592
rect 264980 121576 265032 121582
rect 264978 121544 264980 121553
rect 265032 121544 265034 121553
rect 265176 121514 265204 121887
rect 264978 121479 265034 121488
rect 265164 121508 265216 121514
rect 265164 121450 265216 121456
rect 265162 121136 265218 121145
rect 265162 121071 265218 121080
rect 264978 120728 265034 120737
rect 264978 120663 265034 120672
rect 264992 120290 265020 120663
rect 265070 120320 265126 120329
rect 264980 120284 265032 120290
rect 265070 120255 265126 120264
rect 264980 120226 265032 120232
rect 265084 120154 265112 120255
rect 265176 120222 265204 121071
rect 265164 120216 265216 120222
rect 265164 120158 265216 120164
rect 265072 120148 265124 120154
rect 265072 120090 265124 120096
rect 264978 119776 265034 119785
rect 264978 119711 265034 119720
rect 264992 118726 265020 119711
rect 264980 118720 265032 118726
rect 264980 118662 265032 118668
rect 264978 118552 265034 118561
rect 264978 118487 265034 118496
rect 264992 117366 265020 118487
rect 265070 117736 265126 117745
rect 265070 117671 265126 117680
rect 265084 117434 265112 117671
rect 265072 117428 265124 117434
rect 265072 117370 265124 117376
rect 264980 117360 265032 117366
rect 264980 117302 265032 117308
rect 265162 117192 265218 117201
rect 265162 117127 265218 117136
rect 264978 116784 265034 116793
rect 264978 116719 265034 116728
rect 264992 116210 265020 116719
rect 265070 116376 265126 116385
rect 265070 116311 265126 116320
rect 264980 116204 265032 116210
rect 264980 116146 265032 116152
rect 264980 116068 265032 116074
rect 264980 116010 265032 116016
rect 264992 115977 265020 116010
rect 265084 116006 265112 116311
rect 265176 116142 265204 117127
rect 265164 116136 265216 116142
rect 265164 116078 265216 116084
rect 265072 116000 265124 116006
rect 264978 115968 265034 115977
rect 265072 115942 265124 115948
rect 264978 115903 265034 115912
rect 264978 115560 265034 115569
rect 264978 115495 265034 115504
rect 264992 114578 265020 115495
rect 264980 114572 265032 114578
rect 264980 114514 265032 114520
rect 265070 112976 265126 112985
rect 265070 112911 265126 112920
rect 264978 112568 265034 112577
rect 264978 112503 265034 112512
rect 264992 111926 265020 112503
rect 264980 111920 265032 111926
rect 264980 111862 265032 111868
rect 265084 111858 265112 112911
rect 265162 112024 265218 112033
rect 265162 111959 265164 111968
rect 265216 111959 265218 111968
rect 265164 111930 265216 111936
rect 265072 111852 265124 111858
rect 265072 111794 265124 111800
rect 265070 111616 265126 111625
rect 265070 111551 265126 111560
rect 264978 110800 265034 110809
rect 264978 110735 265034 110744
rect 264992 110566 265020 110735
rect 264980 110560 265032 110566
rect 264980 110502 265032 110508
rect 265084 110498 265112 111551
rect 265162 111208 265218 111217
rect 265162 111143 265218 111152
rect 265176 110634 265204 111143
rect 265164 110628 265216 110634
rect 265164 110570 265216 110576
rect 265072 110492 265124 110498
rect 265072 110434 265124 110440
rect 264428 110424 264480 110430
rect 264428 110366 264480 110372
rect 265070 110392 265126 110401
rect 265070 110327 265126 110336
rect 264978 109984 265034 109993
rect 264978 109919 265034 109928
rect 264992 109138 265020 109919
rect 264980 109132 265032 109138
rect 264980 109074 265032 109080
rect 265084 109070 265112 110327
rect 265162 109576 265218 109585
rect 265162 109511 265218 109520
rect 265176 109206 265204 109511
rect 265164 109200 265216 109206
rect 265164 109142 265216 109148
rect 265072 109064 265124 109070
rect 265072 109006 265124 109012
rect 265162 109032 265218 109041
rect 265162 108967 265218 108976
rect 265070 108624 265126 108633
rect 265070 108559 265126 108568
rect 264518 108216 264574 108225
rect 264518 108151 264574 108160
rect 264426 106448 264482 106457
rect 264426 106383 264482 106392
rect 264440 76634 264468 106383
rect 264532 87718 264560 108151
rect 265084 107914 265112 108559
rect 265072 107908 265124 107914
rect 265072 107850 265124 107856
rect 264980 107840 265032 107846
rect 264978 107808 264980 107817
rect 265032 107808 265034 107817
rect 265176 107778 265204 108967
rect 264978 107743 265034 107752
rect 265164 107772 265216 107778
rect 265164 107714 265216 107720
rect 265070 107400 265126 107409
rect 265070 107335 265126 107344
rect 264978 106992 265034 107001
rect 264978 106927 265034 106936
rect 264992 106486 265020 106927
rect 264980 106480 265032 106486
rect 264980 106422 265032 106428
rect 265084 106418 265112 107335
rect 265072 106412 265124 106418
rect 265072 106354 265124 106360
rect 265438 106040 265494 106049
rect 265438 105975 265494 105984
rect 264978 105632 265034 105641
rect 264978 105567 265034 105576
rect 264992 104922 265020 105567
rect 265070 105224 265126 105233
rect 265070 105159 265126 105168
rect 265084 105058 265112 105159
rect 265072 105052 265124 105058
rect 265072 104994 265124 105000
rect 265452 104990 265480 105975
rect 265440 104984 265492 104990
rect 265440 104926 265492 104932
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 265162 104816 265218 104825
rect 265162 104751 265218 104760
rect 265070 104408 265126 104417
rect 265070 104343 265126 104352
rect 264978 103864 265034 103873
rect 264978 103799 265034 103808
rect 264992 103562 265020 103799
rect 265084 103698 265112 104343
rect 265072 103692 265124 103698
rect 265072 103634 265124 103640
rect 265176 103630 265204 104751
rect 265164 103624 265216 103630
rect 265164 103566 265216 103572
rect 264980 103556 265032 103562
rect 264980 103498 265032 103504
rect 265254 103456 265310 103465
rect 265254 103391 265310 103400
rect 265070 103048 265126 103057
rect 265070 102983 265126 102992
rect 265084 102406 265112 102983
rect 265162 102640 265218 102649
rect 265162 102575 265218 102584
rect 265072 102400 265124 102406
rect 265072 102342 265124 102348
rect 264980 102332 265032 102338
rect 264980 102274 265032 102280
rect 264992 102241 265020 102274
rect 265176 102270 265204 102575
rect 265164 102264 265216 102270
rect 264978 102232 265034 102241
rect 265164 102206 265216 102212
rect 265268 102202 265296 103391
rect 264978 102167 265034 102176
rect 265256 102196 265308 102202
rect 265256 102138 265308 102144
rect 265346 101824 265402 101833
rect 265346 101759 265402 101768
rect 264978 101280 265034 101289
rect 264978 101215 265034 101224
rect 264992 100774 265020 101215
rect 265072 100904 265124 100910
rect 265070 100872 265072 100881
rect 265124 100872 265126 100881
rect 265360 100842 265388 101759
rect 265070 100807 265126 100816
rect 265348 100836 265400 100842
rect 265348 100778 265400 100784
rect 264980 100768 265032 100774
rect 264980 100710 265032 100716
rect 265070 100056 265126 100065
rect 265070 99991 265126 100000
rect 264978 99648 265034 99657
rect 264978 99583 265034 99592
rect 264992 99414 265020 99583
rect 265084 99482 265112 99991
rect 265072 99476 265124 99482
rect 265072 99418 265124 99424
rect 264980 99408 265032 99414
rect 264980 99350 265032 99356
rect 265070 99240 265126 99249
rect 265070 99175 265126 99184
rect 264978 98696 265034 98705
rect 264978 98631 265034 98640
rect 264992 98122 265020 98631
rect 264980 98116 265032 98122
rect 264980 98058 265032 98064
rect 265084 98054 265112 99175
rect 265072 98048 265124 98054
rect 265072 97990 265124 97996
rect 264978 97880 265034 97889
rect 264978 97815 265034 97824
rect 264992 97306 265020 97815
rect 265162 97472 265218 97481
rect 265162 97407 265218 97416
rect 264980 97300 265032 97306
rect 264980 97242 265032 97248
rect 265070 97064 265126 97073
rect 265070 96999 265126 97008
rect 264980 96824 265032 96830
rect 264980 96766 265032 96772
rect 264992 96665 265020 96766
rect 265084 96694 265112 96999
rect 265176 96762 265204 97407
rect 265164 96756 265216 96762
rect 265164 96698 265216 96704
rect 265072 96688 265124 96694
rect 264978 96656 265034 96665
rect 265072 96630 265124 96636
rect 264978 96591 265034 96600
rect 264978 96248 265034 96257
rect 264978 96183 265034 96192
rect 264992 95266 265020 96183
rect 264980 95260 265032 95266
rect 264980 95202 265032 95208
rect 264520 87712 264572 87718
rect 264520 87654 264572 87660
rect 265636 80714 265664 132631
rect 265728 127634 265756 143783
rect 265820 131782 265848 147727
rect 266084 147698 266136 147704
rect 265898 142216 265954 142225
rect 265898 142151 265954 142160
rect 265912 132666 265940 142151
rect 267278 138680 267334 138689
rect 267278 138615 267334 138624
rect 265900 132660 265952 132666
rect 265900 132602 265952 132608
rect 265808 131776 265860 131782
rect 265808 131718 265860 131724
rect 267094 131472 267150 131481
rect 267094 131407 267150 131416
rect 265716 127628 265768 127634
rect 265716 127570 265768 127576
rect 265806 127528 265862 127537
rect 265806 127463 265862 127472
rect 265714 122904 265770 122913
rect 265714 122839 265770 122848
rect 265728 94518 265756 122839
rect 265820 116657 265848 127463
rect 267002 118144 267058 118153
rect 267002 118079 267058 118088
rect 265806 116648 265862 116657
rect 265806 116583 265862 116592
rect 265806 114608 265862 114617
rect 265806 114543 265862 114552
rect 265716 94512 265768 94518
rect 265716 94454 265768 94460
rect 265820 90370 265848 114543
rect 265808 90364 265860 90370
rect 265808 90306 265860 90312
rect 265624 80708 265676 80714
rect 265624 80650 265676 80656
rect 264428 76628 264480 76634
rect 264428 76570 264480 76576
rect 264336 71052 264388 71058
rect 264336 70994 264388 71000
rect 267016 21418 267044 118079
rect 267108 62830 267136 131407
rect 267186 131064 267242 131073
rect 267186 130999 267242 131008
rect 267200 77994 267228 130999
rect 267292 115258 267320 138615
rect 280172 137057 280200 210394
rect 280344 177336 280396 177342
rect 280344 177278 280396 177284
rect 280252 176520 280304 176526
rect 280252 176462 280304 176468
rect 280264 156369 280292 176462
rect 280356 163985 280384 177278
rect 280816 176594 280844 276014
rect 282184 224256 282236 224262
rect 282184 224198 282236 224204
rect 282196 185638 282224 224198
rect 282184 185632 282236 185638
rect 282184 185574 282236 185580
rect 281540 181756 281592 181762
rect 281540 181698 281592 181704
rect 280804 176588 280856 176594
rect 280804 176530 280856 176536
rect 280436 176112 280488 176118
rect 280436 176054 280488 176060
rect 280448 170921 280476 176054
rect 280434 170912 280490 170921
rect 280434 170847 280490 170856
rect 280342 163976 280398 163985
rect 280342 163911 280398 163920
rect 281552 157049 281580 181698
rect 281632 176044 281684 176050
rect 281632 175986 281684 175992
rect 281538 157040 281594 157049
rect 281538 156975 281594 156984
rect 280250 156360 280306 156369
rect 280250 156295 280306 156304
rect 281644 152425 281672 175986
rect 281816 175976 281868 175982
rect 281816 175918 281868 175924
rect 281724 173596 281776 173602
rect 281724 173538 281776 173544
rect 281736 173233 281764 173538
rect 281722 173224 281778 173233
rect 281722 173159 281778 173168
rect 281724 170672 281776 170678
rect 281724 170614 281776 170620
rect 281736 170105 281764 170614
rect 281722 170096 281778 170105
rect 281722 170031 281778 170040
rect 281828 161474 281856 175918
rect 282644 172440 282696 172446
rect 282642 172408 282644 172417
rect 282696 172408 282698 172417
rect 282642 172343 282698 172352
rect 282734 169416 282790 169425
rect 282734 169351 282790 169360
rect 282748 168774 282776 169351
rect 282736 168768 282788 168774
rect 282736 168710 282788 168716
rect 282828 168700 282880 168706
rect 282828 168642 282880 168648
rect 282840 168609 282868 168642
rect 282826 168600 282882 168609
rect 282826 168535 282882 168544
rect 282736 168360 282788 168366
rect 282736 168302 282788 168308
rect 282748 167113 282776 168302
rect 282828 168292 282880 168298
rect 282828 168234 282880 168240
rect 282840 167793 282868 168234
rect 282826 167784 282882 167793
rect 282826 167719 282882 167728
rect 282734 167104 282790 167113
rect 282734 167039 282790 167048
rect 282000 165572 282052 165578
rect 282000 165514 282052 165520
rect 282012 164801 282040 165514
rect 282828 165504 282880 165510
rect 282826 165472 282828 165481
rect 282880 165472 282882 165481
rect 282826 165407 282882 165416
rect 281998 164792 282054 164801
rect 281998 164727 282054 164736
rect 282092 162852 282144 162858
rect 282092 162794 282144 162800
rect 282104 162489 282132 162794
rect 282090 162480 282146 162489
rect 282090 162415 282146 162424
rect 281736 161446 281856 161474
rect 281736 155553 281764 161446
rect 282460 161220 282512 161226
rect 282460 161162 282512 161168
rect 282472 160177 282500 161162
rect 282826 160848 282882 160857
rect 282932 160834 282960 283562
rect 283472 181484 283524 181490
rect 283472 181426 283524 181432
rect 283196 180192 283248 180198
rect 283196 180134 283248 180140
rect 283012 176656 283064 176662
rect 283010 176624 283012 176633
rect 283064 176624 283066 176633
rect 283010 176559 283066 176568
rect 283208 176474 283236 180134
rect 283380 178696 283432 178702
rect 283380 178638 283432 178644
rect 282882 160806 282960 160834
rect 283024 176446 283236 176474
rect 282826 160783 282882 160792
rect 282458 160168 282514 160177
rect 282458 160103 282514 160112
rect 282092 160064 282144 160070
rect 282092 160006 282144 160012
rect 282104 159361 282132 160006
rect 282090 159352 282146 159361
rect 282090 159287 282146 159296
rect 282828 158704 282880 158710
rect 282828 158646 282880 158652
rect 282840 158545 282868 158646
rect 282826 158536 282882 158545
rect 282826 158471 282882 158480
rect 281722 155544 281778 155553
rect 281722 155479 281778 155488
rect 281724 154556 281776 154562
rect 281724 154498 281776 154504
rect 281736 154057 281764 154498
rect 281722 154048 281778 154057
rect 281722 153983 281778 153992
rect 281630 152416 281686 152425
rect 281630 152351 281686 152360
rect 282828 151768 282880 151774
rect 282826 151736 282828 151745
rect 282880 151736 282882 151745
rect 282826 151671 282882 151680
rect 282644 151292 282696 151298
rect 282644 151234 282696 151240
rect 282656 150929 282684 151234
rect 282642 150920 282698 150929
rect 282642 150855 282698 150864
rect 282828 150408 282880 150414
rect 282828 150350 282880 150356
rect 282840 150113 282868 150350
rect 282826 150104 282882 150113
rect 282826 150039 282882 150048
rect 281724 149660 281776 149666
rect 281724 149602 281776 149608
rect 281736 149433 281764 149602
rect 281722 149424 281778 149433
rect 281722 149359 281778 149368
rect 282736 149048 282788 149054
rect 282736 148990 282788 148996
rect 282748 147801 282776 148990
rect 282828 148980 282880 148986
rect 282828 148922 282880 148928
rect 282840 148617 282868 148922
rect 282826 148608 282882 148617
rect 282826 148543 282882 148552
rect 282734 147792 282790 147801
rect 282734 147727 282790 147736
rect 282826 146296 282882 146305
rect 282000 146260 282052 146266
rect 282826 146231 282882 146240
rect 282000 146202 282052 146208
rect 282012 145489 282040 146202
rect 282840 146198 282868 146231
rect 282828 146192 282880 146198
rect 282828 146134 282880 146140
rect 281998 145480 282054 145489
rect 281998 145415 282054 145424
rect 282828 144900 282880 144906
rect 282828 144842 282880 144848
rect 282840 143993 282868 144842
rect 282826 143984 282882 143993
rect 282826 143919 282882 143928
rect 281632 143540 281684 143546
rect 281632 143482 281684 143488
rect 281644 142497 281672 143482
rect 281630 142488 281686 142497
rect 281630 142423 281686 142432
rect 282736 142112 282788 142118
rect 282736 142054 282788 142060
rect 282748 140865 282776 142054
rect 282828 142044 282880 142050
rect 282828 141986 282880 141992
rect 282840 141681 282868 141986
rect 282826 141672 282882 141681
rect 282826 141607 282882 141616
rect 282828 141432 282880 141438
rect 282828 141374 282880 141380
rect 282734 140856 282790 140865
rect 282734 140791 282790 140800
rect 281908 140752 281960 140758
rect 281908 140694 281960 140700
rect 281920 140185 281948 140694
rect 281906 140176 281962 140185
rect 281906 140111 281962 140120
rect 282840 139369 282868 141374
rect 282826 139360 282882 139369
rect 282826 139295 282882 139304
rect 282828 137964 282880 137970
rect 282828 137906 282880 137912
rect 282840 137873 282868 137906
rect 282826 137864 282882 137873
rect 282826 137799 282882 137808
rect 280158 137048 280214 137057
rect 280158 136983 280214 136992
rect 282368 136604 282420 136610
rect 282368 136546 282420 136552
rect 282380 135561 282408 136546
rect 282552 136400 282604 136406
rect 282550 136368 282552 136377
rect 282604 136368 282606 136377
rect 282550 136303 282606 136312
rect 282366 135552 282422 135561
rect 282366 135487 282422 135496
rect 283024 132494 283052 176446
rect 283392 176338 283420 178638
rect 283116 176310 283420 176338
rect 283116 133249 283144 176310
rect 283484 170678 283512 181426
rect 284312 173602 284340 283834
rect 285680 269136 285732 269142
rect 285680 269078 285732 269084
rect 284392 204944 284444 204950
rect 284392 204886 284444 204892
rect 284300 173596 284352 173602
rect 284300 173538 284352 173544
rect 283472 170672 283524 170678
rect 283472 170614 283524 170620
rect 283102 133240 283158 133249
rect 283102 133175 283158 133184
rect 282932 132466 283052 132494
rect 282736 132456 282788 132462
rect 282736 132398 282788 132404
rect 282826 132424 282882 132433
rect 282748 131753 282776 132398
rect 282826 132359 282828 132368
rect 282880 132359 282882 132368
rect 282828 132330 282880 132336
rect 282734 131744 282790 131753
rect 282734 131679 282790 131688
rect 282828 131096 282880 131102
rect 282828 131038 282880 131044
rect 282184 131028 282236 131034
rect 282184 130970 282236 130976
rect 282196 130121 282224 130970
rect 282840 130937 282868 131038
rect 282826 130928 282882 130937
rect 282826 130863 282882 130872
rect 282182 130112 282238 130121
rect 282182 130047 282238 130056
rect 282826 128616 282882 128625
rect 282932 128602 282960 132466
rect 282882 128574 282960 128602
rect 282826 128551 282882 128560
rect 281724 128308 281776 128314
rect 281724 128250 281776 128256
rect 281736 127809 281764 128250
rect 282828 128240 282880 128246
rect 282828 128182 282880 128188
rect 281722 127800 281778 127809
rect 281722 127735 281778 127744
rect 282840 127129 282868 128182
rect 282826 127120 282882 127129
rect 282826 127055 282882 127064
rect 281908 126948 281960 126954
rect 281908 126890 281960 126896
rect 281920 126313 281948 126890
rect 281906 126304 281962 126313
rect 281906 126239 281962 126248
rect 282828 125588 282880 125594
rect 282828 125530 282880 125536
rect 282736 125520 282788 125526
rect 282840 125497 282868 125530
rect 282736 125462 282788 125468
rect 282826 125488 282882 125497
rect 282748 124817 282776 125462
rect 282826 125423 282882 125432
rect 282734 124808 282790 124817
rect 282734 124743 282790 124752
rect 282644 124160 282696 124166
rect 282644 124102 282696 124108
rect 282656 123185 282684 124102
rect 282828 124092 282880 124098
rect 282828 124034 282880 124040
rect 282840 124001 282868 124034
rect 282826 123992 282882 124001
rect 282826 123927 282882 123936
rect 282736 123480 282788 123486
rect 282736 123422 282788 123428
rect 282642 123176 282698 123185
rect 282642 123111 282698 123120
rect 281540 121372 281592 121378
rect 281540 121314 281592 121320
rect 281552 120873 281580 121314
rect 281538 120864 281594 120873
rect 281538 120799 281594 120808
rect 282748 120193 282776 123422
rect 282828 122800 282880 122806
rect 282828 122742 282880 122748
rect 282840 121689 282868 122742
rect 282826 121680 282882 121689
rect 282826 121615 282882 121624
rect 284404 121378 284432 204886
rect 284484 185564 284536 185570
rect 284484 185506 284536 185512
rect 284392 121372 284444 121378
rect 284392 121314 284444 121320
rect 282734 120184 282790 120193
rect 282734 120119 282790 120128
rect 282092 120080 282144 120086
rect 282092 120022 282144 120028
rect 282104 119377 282132 120022
rect 282090 119368 282146 119377
rect 282090 119303 282146 119312
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282736 118584 282788 118590
rect 282840 118561 282868 118594
rect 282736 118526 282788 118532
rect 282826 118552 282882 118561
rect 282748 117881 282776 118526
rect 282826 118487 282882 118496
rect 282734 117872 282790 117881
rect 282734 117807 282790 117816
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282736 117224 282788 117230
rect 282736 117166 282788 117172
rect 282748 116385 282776 117166
rect 282840 117065 282868 117234
rect 282826 117056 282882 117065
rect 282826 116991 282882 117000
rect 282734 116376 282790 116385
rect 282734 116311 282790 116320
rect 281724 115932 281776 115938
rect 281724 115874 281776 115880
rect 267280 115252 267332 115258
rect 267280 115194 267332 115200
rect 281736 114753 281764 115874
rect 282092 115864 282144 115870
rect 282092 115806 282144 115812
rect 282104 115569 282132 115806
rect 282090 115560 282146 115569
rect 282090 115495 282146 115504
rect 281722 114744 281778 114753
rect 281722 114679 281778 114688
rect 282828 114504 282880 114510
rect 282828 114446 282880 114452
rect 282736 114436 282788 114442
rect 282736 114378 282788 114384
rect 267646 113384 267702 113393
rect 267646 113319 267702 113328
rect 267660 94518 267688 113319
rect 282748 113257 282776 114378
rect 282840 114073 282868 114446
rect 282826 114064 282882 114073
rect 282826 113999 282882 114008
rect 282734 113248 282790 113257
rect 282734 113183 282790 113192
rect 282092 113144 282144 113150
rect 282092 113086 282144 113092
rect 282104 112441 282132 113086
rect 282090 112432 282146 112441
rect 282090 112367 282146 112376
rect 282736 111784 282788 111790
rect 282736 111726 282788 111732
rect 282826 111752 282882 111761
rect 282748 110945 282776 111726
rect 282826 111687 282828 111696
rect 282880 111687 282882 111696
rect 282828 111658 282880 111664
rect 282734 110936 282790 110945
rect 282734 110871 282790 110880
rect 282092 110424 282144 110430
rect 282092 110366 282144 110372
rect 282104 110129 282132 110366
rect 282276 110356 282328 110362
rect 282276 110298 282328 110304
rect 282090 110120 282146 110129
rect 282090 110055 282146 110064
rect 282288 109449 282316 110298
rect 282274 109440 282330 109449
rect 282274 109375 282330 109384
rect 281724 108996 281776 109002
rect 281724 108938 281776 108944
rect 281736 107817 281764 108938
rect 282092 108928 282144 108934
rect 282092 108870 282144 108876
rect 282104 108633 282132 108870
rect 282090 108624 282146 108633
rect 282090 108559 282146 108568
rect 281722 107808 281778 107817
rect 281722 107743 281778 107752
rect 284496 106282 284524 185506
rect 284576 179036 284628 179042
rect 284576 178978 284628 178984
rect 284588 149666 284616 178978
rect 284576 149660 284628 149666
rect 284576 149602 284628 149608
rect 285692 126954 285720 269078
rect 287060 258188 287112 258194
rect 287060 258130 287112 258136
rect 285772 221468 285824 221474
rect 285772 221410 285824 221416
rect 285784 136406 285812 221410
rect 285864 188352 285916 188358
rect 285864 188294 285916 188300
rect 285876 151298 285904 188294
rect 285956 185632 286008 185638
rect 285956 185574 286008 185580
rect 285968 172446 285996 185574
rect 285956 172440 286008 172446
rect 285956 172382 286008 172388
rect 285864 151292 285916 151298
rect 285864 151234 285916 151240
rect 287072 148986 287100 258130
rect 288624 239488 288676 239494
rect 288624 239430 288676 239436
rect 288532 213240 288584 213246
rect 288532 213182 288584 213188
rect 287244 186992 287296 186998
rect 287244 186934 287296 186940
rect 287152 182844 287204 182850
rect 287152 182786 287204 182792
rect 287060 148980 287112 148986
rect 287060 148922 287112 148928
rect 285772 136400 285824 136406
rect 285772 136342 285824 136348
rect 285680 126948 285732 126954
rect 285680 126890 285732 126896
rect 281540 106276 281592 106282
rect 281540 106218 281592 106224
rect 284484 106276 284536 106282
rect 284484 106218 284536 106224
rect 281552 105505 281580 106218
rect 281538 105496 281594 105505
rect 281538 105431 281594 105440
rect 282828 104848 282880 104854
rect 282828 104790 282880 104796
rect 282840 104009 282868 104790
rect 282826 104000 282882 104009
rect 282826 103935 282882 103944
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282840 102513 282868 103430
rect 282826 102504 282882 102513
rect 282826 102439 282882 102448
rect 281814 101688 281870 101697
rect 281814 101623 281870 101632
rect 281538 100872 281594 100881
rect 281538 100807 281594 100816
rect 279330 98152 279386 98161
rect 279330 98087 279386 98096
rect 279344 96422 279372 98087
rect 279332 96416 279384 96422
rect 279332 96358 279384 96364
rect 279240 96348 279292 96354
rect 279240 96290 279292 96296
rect 279252 96121 279280 96290
rect 279238 96112 279294 96121
rect 267648 94512 267700 94518
rect 267648 94454 267700 94460
rect 269120 94512 269172 94518
rect 269120 94454 269172 94460
rect 270590 94480 270646 94489
rect 267188 77988 267240 77994
rect 267188 77930 267240 77936
rect 267096 62824 267148 62830
rect 267096 62766 267148 62772
rect 269132 47598 269160 94454
rect 270590 94415 270646 94424
rect 269120 47592 269172 47598
rect 269120 47534 269172 47540
rect 270604 28286 270632 94415
rect 270972 93702 271000 96084
rect 276952 93770 276980 96084
rect 279238 96047 279294 96056
rect 281552 95169 281580 100807
rect 281724 100700 281776 100706
rect 281724 100642 281776 100648
rect 281736 100201 281764 100642
rect 281722 100192 281778 100201
rect 281722 100127 281778 100136
rect 281538 95160 281594 95169
rect 281538 95095 281594 95104
rect 281828 93838 281856 101623
rect 282826 99376 282882 99385
rect 282826 99311 282828 99320
rect 282880 99311 282882 99320
rect 282828 99282 282880 99288
rect 282184 97980 282236 97986
rect 282184 97922 282236 97928
rect 282196 97073 282224 97922
rect 287164 97918 287192 182786
rect 287256 168706 287284 186934
rect 288440 177608 288492 177614
rect 288440 177550 288492 177556
rect 287336 176588 287388 176594
rect 287336 176530 287388 176536
rect 287244 168700 287296 168706
rect 287244 168642 287296 168648
rect 287348 161226 287376 176530
rect 288452 168298 288480 177550
rect 288440 168292 288492 168298
rect 288440 168234 288492 168240
rect 287336 161220 287388 161226
rect 287336 161162 287388 161168
rect 288544 117230 288572 213182
rect 288636 168774 288664 239430
rect 289820 234048 289872 234054
rect 289820 233990 289872 233996
rect 288716 229832 288768 229838
rect 288716 229774 288768 229780
rect 288624 168768 288676 168774
rect 288624 168710 288676 168716
rect 288728 118590 288756 229774
rect 289832 118658 289860 233990
rect 289912 203584 289964 203590
rect 289912 203526 289964 203532
rect 289924 128246 289952 203526
rect 290096 184204 290148 184210
rect 290096 184146 290148 184152
rect 290004 178968 290056 178974
rect 290004 178910 290056 178916
rect 290016 140758 290044 178910
rect 290108 150414 290136 184146
rect 290096 150408 290148 150414
rect 290096 150350 290148 150356
rect 291212 146198 291240 285738
rect 295340 273284 295392 273290
rect 295340 273226 295392 273232
rect 294052 258120 294104 258126
rect 294052 258062 294104 258068
rect 293960 234116 294012 234122
rect 293960 234058 294012 234064
rect 291292 228472 291344 228478
rect 291292 228414 291344 228420
rect 291200 146192 291252 146198
rect 291200 146134 291252 146140
rect 290004 140752 290056 140758
rect 290004 140694 290056 140700
rect 289912 128240 289964 128246
rect 289912 128182 289964 128188
rect 291304 120086 291332 228414
rect 292580 227044 292632 227050
rect 292580 226986 292632 226992
rect 291384 198008 291436 198014
rect 291384 197950 291436 197956
rect 291292 120080 291344 120086
rect 291292 120022 291344 120028
rect 289820 118652 289872 118658
rect 289820 118594 289872 118600
rect 288716 118584 288768 118590
rect 288716 118526 288768 118532
rect 288532 117224 288584 117230
rect 288532 117166 288584 117172
rect 291396 100706 291424 197950
rect 291476 185700 291528 185706
rect 291476 185642 291528 185648
rect 291488 141438 291516 185642
rect 291476 141432 291528 141438
rect 291476 141374 291528 141380
rect 292592 122806 292620 226986
rect 292764 192500 292816 192506
rect 292764 192442 292816 192448
rect 292672 180260 292724 180266
rect 292672 180202 292724 180208
rect 292580 122800 292632 122806
rect 292580 122742 292632 122748
rect 292684 110362 292712 180202
rect 292776 149054 292804 192442
rect 292856 180124 292908 180130
rect 292856 180066 292908 180072
rect 292868 160070 292896 180066
rect 292856 160064 292908 160070
rect 292856 160006 292908 160012
rect 292764 149048 292816 149054
rect 292764 148990 292816 148996
rect 292672 110356 292724 110362
rect 292672 110298 292724 110304
rect 293972 108934 294000 234058
rect 294064 158710 294092 258062
rect 294144 180328 294196 180334
rect 294144 180270 294196 180276
rect 294052 158704 294104 158710
rect 294052 158646 294104 158652
rect 293960 108928 294012 108934
rect 293960 108870 294012 108876
rect 291384 100700 291436 100706
rect 291384 100642 291436 100648
rect 294156 97986 294184 180270
rect 294236 177472 294288 177478
rect 294236 177414 294288 177420
rect 294248 144906 294276 177414
rect 294236 144900 294288 144906
rect 294236 144842 294288 144848
rect 295352 132394 295380 273226
rect 295432 235340 295484 235346
rect 295432 235282 295484 235288
rect 295340 132388 295392 132394
rect 295340 132330 295392 132336
rect 295444 128314 295472 235282
rect 296812 215960 296864 215966
rect 296812 215902 296864 215908
rect 296720 211812 296772 211818
rect 296720 211754 296772 211760
rect 295616 181620 295668 181626
rect 295616 181562 295668 181568
rect 295524 178832 295576 178838
rect 295524 178774 295576 178780
rect 295432 128308 295484 128314
rect 295432 128250 295484 128256
rect 295536 124098 295564 178774
rect 295628 162858 295656 181562
rect 295616 162852 295668 162858
rect 295616 162794 295668 162800
rect 295524 124092 295576 124098
rect 295524 124034 295576 124040
rect 296732 115870 296760 211754
rect 296824 165510 296852 215902
rect 296904 181688 296956 181694
rect 296904 181630 296956 181636
rect 296812 165504 296864 165510
rect 296812 165446 296864 165452
rect 296916 132462 296944 181630
rect 296996 178900 297048 178906
rect 296996 178842 297048 178848
rect 297008 143546 297036 178842
rect 296996 143540 297048 143546
rect 296996 143482 297048 143488
rect 296904 132456 296956 132462
rect 296904 132398 296956 132404
rect 296720 115864 296772 115870
rect 296720 115806 296772 115812
rect 298112 111722 298140 285767
rect 299480 284368 299532 284374
rect 299480 284310 299532 284316
rect 298190 244080 298246 244089
rect 298190 244015 298246 244024
rect 298204 125526 298232 244015
rect 298284 229764 298336 229770
rect 298284 229706 298336 229712
rect 298192 125520 298244 125526
rect 298192 125462 298244 125468
rect 298296 117298 298324 229706
rect 298376 182912 298428 182918
rect 298376 182854 298428 182860
rect 298388 142050 298416 182854
rect 298376 142044 298428 142050
rect 298376 141986 298428 141992
rect 298284 117292 298336 117298
rect 298284 117234 298336 117240
rect 298100 111716 298152 111722
rect 298100 111658 298152 111664
rect 299492 103494 299520 284310
rect 300124 271176 300176 271182
rect 300124 271118 300176 271124
rect 300136 238542 300164 271118
rect 300860 259480 300912 259486
rect 300860 259422 300912 259428
rect 300124 238536 300176 238542
rect 300124 238478 300176 238484
rect 299664 218748 299716 218754
rect 299664 218690 299716 218696
rect 299572 200796 299624 200802
rect 299572 200738 299624 200744
rect 299584 114442 299612 200738
rect 299676 165578 299704 218690
rect 299754 178664 299810 178673
rect 299754 178599 299810 178608
rect 299664 165572 299716 165578
rect 299664 165514 299716 165520
rect 299768 142118 299796 178599
rect 299756 142112 299808 142118
rect 299756 142054 299808 142060
rect 299572 114436 299624 114442
rect 299572 114378 299624 114384
rect 300872 113150 300900 259422
rect 300952 195288 301004 195294
rect 300952 195230 301004 195236
rect 300964 131034 300992 195230
rect 301044 177540 301096 177546
rect 301044 177482 301096 177488
rect 301056 168366 301084 177482
rect 301044 168360 301096 168366
rect 301044 168302 301096 168308
rect 300952 131028 301004 131034
rect 300952 130970 301004 130976
rect 300860 113144 300912 113150
rect 300860 113086 300912 113092
rect 302252 110430 302280 287030
rect 302332 227112 302384 227118
rect 302332 227054 302384 227060
rect 302344 114510 302372 227054
rect 302896 206990 302924 287234
rect 303620 285728 303672 285734
rect 303620 285670 303672 285676
rect 302884 206984 302936 206990
rect 302884 206926 302936 206932
rect 302424 189780 302476 189786
rect 302424 189722 302476 189728
rect 302436 146266 302464 189722
rect 302516 184272 302568 184278
rect 302516 184214 302568 184220
rect 302528 151774 302556 184214
rect 302516 151768 302568 151774
rect 302516 151710 302568 151716
rect 302424 146260 302476 146266
rect 302424 146202 302476 146208
rect 303632 123486 303660 285670
rect 304264 271924 304316 271930
rect 304264 271866 304316 271872
rect 304276 238610 304304 271866
rect 304264 238604 304316 238610
rect 304264 238546 304316 238552
rect 303712 232620 303764 232626
rect 303712 232562 303764 232568
rect 303620 123480 303672 123486
rect 303620 123422 303672 123428
rect 302332 114504 302384 114510
rect 302332 114446 302384 114452
rect 303724 111790 303752 232562
rect 303804 181552 303856 181558
rect 303804 181494 303856 181500
rect 303712 111784 303764 111790
rect 303712 111726 303764 111732
rect 302240 110424 302292 110430
rect 302240 110366 302292 110372
rect 303816 109002 303844 181494
rect 305012 136610 305040 292606
rect 305184 245676 305236 245682
rect 305184 245618 305236 245624
rect 305092 225616 305144 225622
rect 305092 225558 305144 225564
rect 305000 136604 305052 136610
rect 305000 136546 305052 136552
rect 303804 108996 303856 109002
rect 303804 108938 303856 108944
rect 305104 104854 305132 225558
rect 305196 125594 305224 245618
rect 305656 235958 305684 364346
rect 309140 287224 309192 287230
rect 309140 287166 309192 287172
rect 306380 252680 306432 252686
rect 306380 252622 306432 252628
rect 305644 235952 305696 235958
rect 305644 235894 305696 235900
rect 305184 125588 305236 125594
rect 305184 125530 305236 125536
rect 306392 124166 306420 252622
rect 306472 252612 306524 252618
rect 306472 252554 306524 252560
rect 306484 137970 306512 252554
rect 307760 249824 307812 249830
rect 307760 249766 307812 249772
rect 306472 137964 306524 137970
rect 306472 137906 306524 137912
rect 307772 131102 307800 249766
rect 307852 202156 307904 202162
rect 307852 202098 307904 202104
rect 307864 154562 307892 202098
rect 307852 154556 307904 154562
rect 307852 154498 307904 154504
rect 307760 131096 307812 131102
rect 307760 131038 307812 131044
rect 306380 124160 306432 124166
rect 306380 124102 306432 124108
rect 309152 115938 309180 287166
rect 309796 248334 309824 430578
rect 334624 287156 334676 287162
rect 334624 287098 334676 287104
rect 309784 248328 309836 248334
rect 309784 248270 309836 248276
rect 309230 224224 309286 224233
rect 309230 224159 309286 224168
rect 309140 115932 309192 115938
rect 309140 115874 309192 115880
rect 305092 104848 305144 104854
rect 305092 104790 305144 104796
rect 299480 103488 299532 103494
rect 299480 103430 299532 103436
rect 309244 99346 309272 224159
rect 334636 193186 334664 287098
rect 352562 285968 352618 285977
rect 352562 285903 352618 285912
rect 352576 224262 352604 285903
rect 363616 237386 363644 699654
rect 395356 239970 395384 700334
rect 397472 697610 397500 703520
rect 413664 700330 413692 703520
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 397460 697604 397512 697610
rect 397460 697546 397512 697552
rect 429212 293282 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700330 462360 703520
rect 453304 700324 453356 700330
rect 453304 700266 453356 700272
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 429200 293276 429252 293282
rect 429200 293218 429252 293224
rect 453316 240242 453344 700266
rect 478524 699718 478552 703520
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 497464 700324 497516 700330
rect 497464 700266 497516 700272
rect 475384 699712 475436 699718
rect 475384 699654 475436 699660
rect 478512 699712 478564 699718
rect 478512 699654 478564 699660
rect 475396 296002 475424 699654
rect 475384 295996 475436 296002
rect 475384 295938 475436 295944
rect 453304 240236 453356 240242
rect 453304 240178 453356 240184
rect 497476 240038 497504 700266
rect 527192 698970 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 698964 527232 698970
rect 527180 698906 527232 698912
rect 542372 246265 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 582378 697232 582434 697241
rect 582378 697167 582434 697176
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 566464 311908 566516 311914
rect 566464 311850 566516 311856
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 566476 266354 566504 311850
rect 580276 298790 580304 418231
rect 580264 298784 580316 298790
rect 580264 298726 580316 298732
rect 580354 298752 580410 298761
rect 580354 298687 580410 298696
rect 574744 289876 574796 289882
rect 574744 289818 574796 289824
rect 566464 266348 566516 266354
rect 566464 266290 566516 266296
rect 542358 246256 542414 246265
rect 542358 246191 542414 246200
rect 497464 240032 497516 240038
rect 497464 239974 497516 239980
rect 395344 239964 395396 239970
rect 395344 239906 395396 239912
rect 363604 237380 363656 237386
rect 363604 237322 363656 237328
rect 352564 224256 352616 224262
rect 352564 224198 352616 224204
rect 334624 193180 334676 193186
rect 334624 193122 334676 193128
rect 309232 99340 309284 99346
rect 309232 99282 309284 99288
rect 294144 97980 294196 97986
rect 294144 97922 294196 97928
rect 282828 97912 282880 97918
rect 282826 97880 282828 97889
rect 287152 97912 287204 97918
rect 282880 97880 282882 97889
rect 287152 97854 287204 97860
rect 282826 97815 282882 97824
rect 282182 97064 282238 97073
rect 282182 96999 282238 97008
rect 281816 93832 281868 93838
rect 281816 93774 281868 93780
rect 276940 93764 276992 93770
rect 276940 93706 276992 93712
rect 270960 93696 271012 93702
rect 270960 93638 271012 93644
rect 574756 73166 574784 289818
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 580368 271182 580396 298687
rect 582392 294642 582420 697167
rect 583022 683904 583078 683913
rect 583022 683839 583078 683848
rect 582654 670712 582710 670721
rect 582654 670647 582710 670656
rect 582470 644056 582526 644065
rect 582470 643991 582526 644000
rect 582380 294636 582432 294642
rect 582380 294578 582432 294584
rect 582378 284336 582434 284345
rect 582378 284271 582434 284280
rect 580356 271176 580408 271182
rect 580356 271118 580408 271124
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 579618 245576 579674 245585
rect 579618 245511 579674 245520
rect 579632 241534 579660 245511
rect 579620 241528 579672 241534
rect 579620 241470 579672 241476
rect 580264 224256 580316 224262
rect 580264 224198 580316 224204
rect 580276 219065 580304 224198
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 574744 73160 574796 73166
rect 574744 73102 574796 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 270592 28280 270644 28286
rect 270592 28222 270644 28228
rect 267004 21412 267056 21418
rect 267004 21354 267056 21360
rect 582392 19825 582420 284271
rect 582484 240174 582512 643991
rect 582562 630864 582618 630873
rect 582562 630799 582618 630808
rect 582472 240168 582524 240174
rect 582472 240110 582524 240116
rect 582576 240106 582604 630799
rect 582668 290465 582696 670647
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582654 290456 582710 290465
rect 582654 290391 582710 290400
rect 582760 254590 582788 617471
rect 582838 591016 582894 591025
rect 582838 590951 582894 590960
rect 582748 254584 582800 254590
rect 582748 254526 582800 254532
rect 582748 250504 582800 250510
rect 582748 250446 582800 250452
rect 582760 243574 582788 250446
rect 582748 243568 582800 243574
rect 582748 243510 582800 243516
rect 582564 240100 582616 240106
rect 582564 240042 582616 240048
rect 582852 237289 582880 590951
rect 582930 577688 582986 577697
rect 582930 577623 582986 577632
rect 582944 238678 582972 577623
rect 583036 356726 583064 683839
rect 583298 564360 583354 564369
rect 583298 564295 583354 564304
rect 583114 537840 583170 537849
rect 583114 537775 583170 537784
rect 583024 356720 583076 356726
rect 583024 356662 583076 356668
rect 583022 351928 583078 351937
rect 583022 351863 583078 351872
rect 583036 291854 583064 351863
rect 583024 291848 583076 291854
rect 583024 291790 583076 291796
rect 583024 288448 583076 288454
rect 583024 288390 583076 288396
rect 582932 238672 582984 238678
rect 582932 238614 582984 238620
rect 582838 237280 582894 237289
rect 582838 237215 582894 237224
rect 582656 236700 582708 236706
rect 582656 236642 582708 236648
rect 582472 235272 582524 235278
rect 582472 235214 582524 235220
rect 582378 19816 582434 19825
rect 582378 19751 582434 19760
rect 582484 6633 582512 235214
rect 582564 231124 582616 231130
rect 582564 231066 582616 231072
rect 582576 33153 582604 231066
rect 582668 46345 582696 236642
rect 582748 233912 582800 233918
rect 582748 233854 582800 233860
rect 582760 59673 582788 233854
rect 582840 209092 582892 209098
rect 582840 209034 582892 209040
rect 582852 86193 582880 209034
rect 583036 112849 583064 288390
rect 583128 238406 583156 537775
rect 583206 524512 583262 524521
rect 583206 524447 583262 524456
rect 583220 243545 583248 524447
rect 583312 300150 583340 564295
rect 583574 510776 583630 510785
rect 583574 510711 583630 510720
rect 583390 484664 583446 484673
rect 583390 484599 583446 484608
rect 583300 300144 583352 300150
rect 583300 300086 583352 300092
rect 583300 257372 583352 257378
rect 583300 257314 583352 257320
rect 583206 243536 583262 243545
rect 583206 243471 583262 243480
rect 583116 238400 583168 238406
rect 583116 238342 583168 238348
rect 583022 112840 583078 112849
rect 583022 112775 583078 112784
rect 583312 99521 583340 257314
rect 583404 256698 583432 484599
rect 583588 380186 583616 510711
rect 583850 471064 583906 471073
rect 583850 470999 583906 471008
rect 583576 380180 583628 380186
rect 583576 380122 583628 380128
rect 583574 378176 583630 378185
rect 583574 378111 583630 378120
rect 583588 282878 583616 378111
rect 583758 324728 583814 324737
rect 583758 324663 583814 324672
rect 583668 292596 583720 292602
rect 583668 292538 583720 292544
rect 583576 282872 583628 282878
rect 583576 282814 583628 282820
rect 583576 278792 583628 278798
rect 583576 278734 583628 278740
rect 583484 277432 583536 277438
rect 583484 277374 583536 277380
rect 583392 256692 583444 256698
rect 583392 256634 583444 256640
rect 583392 251252 583444 251258
rect 583392 251194 583444 251200
rect 583404 165889 583432 251194
rect 583390 165880 583446 165889
rect 583390 165815 583446 165824
rect 583496 161474 583524 277374
rect 583404 161446 583524 161474
rect 583404 152697 583432 161446
rect 583390 152688 583446 152697
rect 583390 152623 583446 152632
rect 583392 139392 583444 139398
rect 583390 139360 583392 139369
rect 583444 139360 583446 139369
rect 583390 139295 583446 139304
rect 583588 126585 583616 278734
rect 583680 179489 583708 292538
rect 583772 248402 583800 324663
rect 583864 276010 583892 470999
rect 583852 276004 583904 276010
rect 583852 275946 583904 275952
rect 583852 267776 583904 267782
rect 583852 267718 583904 267724
rect 583760 248396 583812 248402
rect 583760 248338 583812 248344
rect 583864 243642 583892 267718
rect 583852 243636 583904 243642
rect 583852 243578 583904 243584
rect 583760 243568 583812 243574
rect 583812 243516 583984 243522
rect 583760 243510 583984 243516
rect 583772 243494 583984 243510
rect 583852 243432 583904 243438
rect 583852 243374 583904 243380
rect 583864 232937 583892 243374
rect 583850 232928 583906 232937
rect 583850 232863 583906 232872
rect 583666 179480 583722 179489
rect 583666 179415 583722 179424
rect 583956 142154 583984 243494
rect 583864 142126 583984 142154
rect 583864 139398 583892 142126
rect 583852 139392 583904 139398
rect 583852 139334 583904 139340
rect 583574 126576 583630 126585
rect 583574 126511 583630 126520
rect 583298 99512 583354 99521
rect 583298 99447 583354 99456
rect 582838 86184 582894 86193
rect 582838 86119 582894 86128
rect 582746 59664 582802 59673
rect 582746 59599 582802 59608
rect 582654 46336 582710 46345
rect 582654 46271 582710 46280
rect 582562 33144 582618 33153
rect 582562 33079 582618 33088
rect 582470 6624 582526 6633
rect 582470 6559 582526 6568
rect 264244 2100 264296 2106
rect 264244 2042 264296 2048
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 619132 2834 619168
rect 2778 619112 2780 619132
rect 2780 619112 2832 619132
rect 2832 619112 2834 619132
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 2870 410488 2926 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3514 188808 3570 188864
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 3422 32408 3478 32464
rect 18 19896 74 19952
rect 3422 6432 3478 6488
rect 19246 66816 19302 66872
rect 16486 50224 16542 50280
rect 23386 65456 23442 65512
rect 22006 59880 22062 59936
rect 20626 21256 20682 21312
rect 28906 24112 28962 24168
rect 33046 57160 33102 57216
rect 31666 30912 31722 30968
rect 178682 238448 178738 238504
rect 102046 177520 102102 177576
rect 99470 176704 99526 176760
rect 105726 176704 105782 176760
rect 107014 176740 107016 176760
rect 107016 176740 107068 176760
rect 107068 176740 107070 176760
rect 107014 176704 107070 176740
rect 108118 176704 108174 176760
rect 109590 176704 109646 176760
rect 110694 176704 110750 176760
rect 112258 176704 112314 176760
rect 114466 176704 114522 176760
rect 121274 177248 121330 177304
rect 123298 177248 123354 177304
rect 130934 177520 130990 177576
rect 129462 177248 129518 177304
rect 116950 176704 117006 176760
rect 119526 176704 119582 176760
rect 125966 176704 126022 176760
rect 127162 176704 127218 176760
rect 128174 176704 128230 176760
rect 132406 176704 132462 176760
rect 134430 176704 134486 176760
rect 136086 176724 136142 176760
rect 136086 176704 136088 176724
rect 136088 176704 136140 176724
rect 136140 176704 136142 176724
rect 148230 176704 148286 176760
rect 158902 176704 158958 176760
rect 124494 175616 124550 175672
rect 133142 175616 133198 175672
rect 118422 175480 118478 175536
rect 121918 175480 121974 175536
rect 115754 174936 115810 174992
rect 166262 175344 166318 175400
rect 167642 176976 167698 177032
rect 167918 171536 167974 171592
rect 170402 176840 170458 176896
rect 171782 175480 171838 175536
rect 177302 178064 177358 178120
rect 66166 129240 66222 129296
rect 66074 128016 66130 128072
rect 65982 122576 66038 122632
rect 59266 94968 59322 95024
rect 62026 86808 62082 86864
rect 65890 120808 65946 120864
rect 65982 102312 66038 102368
rect 67454 126248 67510 126304
rect 66166 125160 66222 125216
rect 66074 93744 66130 93800
rect 67546 123528 67602 123584
rect 67454 91024 67510 91080
rect 67638 100680 67694 100736
rect 151634 94832 151690 94888
rect 109038 94696 109094 94752
rect 110694 94696 110750 94752
rect 115846 94696 115902 94752
rect 119434 94696 119490 94752
rect 100574 93472 100630 93528
rect 105542 93472 105598 93528
rect 118238 93472 118294 93528
rect 125414 93472 125470 93528
rect 151542 93492 151598 93528
rect 151542 93472 151544 93492
rect 151544 93472 151596 93492
rect 151596 93472 151598 93492
rect 110142 93200 110198 93256
rect 113822 93200 113878 93256
rect 74814 92384 74870 92440
rect 85854 92384 85910 92440
rect 91466 92384 91522 92440
rect 99010 92384 99066 92440
rect 104438 92384 104494 92440
rect 105726 92384 105782 92440
rect 106738 92384 106794 92440
rect 109590 92420 109592 92440
rect 109592 92420 109644 92440
rect 109644 92420 109646 92440
rect 109590 92384 109646 92420
rect 85026 91704 85082 91760
rect 91006 91840 91062 91896
rect 86774 91568 86830 91624
rect 85026 89528 85082 89584
rect 88062 91160 88118 91216
rect 89166 91160 89222 91216
rect 97354 91704 97410 91760
rect 93122 91160 93178 91216
rect 94410 91160 94466 91216
rect 95146 91160 95202 91216
rect 96342 91160 96398 91216
rect 91006 89664 91062 89720
rect 97814 91160 97870 91216
rect 98734 91160 98790 91216
rect 101862 91704 101918 91760
rect 99102 91160 99158 91216
rect 100206 91160 100262 91216
rect 101954 91296 102010 91352
rect 102046 91160 102102 91216
rect 102874 91160 102930 91216
rect 107566 91160 107622 91216
rect 107934 91160 107990 91216
rect 108946 91160 109002 91216
rect 57886 61376 57942 61432
rect 67546 43424 67602 43480
rect 113270 92404 113326 92440
rect 113270 92384 113272 92404
rect 113272 92384 113324 92404
rect 113324 92384 113326 92404
rect 111338 91160 111394 91216
rect 112074 91160 112130 91216
rect 112718 91160 112774 91216
rect 152094 93472 152150 93528
rect 115754 92384 115810 92440
rect 121182 92384 121238 92440
rect 123022 92384 123078 92440
rect 125782 92384 125838 92440
rect 136178 92384 136234 92440
rect 117134 91704 117190 91760
rect 114466 91160 114522 91216
rect 115018 91160 115074 91216
rect 119710 91160 119766 91216
rect 126610 91568 126666 91624
rect 121274 91160 121330 91216
rect 121918 91160 121974 91216
rect 122746 91160 122802 91216
rect 123298 91160 123354 91216
rect 124126 91160 124182 91216
rect 119986 84768 120042 84824
rect 123298 88168 123354 88224
rect 126886 91160 126942 91216
rect 128266 91160 128322 91216
rect 129646 91160 129702 91216
rect 131026 91160 131082 91216
rect 132406 91160 132462 91216
rect 133786 91160 133842 91216
rect 135166 91160 135222 91216
rect 151726 91160 151782 91216
rect 167826 111732 167828 111752
rect 167828 111732 167880 111752
rect 167880 111732 167882 111752
rect 167826 111696 167882 111732
rect 167826 110064 167882 110120
rect 167826 108704 167882 108760
rect 167734 93880 167790 93936
rect 169022 93608 169078 93664
rect 174634 92112 174690 92168
rect 177394 90888 177450 90944
rect 176014 89528 176070 89584
rect 121090 3304 121146 3360
rect 178774 177112 178830 177168
rect 184846 182824 184902 182880
rect 187514 189624 187570 189680
rect 186226 179968 186282 180024
rect 190366 186904 190422 186960
rect 190274 181464 190330 181520
rect 194414 190984 194470 191040
rect 193126 187040 193182 187096
rect 191746 177248 191802 177304
rect 198554 295296 198610 295352
rect 198554 282920 198610 282976
rect 197450 282376 197506 282432
rect 197358 281580 197414 281616
rect 197358 281560 197360 281580
rect 197360 281560 197412 281580
rect 197412 281560 197414 281580
rect 198646 280744 198702 280800
rect 197174 280200 197230 280256
rect 196990 260888 197046 260944
rect 197082 250824 197138 250880
rect 197358 279384 197414 279440
rect 198002 278568 198058 278624
rect 197358 278024 197414 278080
rect 197450 277208 197506 277264
rect 197266 276664 197322 276720
rect 195886 184184 195942 184240
rect 197358 275848 197414 275904
rect 197358 275032 197414 275088
rect 197450 274488 197506 274544
rect 197358 273672 197414 273728
rect 197450 272312 197506 272368
rect 197450 271496 197506 271552
rect 197358 270952 197414 271008
rect 197450 270136 197506 270192
rect 197358 269320 197414 269376
rect 197450 268776 197506 268832
rect 197358 267960 197414 268016
rect 197910 267144 197966 267200
rect 197358 266600 197414 266656
rect 197450 265784 197506 265840
rect 197358 264424 197414 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197450 262268 197506 262304
rect 197450 262248 197452 262268
rect 197452 262248 197504 262268
rect 197504 262248 197506 262268
rect 197358 261432 197414 261488
rect 197358 260072 197414 260128
rect 197450 259256 197506 259312
rect 197358 258712 197414 258768
rect 197358 257896 197414 257952
rect 197542 257352 197598 257408
rect 197358 256536 197414 256592
rect 197910 255720 197966 255776
rect 197450 255176 197506 255232
rect 197358 254360 197414 254416
rect 197358 253544 197414 253600
rect 198554 272856 198610 272912
rect 198094 265240 198150 265296
rect 198646 263064 198702 263120
rect 198554 259392 198610 259448
rect 198554 253000 198610 253056
rect 198370 251640 198426 251696
rect 197358 250008 197414 250064
rect 197450 249464 197506 249520
rect 197358 248648 197414 248704
rect 197634 247832 197690 247888
rect 197358 247288 197414 247344
rect 197358 245928 197414 245984
rect 197358 243752 197414 243808
rect 197450 242936 197506 242992
rect 197450 242120 197506 242176
rect 197358 241576 197414 241632
rect 198462 246472 198518 246528
rect 198370 225528 198426 225584
rect 198554 181328 198610 181384
rect 197266 178608 197322 178664
rect 199750 245112 199806 245168
rect 199106 241440 199162 241496
rect 199842 244296 199898 244352
rect 200946 284008 201002 284064
rect 201406 284144 201462 284200
rect 202234 288496 202290 288552
rect 207570 287136 207626 287192
rect 211986 285776 212042 285832
rect 218978 699760 219034 699816
rect 216586 291216 216642 291272
rect 217322 285640 217378 285696
rect 217046 284008 217102 284064
rect 219714 288632 219770 288688
rect 220634 286048 220690 286104
rect 220082 284280 220138 284336
rect 221186 285912 221242 285968
rect 223394 290400 223450 290456
rect 226982 290536 227038 290592
rect 228914 284416 228970 284472
rect 231582 284008 231638 284064
rect 233698 284280 233754 284336
rect 238482 286048 238538 286104
rect 243634 284008 243690 284064
rect 204902 283872 204958 283928
rect 210698 283872 210754 283928
rect 211710 283872 211766 283928
rect 217598 283872 217654 283928
rect 222658 283872 222714 283928
rect 224222 283872 224278 283928
rect 225234 283872 225290 283928
rect 226614 283872 226670 283928
rect 229466 283872 229522 283928
rect 231030 283872 231086 283928
rect 244002 279656 244058 279712
rect 244278 278840 244334 278896
rect 244278 260888 244334 260944
rect 244186 244160 244242 244216
rect 204718 240080 204774 240136
rect 204442 237360 204498 237416
rect 205546 240080 205602 240136
rect 180154 93744 180210 93800
rect 184386 89664 184442 89720
rect 189722 88168 189778 88224
rect 206742 185544 206798 185600
rect 206282 178064 206338 178120
rect 208858 238584 208914 238640
rect 211066 192480 211122 192536
rect 212446 178744 212502 178800
rect 213734 206216 213790 206272
rect 216586 208936 216642 208992
rect 219346 240080 219402 240136
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214010 171536 214066 171592
rect 213918 171028 213920 171048
rect 213920 171028 213972 171048
rect 213972 171028 213974 171048
rect 213918 170992 213974 171028
rect 214010 170312 214066 170368
rect 213918 169668 213920 169688
rect 213920 169668 213972 169688
rect 213972 169668 213974 169688
rect 213918 169632 213974 169668
rect 214010 168952 214066 169008
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 214010 167592 214066 167648
rect 213918 166912 213974 166968
rect 214102 166368 214158 166424
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 228178 238584 228234 238640
rect 227626 180104 227682 180160
rect 220910 175888 220966 175944
rect 229742 240080 229798 240136
rect 229098 177928 229154 177984
rect 228362 176024 228418 176080
rect 224222 175788 224224 175808
rect 224224 175788 224276 175808
rect 224276 175788 224278 175808
rect 224222 175752 224278 175788
rect 227626 175752 227682 175808
rect 229190 173712 229246 173768
rect 229098 173304 229154 173360
rect 214562 163648 214618 163704
rect 213918 162968 213974 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 158344 213974 158400
rect 214010 157664 214066 157720
rect 214930 157120 214986 157176
rect 213918 156440 213974 156496
rect 213918 155760 213974 155816
rect 229742 176704 229798 176760
rect 230478 174972 230480 174992
rect 230480 174972 230532 174992
rect 230532 174972 230534 174992
rect 230478 174936 230534 174972
rect 230478 165688 230534 165744
rect 230478 161608 230534 161664
rect 229282 158072 229338 158128
rect 229190 155760 229246 155816
rect 229098 155216 229154 155272
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 214010 153040 214066 153096
rect 213918 152496 213974 152552
rect 214470 151816 214526 151872
rect 215206 151136 215262 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 213918 149776 213974 149832
rect 214010 149096 214066 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 213918 143248 213974 143304
rect 214930 142568 214986 142624
rect 214010 141888 214066 141944
rect 213918 141208 213974 141264
rect 214010 140528 214066 140584
rect 213918 139848 213974 139904
rect 214010 139168 214066 139224
rect 214562 138624 214618 138680
rect 213918 137944 213974 138000
rect 214102 137264 214158 137320
rect 214010 136584 214066 136640
rect 213918 135260 213920 135280
rect 213920 135260 213972 135280
rect 213972 135260 213974 135280
rect 213918 135224 213974 135260
rect 213918 134544 213974 134600
rect 213366 133864 213422 133920
rect 214010 133320 214066 133376
rect 213918 132640 213974 132696
rect 213918 131280 213974 131336
rect 213918 130600 213974 130656
rect 214010 129920 214066 129976
rect 214010 129240 214066 129296
rect 213918 128696 213974 128752
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214102 119992 214158 120048
rect 214010 119448 214066 119504
rect 213918 118804 213920 118824
rect 213920 118804 213972 118824
rect 213972 118804 213974 118824
rect 213918 118768 213974 118804
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 213918 116728 213974 116784
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 213918 104916 213974 104952
rect 213918 104896 213920 104916
rect 213920 104896 213972 104916
rect 213972 104896 213974 104916
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 213458 102856 213514 102912
rect 214654 131960 214710 132016
rect 230478 158616 230534 158672
rect 230662 174256 230718 174312
rect 230570 157664 230626 157720
rect 229834 146240 229890 146296
rect 229742 136856 229798 136912
rect 216034 135904 216090 135960
rect 215022 105576 215078 105632
rect 214838 104216 214894 104272
rect 214562 102720 214618 102776
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 214746 101496 214802 101552
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 214010 96872 214066 96928
rect 214102 96328 214158 96384
rect 214562 88984 214618 89040
rect 215022 94968 215078 95024
rect 214838 91024 214894 91080
rect 214746 86808 214802 86864
rect 216218 116048 216274 116104
rect 229190 97144 229246 97200
rect 229098 97008 229154 97064
rect 229190 96600 229246 96656
rect 224222 93880 224278 93936
rect 222934 91704 222990 91760
rect 232962 238448 233018 238504
rect 231766 185680 231822 185736
rect 231766 175208 231822 175264
rect 231122 174664 231178 174720
rect 231582 172760 231638 172816
rect 231766 172388 231768 172408
rect 231768 172388 231820 172408
rect 231820 172388 231822 172408
rect 231766 172352 231822 172388
rect 231674 171808 231730 171864
rect 231490 171400 231546 171456
rect 231214 170448 231270 170504
rect 231766 170856 231822 170912
rect 231490 169904 231546 169960
rect 231674 169496 231730 169552
rect 231766 168952 231822 169008
rect 231122 168544 231178 168600
rect 231674 168036 231676 168056
rect 231676 168036 231728 168056
rect 231728 168036 231730 168056
rect 231674 168000 231730 168036
rect 231398 167592 231454 167648
rect 231766 167048 231822 167104
rect 231030 166676 231032 166696
rect 231032 166676 231084 166696
rect 231084 166676 231086 166696
rect 231030 166640 231086 166676
rect 230938 164736 230994 164792
rect 231306 166096 231362 166152
rect 231398 165144 231454 165200
rect 231306 164328 231362 164384
rect 231398 163784 231454 163840
rect 231122 162832 231178 162888
rect 231398 162424 231454 162480
rect 230938 161880 230994 161936
rect 231398 161472 231454 161528
rect 231398 160928 231454 160984
rect 230938 160520 230994 160576
rect 231398 160012 231400 160032
rect 231400 160012 231452 160032
rect 231452 160012 231454 160032
rect 231398 159976 231454 160012
rect 230938 159024 230994 159080
rect 231122 156712 231178 156768
rect 230938 154808 230994 154864
rect 231766 157120 231822 157176
rect 231766 154264 231822 154320
rect 231674 153720 231730 153776
rect 231490 153312 231546 153368
rect 231674 152904 231730 152960
rect 231766 152496 231822 152552
rect 231398 151952 231454 152008
rect 230754 149640 230810 149696
rect 230938 150048 230994 150104
rect 230846 149096 230902 149152
rect 230938 145560 230994 145616
rect 230938 142976 230994 143032
rect 231214 151580 231216 151600
rect 231216 151580 231268 151600
rect 231268 151580 231270 151600
rect 231214 151544 231270 151580
rect 231122 148144 231178 148200
rect 231766 148688 231822 148744
rect 231306 144336 231362 144392
rect 231306 142432 231362 142488
rect 231214 135904 231270 135960
rect 231030 134000 231086 134056
rect 231122 133048 231178 133104
rect 230846 127880 230902 127936
rect 230754 124108 230756 124128
rect 230756 124108 230808 124128
rect 230808 124108 230810 124128
rect 230754 124072 230810 124108
rect 230938 123528 230994 123584
rect 231122 125976 231178 126032
rect 230754 121624 230810 121680
rect 230938 119720 230994 119776
rect 230754 118904 230810 118960
rect 230662 116048 230718 116104
rect 229926 113192 229982 113248
rect 230570 110744 230626 110800
rect 230570 109384 230626 109440
rect 230846 107888 230902 107944
rect 230570 105168 230626 105224
rect 230846 104216 230902 104272
rect 231766 146784 231822 146840
rect 232042 150592 232098 150648
rect 231766 145832 231822 145888
rect 231674 144880 231730 144936
rect 231490 143928 231546 143984
rect 231766 141072 231822 141128
rect 231766 140684 231822 140720
rect 231766 140664 231768 140684
rect 231768 140664 231820 140684
rect 231820 140664 231822 140684
rect 231674 140120 231730 140176
rect 231766 138216 231822 138272
rect 231674 137844 231676 137864
rect 231676 137844 231728 137864
rect 231728 137844 231730 137864
rect 231674 137808 231730 137844
rect 231398 135360 231454 135416
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231766 133456 231822 133512
rect 231674 132504 231730 132560
rect 231766 132096 231822 132152
rect 231674 131552 231730 131608
rect 231306 131144 231362 131200
rect 231766 130600 231822 130656
rect 231674 130192 231730 130248
rect 231582 129784 231638 129840
rect 231490 124480 231546 124536
rect 231766 129240 231822 129296
rect 231674 128832 231730 128888
rect 231766 128288 231822 128344
rect 231766 126948 231822 126984
rect 231766 126928 231768 126948
rect 231768 126928 231820 126948
rect 231820 126928 231822 126948
rect 231674 126384 231730 126440
rect 231766 125468 231768 125488
rect 231768 125468 231820 125488
rect 231820 125468 231822 125488
rect 231766 125432 231822 125468
rect 231766 125060 231768 125080
rect 231768 125060 231820 125080
rect 231820 125060 231822 125080
rect 231766 125024 231822 125060
rect 231582 123120 231638 123176
rect 231766 122576 231822 122632
rect 231674 122168 231730 122224
rect 231582 120672 231638 120728
rect 231766 121216 231822 121272
rect 231674 120264 231730 120320
rect 231398 119312 231454 119368
rect 231214 116456 231270 116512
rect 231674 118396 231676 118416
rect 231676 118396 231728 118416
rect 231728 118396 231730 118416
rect 231674 118360 231730 118396
rect 231766 117952 231822 118008
rect 231490 117408 231546 117464
rect 231766 117000 231822 117056
rect 231766 115504 231822 115560
rect 231674 114552 231730 114608
rect 231766 114144 231822 114200
rect 231490 113600 231546 113656
rect 231766 112648 231822 112704
rect 231674 112240 231730 112296
rect 231306 111696 231362 111752
rect 231766 111288 231822 111344
rect 231766 110336 231822 110392
rect 231674 109792 231730 109848
rect 231766 108840 231822 108896
rect 231490 108432 231546 108488
rect 231306 107072 231362 107128
rect 231122 101768 231178 101824
rect 230754 100408 230810 100464
rect 231122 99864 231178 99920
rect 230662 98504 230718 98560
rect 231766 107516 231768 107536
rect 231768 107516 231820 107536
rect 231820 107516 231822 107536
rect 231766 107480 231822 107516
rect 231490 106528 231546 106584
rect 231766 106156 231768 106176
rect 231768 106156 231820 106176
rect 231820 106156 231822 106176
rect 231766 106120 231822 106156
rect 231674 105576 231730 105632
rect 231766 104660 231768 104680
rect 231768 104660 231820 104680
rect 231820 104660 231822 104680
rect 231766 104624 231822 104660
rect 231490 103672 231546 103728
rect 231766 103264 231822 103320
rect 231674 102720 231730 102776
rect 231582 102312 231638 102368
rect 231306 100816 231362 100872
rect 231582 99456 231638 99512
rect 231214 98912 231270 98968
rect 231122 97960 231178 98016
rect 231122 96192 231178 96248
rect 231766 101360 231822 101416
rect 231674 97552 231730 97608
rect 233422 177384 233478 177440
rect 234618 236000 234674 236056
rect 234710 175888 234766 175944
rect 234066 114416 234122 114472
rect 239770 240080 239826 240136
rect 238298 237360 238354 237416
rect 240598 240116 240600 240136
rect 240600 240116 240652 240136
rect 240652 240116 240654 240136
rect 240598 240080 240654 240116
rect 238850 182960 238906 183016
rect 240230 178608 240286 178664
rect 241518 176432 241574 176488
rect 241150 141344 241206 141400
rect 244186 234640 244242 234696
rect 241242 137264 241298 137320
rect 245750 290536 245806 290592
rect 245658 283736 245714 283792
rect 245934 282376 245990 282432
rect 246026 281560 246082 281616
rect 246026 281016 246082 281072
rect 245934 280220 245990 280256
rect 245934 280200 245936 280220
rect 245936 280200 245988 280220
rect 245988 280200 245990 280220
rect 245934 279384 245990 279440
rect 245934 278024 245990 278080
rect 245934 277480 245990 277536
rect 246026 276664 246082 276720
rect 245934 275848 245990 275904
rect 245934 275340 245936 275360
rect 245936 275340 245988 275360
rect 245988 275340 245990 275360
rect 245934 275304 245990 275340
rect 246026 274488 246082 274544
rect 245934 273672 245990 273728
rect 246026 273128 246082 273184
rect 245934 272312 245990 272368
rect 246026 271496 246082 271552
rect 245934 270952 245990 271008
rect 245934 269592 245990 269648
rect 246026 268776 246082 268832
rect 245934 267960 245990 268016
rect 246026 267416 246082 267472
rect 245842 265784 245898 265840
rect 245934 265240 245990 265296
rect 245934 264424 245990 264480
rect 245750 263880 245806 263936
rect 245658 263064 245714 263120
rect 244370 250824 244426 250880
rect 245934 262268 245990 262304
rect 245934 262248 245936 262268
rect 245936 262248 245988 262268
rect 245988 262248 245990 262268
rect 245842 261704 245898 261760
rect 245750 255992 245806 256048
rect 246118 260072 246174 260128
rect 245934 259528 245990 259584
rect 246026 258712 246082 258768
rect 245934 258168 245990 258224
rect 245934 257352 245990 257408
rect 245934 255176 245990 255232
rect 245842 254360 245898 254416
rect 245934 253816 245990 253872
rect 245842 253000 245898 253056
rect 245934 252184 245990 252240
rect 245934 251640 245990 251696
rect 245842 250280 245898 250336
rect 245934 249464 245990 249520
rect 245842 248104 245898 248160
rect 245934 247288 245990 247344
rect 245934 245928 245990 245984
rect 246026 245112 246082 245168
rect 245934 244568 245990 244624
rect 245842 243752 245898 243808
rect 245842 242392 245898 242448
rect 245750 241576 245806 241632
rect 245934 240760 245990 240816
rect 246394 266600 246450 266656
rect 246394 256536 246450 256592
rect 246302 242936 246358 242992
rect 246486 246472 246542 246528
rect 247130 270136 247186 270192
rect 257526 84768 257582 84824
rect 264242 182824 264298 182880
rect 265622 178608 265678 178664
rect 264334 177248 264390 177304
rect 271142 177384 271198 177440
rect 298098 285776 298154 285832
rect 278778 176024 278834 176080
rect 264978 175616 265034 175672
rect 265254 175208 265310 175264
rect 264978 174800 265034 174856
rect 265070 174392 265126 174448
rect 265162 173984 265218 174040
rect 264978 173576 265034 173632
rect 265070 173032 265126 173088
rect 264518 172624 264574 172680
rect 264242 162832 264298 162888
rect 264334 135224 264390 135280
rect 264242 118904 264298 118960
rect 264978 172216 265034 172272
rect 265070 171808 265126 171864
rect 264978 171400 265034 171456
rect 265070 170992 265126 171048
rect 264978 170040 265034 170096
rect 265162 170448 265218 170504
rect 265070 169632 265126 169688
rect 264978 169224 265034 169280
rect 265162 168816 265218 168872
rect 265254 168408 265310 168464
rect 265162 167864 265218 167920
rect 264978 167456 265034 167512
rect 265070 167048 265126 167104
rect 265162 166640 265218 166696
rect 265070 166232 265126 166288
rect 264978 165824 265034 165880
rect 264978 165280 265034 165336
rect 265070 164872 265126 164928
rect 265622 164464 265678 164520
rect 265162 164056 265218 164112
rect 265070 163648 265126 163704
rect 264978 163240 265034 163296
rect 265162 162288 265218 162344
rect 264978 161880 265034 161936
rect 265070 161472 265126 161528
rect 265070 161064 265126 161120
rect 264978 160248 265034 160304
rect 265162 160656 265218 160712
rect 265070 159704 265126 159760
rect 264978 159296 265034 159352
rect 265162 158908 265218 158944
rect 265162 158888 265164 158908
rect 265164 158888 265216 158908
rect 265216 158888 265218 158908
rect 265162 158480 265218 158536
rect 265070 158072 265126 158128
rect 264978 157664 265034 157720
rect 265162 157120 265218 157176
rect 265070 156712 265126 156768
rect 264978 156304 265034 156360
rect 265070 155896 265126 155952
rect 264978 155488 265034 155544
rect 279330 175208 279386 175264
rect 279330 162152 279386 162208
rect 279330 155216 279386 155272
rect 265162 155080 265218 155136
rect 265070 154128 265126 154184
rect 264978 153312 265034 153368
rect 265346 154536 265402 154592
rect 265162 153720 265218 153776
rect 265070 152904 265126 152960
rect 264978 151952 265034 152008
rect 265254 152496 265310 152552
rect 279422 153720 279478 153776
rect 264978 150728 265034 150784
rect 265070 150320 265126 150376
rect 264978 149504 265034 149560
rect 266082 151544 266138 151600
rect 265346 151136 265402 151192
rect 265070 148960 265126 149016
rect 264978 148144 265034 148200
rect 265162 148552 265218 148608
rect 265070 147328 265126 147384
rect 264978 146376 265034 146432
rect 265438 149912 265494 149968
rect 265806 147736 265862 147792
rect 265254 146920 265310 146976
rect 265162 145968 265218 146024
rect 265070 145560 265126 145616
rect 264978 145152 265034 145208
rect 265070 144744 265126 144800
rect 264978 144336 265034 144392
rect 265714 143792 265770 143848
rect 265162 143384 265218 143440
rect 264978 142976 265034 143032
rect 265070 142568 265126 142624
rect 265070 141752 265126 141808
rect 265162 141208 265218 141264
rect 264978 140800 265034 140856
rect 264978 139984 265034 140040
rect 265070 139168 265126 139224
rect 264978 138216 265034 138272
rect 265254 137808 265310 137864
rect 265070 137400 265126 137456
rect 264978 136992 265034 137048
rect 265162 136584 265218 136640
rect 265070 136176 265126 136232
rect 264978 135632 265034 135688
rect 265162 134816 265218 134872
rect 265070 134408 265126 134464
rect 264978 134020 265034 134056
rect 264978 134000 264980 134020
rect 264980 134000 265032 134020
rect 265032 134000 265034 134020
rect 264978 133592 265034 133648
rect 265070 133048 265126 133104
rect 265622 132640 265678 132696
rect 265070 130464 265126 130520
rect 264978 130056 265034 130112
rect 265070 129648 265126 129704
rect 264978 129240 265034 129296
rect 264978 127064 265034 127120
rect 265162 126656 265218 126712
rect 265070 126248 265126 126304
rect 264978 125840 265034 125896
rect 265162 125296 265218 125352
rect 265070 124888 265126 124944
rect 264978 124480 265034 124536
rect 265162 124072 265218 124128
rect 265070 123664 265126 123720
rect 264978 123256 265034 123312
rect 265070 122304 265126 122360
rect 265162 121896 265218 121952
rect 264978 121524 264980 121544
rect 264980 121524 265032 121544
rect 265032 121524 265034 121544
rect 264978 121488 265034 121524
rect 265162 121080 265218 121136
rect 264978 120672 265034 120728
rect 265070 120264 265126 120320
rect 264978 119720 265034 119776
rect 264978 118496 265034 118552
rect 265070 117680 265126 117736
rect 265162 117136 265218 117192
rect 264978 116728 265034 116784
rect 265070 116320 265126 116376
rect 264978 115912 265034 115968
rect 264978 115504 265034 115560
rect 265070 112920 265126 112976
rect 264978 112512 265034 112568
rect 265162 111988 265218 112024
rect 265162 111968 265164 111988
rect 265164 111968 265216 111988
rect 265216 111968 265218 111988
rect 265070 111560 265126 111616
rect 264978 110744 265034 110800
rect 265162 111152 265218 111208
rect 265070 110336 265126 110392
rect 264978 109928 265034 109984
rect 265162 109520 265218 109576
rect 265162 108976 265218 109032
rect 265070 108568 265126 108624
rect 264518 108160 264574 108216
rect 264426 106392 264482 106448
rect 264978 107788 264980 107808
rect 264980 107788 265032 107808
rect 265032 107788 265034 107808
rect 264978 107752 265034 107788
rect 265070 107344 265126 107400
rect 264978 106936 265034 106992
rect 265438 105984 265494 106040
rect 264978 105576 265034 105632
rect 265070 105168 265126 105224
rect 265162 104760 265218 104816
rect 265070 104352 265126 104408
rect 264978 103808 265034 103864
rect 265254 103400 265310 103456
rect 265070 102992 265126 103048
rect 265162 102584 265218 102640
rect 264978 102176 265034 102232
rect 265346 101768 265402 101824
rect 264978 101224 265034 101280
rect 265070 100852 265072 100872
rect 265072 100852 265124 100872
rect 265124 100852 265126 100872
rect 265070 100816 265126 100852
rect 265070 100000 265126 100056
rect 264978 99592 265034 99648
rect 265070 99184 265126 99240
rect 264978 98640 265034 98696
rect 264978 97824 265034 97880
rect 265162 97416 265218 97472
rect 265070 97008 265126 97064
rect 264978 96600 265034 96656
rect 264978 96192 265034 96248
rect 265898 142160 265954 142216
rect 267278 138624 267334 138680
rect 267094 131416 267150 131472
rect 265806 127472 265862 127528
rect 265714 122848 265770 122904
rect 267002 118088 267058 118144
rect 265806 116592 265862 116648
rect 265806 114552 265862 114608
rect 267186 131008 267242 131064
rect 280434 170856 280490 170912
rect 280342 163920 280398 163976
rect 281538 156984 281594 157040
rect 280250 156304 280306 156360
rect 281722 173168 281778 173224
rect 281722 170040 281778 170096
rect 282642 172388 282644 172408
rect 282644 172388 282696 172408
rect 282696 172388 282698 172408
rect 282642 172352 282698 172388
rect 282734 169360 282790 169416
rect 282826 168544 282882 168600
rect 282826 167728 282882 167784
rect 282734 167048 282790 167104
rect 282826 165452 282828 165472
rect 282828 165452 282880 165472
rect 282880 165452 282882 165472
rect 282826 165416 282882 165452
rect 281998 164736 282054 164792
rect 282090 162424 282146 162480
rect 282826 160792 282882 160848
rect 283010 176604 283012 176624
rect 283012 176604 283064 176624
rect 283064 176604 283066 176624
rect 283010 176568 283066 176604
rect 282458 160112 282514 160168
rect 282090 159296 282146 159352
rect 282826 158480 282882 158536
rect 281722 155488 281778 155544
rect 281722 153992 281778 154048
rect 281630 152360 281686 152416
rect 282826 151716 282828 151736
rect 282828 151716 282880 151736
rect 282880 151716 282882 151736
rect 282826 151680 282882 151716
rect 282642 150864 282698 150920
rect 282826 150048 282882 150104
rect 281722 149368 281778 149424
rect 282826 148552 282882 148608
rect 282734 147736 282790 147792
rect 282826 146240 282882 146296
rect 281998 145424 282054 145480
rect 282826 143928 282882 143984
rect 281630 142432 281686 142488
rect 282826 141616 282882 141672
rect 282734 140800 282790 140856
rect 281906 140120 281962 140176
rect 282826 139304 282882 139360
rect 282826 137808 282882 137864
rect 280158 136992 280214 137048
rect 282550 136348 282552 136368
rect 282552 136348 282604 136368
rect 282604 136348 282606 136368
rect 282550 136312 282606 136348
rect 282366 135496 282422 135552
rect 283102 133184 283158 133240
rect 282826 132388 282882 132424
rect 282826 132368 282828 132388
rect 282828 132368 282880 132388
rect 282880 132368 282882 132388
rect 282734 131688 282790 131744
rect 282826 130872 282882 130928
rect 282182 130056 282238 130112
rect 282826 128560 282882 128616
rect 281722 127744 281778 127800
rect 282826 127064 282882 127120
rect 281906 126248 281962 126304
rect 282826 125432 282882 125488
rect 282734 124752 282790 124808
rect 282826 123936 282882 123992
rect 282642 123120 282698 123176
rect 281538 120808 281594 120864
rect 282826 121624 282882 121680
rect 282734 120128 282790 120184
rect 282090 119312 282146 119368
rect 282826 118496 282882 118552
rect 282734 117816 282790 117872
rect 282826 117000 282882 117056
rect 282734 116320 282790 116376
rect 282090 115504 282146 115560
rect 281722 114688 281778 114744
rect 267646 113328 267702 113384
rect 282826 114008 282882 114064
rect 282734 113192 282790 113248
rect 282090 112376 282146 112432
rect 282826 111716 282882 111752
rect 282826 111696 282828 111716
rect 282828 111696 282880 111716
rect 282880 111696 282882 111716
rect 282734 110880 282790 110936
rect 282090 110064 282146 110120
rect 282274 109384 282330 109440
rect 282090 108568 282146 108624
rect 281722 107752 281778 107808
rect 281538 105440 281594 105496
rect 282826 103944 282882 104000
rect 282826 102448 282882 102504
rect 281814 101632 281870 101688
rect 281538 100816 281594 100872
rect 279330 98096 279386 98152
rect 270590 94424 270646 94480
rect 279238 96056 279294 96112
rect 281722 100136 281778 100192
rect 281538 95104 281594 95160
rect 282826 99340 282882 99376
rect 282826 99320 282828 99340
rect 282828 99320 282880 99340
rect 282880 99320 282882 99340
rect 298190 244024 298246 244080
rect 299754 178608 299810 178664
rect 309230 224168 309286 224224
rect 352562 285912 352618 285968
rect 582378 697176 582434 697232
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 579618 365064 579674 365120
rect 579986 312024 580042 312080
rect 580354 298696 580410 298752
rect 542358 246200 542414 246256
rect 282826 97860 282828 97880
rect 282828 97860 282880 97880
rect 282880 97860 282882 97880
rect 282826 97824 282882 97860
rect 282182 97008 282238 97064
rect 579802 272176 579858 272232
rect 583022 683848 583078 683904
rect 582654 670656 582710 670712
rect 582470 644000 582526 644056
rect 582378 284280 582434 284336
rect 580170 258848 580226 258904
rect 579618 245520 579674 245576
rect 580262 219000 580318 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 72936 580226 72992
rect 582562 630808 582618 630864
rect 582746 617480 582802 617536
rect 582654 290400 582710 290456
rect 582838 590960 582894 591016
rect 582930 577632 582986 577688
rect 583298 564304 583354 564360
rect 583114 537784 583170 537840
rect 583022 351872 583078 351928
rect 582838 237224 582894 237280
rect 582378 19760 582434 19816
rect 583206 524456 583262 524512
rect 583574 510720 583630 510776
rect 583390 484608 583446 484664
rect 583206 243480 583262 243536
rect 583022 112784 583078 112840
rect 583850 471008 583906 471064
rect 583574 378120 583630 378176
rect 583758 324672 583814 324728
rect 583390 165824 583446 165880
rect 583390 152632 583446 152688
rect 583390 139340 583392 139360
rect 583392 139340 583444 139360
rect 583444 139340 583446 139360
rect 583390 139304 583446 139340
rect 583850 232872 583906 232928
rect 583666 179424 583722 179480
rect 583574 126520 583630 126576
rect 583298 99456 583354 99512
rect 582838 86128 582894 86184
rect 582746 59608 582802 59664
rect 582654 46280 582710 46336
rect 582562 33088 582618 33144
rect 582470 6568 582526 6624
<< metal3 >>
rect 213126 699756 213132 699820
rect 213196 699818 213202 699820
rect 218973 699818 219039 699821
rect 213196 699816 219039 699818
rect 213196 699760 218978 699816
rect 219034 699760 219039 699816
rect 213196 699758 219039 699760
rect 213196 699756 213202 699758
rect 218973 699755 219039 699758
rect -960 697220 480 697460
rect 582373 697234 582439 697237
rect 583520 697234 584960 697324
rect 582373 697232 584960 697234
rect 582373 697176 582378 697232
rect 582434 697176 584960 697232
rect 582373 697174 584960 697176
rect 582373 697171 582439 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 583017 683906 583083 683909
rect 583520 683906 584960 683996
rect 583017 683904 584960 683906
rect 583017 683848 583022 683904
rect 583078 683848 584960 683904
rect 583017 683846 584960 683848
rect 583017 683843 583083 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582649 670714 582715 670717
rect 583520 670714 584960 670804
rect 582649 670712 584960 670714
rect 582649 670656 582654 670712
rect 582710 670656 584960 670712
rect 582649 670654 584960 670656
rect 582649 670651 582715 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582465 644058 582531 644061
rect 583520 644058 584960 644148
rect 582465 644056 584960 644058
rect 582465 644000 582470 644056
rect 582526 644000 584960 644056
rect 582465 643998 584960 644000
rect 582465 643995 582531 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 582557 630866 582623 630869
rect 583520 630866 584960 630956
rect 582557 630864 584960 630866
rect 582557 630808 582562 630864
rect 582618 630808 584960 630864
rect 582557 630806 584960 630808
rect 582557 630803 582623 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582833 591018 582899 591021
rect 583520 591018 584960 591108
rect 582833 591016 584960 591018
rect 582833 590960 582838 591016
rect 582894 590960 584960 591016
rect 582833 590958 584960 590960
rect 582833 590955 582899 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 582925 577690 582991 577693
rect 583520 577690 584960 577780
rect 582925 577688 584960 577690
rect 582925 577632 582930 577688
rect 582986 577632 584960 577688
rect 582925 577630 584960 577632
rect 582925 577627 582991 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 583293 564362 583359 564365
rect 583520 564362 584960 564452
rect 583293 564360 584960 564362
rect 583293 564304 583298 564360
rect 583354 564304 584960 564360
rect 583293 564302 584960 564304
rect 583293 564299 583359 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583109 537842 583175 537845
rect 583520 537842 584960 537932
rect 583109 537840 584960 537842
rect 583109 537784 583114 537840
rect 583170 537784 584960 537840
rect 583109 537782 584960 537784
rect 583109 537779 583175 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 583201 524514 583267 524517
rect 583520 524514 584960 524604
rect 583201 524512 584960 524514
rect 583201 524456 583206 524512
rect 583262 524456 584960 524512
rect 583201 524454 584960 524456
rect 583201 524451 583267 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 583520 511322 584960 511412
rect 583342 511262 584960 511322
rect 583342 511186 583402 511262
rect 583520 511186 584960 511262
rect 583342 511172 584960 511186
rect 583342 511126 583586 511172
rect 583526 510781 583586 511126
rect 583526 510776 583635 510781
rect 583526 510720 583574 510776
rect 583630 510720 583635 510776
rect 583526 510718 583635 510720
rect 583569 510715 583635 510718
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583385 484666 583451 484669
rect 583520 484666 584960 484756
rect 583385 484664 584960 484666
rect 583385 484608 583390 484664
rect 583446 484608 584960 484664
rect 583385 484606 584960 484608
rect 583385 484603 583451 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 583520 471474 584960 471564
rect 583342 471414 584960 471474
rect 583342 471338 583402 471414
rect 583520 471338 584960 471414
rect 583342 471324 584960 471338
rect 583342 471278 583770 471324
rect 583710 471066 583770 471278
rect 583845 471066 583911 471069
rect 583710 471064 583911 471066
rect 583710 471008 583850 471064
rect 583906 471008 583911 471064
rect 583710 471006 583911 471008
rect 583845 471003 583911 471006
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378450 584960 378540
rect 583342 378390 584960 378450
rect 583342 378314 583402 378390
rect 583520 378314 584960 378390
rect 583342 378300 584960 378314
rect 583342 378254 583586 378300
rect 583526 378181 583586 378254
rect 583526 378176 583635 378181
rect 583526 378120 583574 378176
rect 583630 378120 583635 378176
rect 583526 378118 583635 378120
rect 583569 378115 583635 378118
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 583017 351930 583083 351933
rect 583520 351930 584960 352020
rect 583017 351928 584960 351930
rect 583017 351872 583022 351928
rect 583078 351872 584960 351928
rect 583017 351870 584960 351872
rect 583017 351867 583083 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325274 584960 325364
rect 583342 325214 584960 325274
rect 583342 325138 583402 325214
rect 583520 325138 584960 325214
rect 583342 325124 584960 325138
rect 583342 325078 583770 325124
rect 583710 324733 583770 325078
rect 583710 324728 583819 324733
rect 583710 324672 583758 324728
rect 583814 324672 583819 324728
rect 583710 324670 583819 324672
rect 583753 324667 583819 324670
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 580349 298754 580415 298757
rect 583520 298754 584960 298844
rect 580349 298752 584960 298754
rect 580349 298696 580354 298752
rect 580410 298696 584960 298752
rect 580349 298694 584960 298696
rect 580349 298691 580415 298694
rect 583520 298604 584960 298694
rect 198549 295354 198615 295357
rect 285622 295354 285628 295356
rect 198549 295352 285628 295354
rect 198549 295296 198554 295352
rect 198610 295296 285628 295352
rect 198549 295294 285628 295296
rect 198549 295291 198615 295294
rect 285622 295292 285628 295294
rect 285692 295292 285698 295356
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 216581 291274 216647 291277
rect 248454 291274 248460 291276
rect 216581 291272 248460 291274
rect 216581 291216 216586 291272
rect 216642 291216 248460 291272
rect 216581 291214 248460 291216
rect 216581 291211 216647 291214
rect 248454 291212 248460 291214
rect 248524 291212 248530 291276
rect 226977 290594 227043 290597
rect 245745 290594 245811 290597
rect 226977 290592 245811 290594
rect 226977 290536 226982 290592
rect 227038 290536 245750 290592
rect 245806 290536 245811 290592
rect 226977 290534 245811 290536
rect 226977 290531 227043 290534
rect 245745 290531 245811 290534
rect 223389 290458 223455 290461
rect 582649 290458 582715 290461
rect 223389 290456 582715 290458
rect 223389 290400 223394 290456
rect 223450 290400 582654 290456
rect 582710 290400 582715 290456
rect 223389 290398 582715 290400
rect 223389 290395 223455 290398
rect 582649 290395 582715 290398
rect 219709 288690 219775 288693
rect 278814 288690 278820 288692
rect 219709 288688 278820 288690
rect 219709 288632 219714 288688
rect 219770 288632 278820 288688
rect 219709 288630 278820 288632
rect 219709 288627 219775 288630
rect 278814 288628 278820 288630
rect 278884 288628 278890 288692
rect 202229 288554 202295 288557
rect 288382 288554 288388 288556
rect 202229 288552 288388 288554
rect 202229 288496 202234 288552
rect 202290 288496 288388 288552
rect 202229 288494 288388 288496
rect 202229 288491 202295 288494
rect 288382 288492 288388 288494
rect 288452 288492 288458 288556
rect 207565 287194 207631 287197
rect 280286 287194 280292 287196
rect 207565 287192 280292 287194
rect 207565 287136 207570 287192
rect 207626 287136 280292 287192
rect 207565 287134 280292 287136
rect 207565 287131 207631 287134
rect 280286 287132 280292 287134
rect 280356 287132 280362 287196
rect 220629 286106 220695 286109
rect 228214 286106 228220 286108
rect 220629 286104 228220 286106
rect 220629 286048 220634 286104
rect 220690 286048 228220 286104
rect 220629 286046 228220 286048
rect 220629 286043 220695 286046
rect 228214 286044 228220 286046
rect 228284 286044 228290 286108
rect 238477 286106 238543 286109
rect 244406 286106 244412 286108
rect 238477 286104 244412 286106
rect 238477 286048 238482 286104
rect 238538 286048 244412 286104
rect 238477 286046 244412 286048
rect 238477 286043 238543 286046
rect 244406 286044 244412 286046
rect 244476 286044 244482 286108
rect 221181 285970 221247 285973
rect 352557 285970 352623 285973
rect 221181 285968 352623 285970
rect 221181 285912 221186 285968
rect 221242 285912 352562 285968
rect 352618 285912 352623 285968
rect 221181 285910 352623 285912
rect 221181 285907 221247 285910
rect 352557 285907 352623 285910
rect 211981 285834 212047 285837
rect 298093 285834 298159 285837
rect 211981 285832 298159 285834
rect 211981 285776 211986 285832
rect 212042 285776 298098 285832
rect 298154 285776 298159 285832
rect 211981 285774 298159 285776
rect 211981 285771 212047 285774
rect 298093 285771 298159 285774
rect 217317 285698 217383 285701
rect 220854 285698 220860 285700
rect 217317 285696 220860 285698
rect 217317 285640 217322 285696
rect 217378 285640 220860 285696
rect 217317 285638 220860 285640
rect 217317 285635 217383 285638
rect 220854 285636 220860 285638
rect 220924 285636 220930 285700
rect 583520 285276 584960 285516
rect 228909 284474 228975 284477
rect 287094 284474 287100 284476
rect 228909 284472 287100 284474
rect 228909 284416 228914 284472
rect 228970 284416 287100 284472
rect 228909 284414 287100 284416
rect 228909 284411 228975 284414
rect 287094 284412 287100 284414
rect 287164 284412 287170 284476
rect 220077 284338 220143 284341
rect 233182 284338 233188 284340
rect 220077 284336 233188 284338
rect 220077 284280 220082 284336
rect 220138 284280 233188 284336
rect 220077 284278 233188 284280
rect 220077 284275 220143 284278
rect 233182 284276 233188 284278
rect 233252 284276 233258 284340
rect 233693 284338 233759 284341
rect 582373 284338 582439 284341
rect 233693 284336 582439 284338
rect 233693 284280 233698 284336
rect 233754 284280 582378 284336
rect 582434 284280 582439 284336
rect 233693 284278 582439 284280
rect 233693 284275 233759 284278
rect 582373 284275 582439 284278
rect 201401 284202 201467 284205
rect 200806 284200 201467 284202
rect 200806 284144 201406 284200
rect 201462 284144 201467 284200
rect 200806 284142 201467 284144
rect 200806 283764 200866 284142
rect 201401 284139 201467 284142
rect 200941 284066 201007 284069
rect 201350 284066 201356 284068
rect 200941 284064 201356 284066
rect 200941 284008 200946 284064
rect 201002 284008 201356 284064
rect 200941 284006 201356 284008
rect 200941 284003 201007 284006
rect 201350 284004 201356 284006
rect 201420 284004 201426 284068
rect 217041 284066 217107 284069
rect 218094 284066 218100 284068
rect 217041 284064 218100 284066
rect 217041 284008 217046 284064
rect 217102 284008 218100 284064
rect 217041 284006 218100 284008
rect 217041 284003 217107 284006
rect 218094 284004 218100 284006
rect 218164 284004 218170 284068
rect 231577 284066 231643 284069
rect 231710 284066 231716 284068
rect 231577 284064 231716 284066
rect 231577 284008 231582 284064
rect 231638 284008 231716 284064
rect 231577 284006 231716 284008
rect 231577 284003 231643 284006
rect 231710 284004 231716 284006
rect 231780 284004 231786 284068
rect 243629 284066 243695 284069
rect 244222 284066 244228 284068
rect 243629 284064 244228 284066
rect 243629 284008 243634 284064
rect 243690 284008 244228 284064
rect 243629 284006 244228 284008
rect 243629 284003 243695 284006
rect 244222 284004 244228 284006
rect 244292 284004 244298 284068
rect 204897 283932 204963 283933
rect 204846 283930 204852 283932
rect 204806 283870 204852 283930
rect 204916 283928 204963 283932
rect 204958 283872 204963 283928
rect 204846 283868 204852 283870
rect 204916 283868 204963 283872
rect 204897 283867 204963 283868
rect 210693 283932 210759 283933
rect 210693 283928 210740 283932
rect 210804 283930 210810 283932
rect 211705 283930 211771 283933
rect 217593 283932 217659 283933
rect 212390 283930 212396 283932
rect 210693 283872 210698 283928
rect 210693 283868 210740 283872
rect 210804 283870 210850 283930
rect 211705 283928 212396 283930
rect 211705 283872 211710 283928
rect 211766 283872 212396 283928
rect 211705 283870 212396 283872
rect 210804 283868 210810 283870
rect 210693 283867 210759 283868
rect 211705 283867 211771 283870
rect 212390 283868 212396 283870
rect 212460 283868 212466 283932
rect 217542 283930 217548 283932
rect 217502 283870 217548 283930
rect 217612 283928 217659 283932
rect 217654 283872 217659 283928
rect 217542 283868 217548 283870
rect 217612 283868 217659 283872
rect 217593 283867 217659 283868
rect 222653 283930 222719 283933
rect 224217 283932 224283 283933
rect 223430 283930 223436 283932
rect 222653 283928 223436 283930
rect 222653 283872 222658 283928
rect 222714 283872 223436 283928
rect 222653 283870 223436 283872
rect 222653 283867 222719 283870
rect 223430 283868 223436 283870
rect 223500 283868 223506 283932
rect 224166 283930 224172 283932
rect 224126 283870 224172 283930
rect 224236 283928 224283 283932
rect 224278 283872 224283 283928
rect 224166 283868 224172 283870
rect 224236 283868 224283 283872
rect 224217 283867 224283 283868
rect 225229 283930 225295 283933
rect 226190 283930 226196 283932
rect 225229 283928 226196 283930
rect 225229 283872 225234 283928
rect 225290 283872 226196 283928
rect 225229 283870 226196 283872
rect 225229 283867 225295 283870
rect 226190 283868 226196 283870
rect 226260 283868 226266 283932
rect 226374 283868 226380 283932
rect 226444 283930 226450 283932
rect 226609 283930 226675 283933
rect 226444 283928 226675 283930
rect 226444 283872 226614 283928
rect 226670 283872 226675 283928
rect 226444 283870 226675 283872
rect 226444 283868 226450 283870
rect 226609 283867 226675 283870
rect 229461 283930 229527 283933
rect 229686 283930 229692 283932
rect 229461 283928 229692 283930
rect 229461 283872 229466 283928
rect 229522 283872 229692 283928
rect 229461 283870 229692 283872
rect 229461 283867 229527 283870
rect 229686 283868 229692 283870
rect 229756 283868 229762 283932
rect 231025 283930 231091 283933
rect 231526 283930 231532 283932
rect 231025 283928 231532 283930
rect 231025 283872 231030 283928
rect 231086 283872 231532 283928
rect 231025 283870 231532 283872
rect 231025 283867 231091 283870
rect 231526 283868 231532 283870
rect 231596 283868 231602 283932
rect 245653 283794 245719 283797
rect 244076 283792 245719 283794
rect 244076 283736 245658 283792
rect 245714 283736 245719 283792
rect 244076 283734 245719 283736
rect 245653 283731 245719 283734
rect 249742 283250 249748 283252
rect 244076 283190 249748 283250
rect 249742 283188 249748 283190
rect 249812 283188 249818 283252
rect 198549 282978 198615 282981
rect 198549 282976 200284 282978
rect 198549 282920 198554 282976
rect 198610 282920 200284 282976
rect 198549 282918 200284 282920
rect 198549 282915 198615 282918
rect 197445 282434 197511 282437
rect 245929 282434 245995 282437
rect 197445 282432 200284 282434
rect 197445 282376 197450 282432
rect 197506 282376 200284 282432
rect 197445 282374 200284 282376
rect 244076 282432 245995 282434
rect 244076 282376 245934 282432
rect 245990 282376 245995 282432
rect 244076 282374 245995 282376
rect 197445 282371 197511 282374
rect 245929 282371 245995 282374
rect 197353 281618 197419 281621
rect 246021 281618 246087 281621
rect 197353 281616 200284 281618
rect 197353 281560 197358 281616
rect 197414 281560 200284 281616
rect 197353 281558 200284 281560
rect 244076 281616 246087 281618
rect 244076 281560 246026 281616
rect 246082 281560 246087 281616
rect 244076 281558 246087 281560
rect 197353 281555 197419 281558
rect 246021 281555 246087 281558
rect 246021 281074 246087 281077
rect 244076 281072 246087 281074
rect 244076 281016 246026 281072
rect 246082 281016 246087 281072
rect 244076 281014 246087 281016
rect 246021 281011 246087 281014
rect 198641 280802 198707 280805
rect 198641 280800 200284 280802
rect 198641 280744 198646 280800
rect 198702 280744 200284 280800
rect 198641 280742 200284 280744
rect 198641 280739 198707 280742
rect 197169 280258 197235 280261
rect 245929 280258 245995 280261
rect 197169 280256 200284 280258
rect -960 279972 480 280212
rect 197169 280200 197174 280256
rect 197230 280200 200284 280256
rect 197169 280198 200284 280200
rect 244076 280256 245995 280258
rect 244076 280200 245934 280256
rect 245990 280200 245995 280256
rect 244076 280198 245995 280200
rect 197169 280195 197235 280198
rect 245929 280195 245995 280198
rect 243997 279714 244063 279717
rect 281574 279714 281580 279716
rect 243997 279712 281580 279714
rect 243997 279656 244002 279712
rect 244058 279656 281580 279712
rect 243997 279654 281580 279656
rect 243997 279651 244063 279654
rect 281574 279652 281580 279654
rect 281644 279652 281650 279716
rect 197353 279442 197419 279445
rect 245929 279442 245995 279445
rect 197353 279440 200284 279442
rect 197353 279384 197358 279440
rect 197414 279384 200284 279440
rect 197353 279382 200284 279384
rect 244076 279440 245995 279442
rect 244076 279384 245934 279440
rect 245990 279384 245995 279440
rect 244076 279382 245995 279384
rect 197353 279379 197419 279382
rect 245929 279379 245995 279382
rect 244273 278898 244339 278901
rect 244076 278896 244339 278898
rect 244076 278840 244278 278896
rect 244334 278840 244339 278896
rect 244076 278838 244339 278840
rect 244273 278835 244339 278838
rect 197997 278626 198063 278629
rect 197997 278624 200284 278626
rect 197997 278568 198002 278624
rect 198058 278568 200284 278624
rect 197997 278566 200284 278568
rect 197997 278563 198063 278566
rect 197353 278082 197419 278085
rect 245929 278082 245995 278085
rect 197353 278080 200284 278082
rect 197353 278024 197358 278080
rect 197414 278024 200284 278080
rect 197353 278022 200284 278024
rect 244076 278080 245995 278082
rect 244076 278024 245934 278080
rect 245990 278024 245995 278080
rect 244076 278022 245995 278024
rect 197353 278019 197419 278022
rect 245929 278019 245995 278022
rect 245929 277538 245995 277541
rect 244076 277536 245995 277538
rect 244076 277480 245934 277536
rect 245990 277480 245995 277536
rect 244076 277478 245995 277480
rect 245929 277475 245995 277478
rect 197445 277266 197511 277269
rect 197445 277264 200284 277266
rect 197445 277208 197450 277264
rect 197506 277208 200284 277264
rect 197445 277206 200284 277208
rect 197445 277203 197511 277206
rect 197261 276722 197327 276725
rect 246021 276722 246087 276725
rect 197261 276720 200284 276722
rect 197261 276664 197266 276720
rect 197322 276664 200284 276720
rect 197261 276662 200284 276664
rect 244076 276720 246087 276722
rect 244076 276664 246026 276720
rect 246082 276664 246087 276720
rect 244076 276662 246087 276664
rect 197261 276659 197327 276662
rect 246021 276659 246087 276662
rect 197353 275906 197419 275909
rect 245929 275906 245995 275909
rect 197353 275904 200284 275906
rect 197353 275848 197358 275904
rect 197414 275848 200284 275904
rect 197353 275846 200284 275848
rect 244076 275904 245995 275906
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 197353 275843 197419 275846
rect 245929 275843 245995 275846
rect 245929 275362 245995 275365
rect 244076 275360 245995 275362
rect 244076 275304 245934 275360
rect 245990 275304 245995 275360
rect 244076 275302 245995 275304
rect 245929 275299 245995 275302
rect 197353 275090 197419 275093
rect 197353 275088 200284 275090
rect 197353 275032 197358 275088
rect 197414 275032 200284 275088
rect 197353 275030 200284 275032
rect 197353 275027 197419 275030
rect 197445 274546 197511 274549
rect 246021 274546 246087 274549
rect 197445 274544 200284 274546
rect 197445 274488 197450 274544
rect 197506 274488 200284 274544
rect 197445 274486 200284 274488
rect 244076 274544 246087 274546
rect 244076 274488 246026 274544
rect 246082 274488 246087 274544
rect 244076 274486 246087 274488
rect 197445 274483 197511 274486
rect 246021 274483 246087 274486
rect 197353 273730 197419 273733
rect 245929 273730 245995 273733
rect 197353 273728 200284 273730
rect 197353 273672 197358 273728
rect 197414 273672 200284 273728
rect 197353 273670 200284 273672
rect 244076 273728 245995 273730
rect 244076 273672 245934 273728
rect 245990 273672 245995 273728
rect 244076 273670 245995 273672
rect 197353 273667 197419 273670
rect 245929 273667 245995 273670
rect 246021 273186 246087 273189
rect 244076 273184 246087 273186
rect 244076 273128 246026 273184
rect 246082 273128 246087 273184
rect 244076 273126 246087 273128
rect 246021 273123 246087 273126
rect 198549 272914 198615 272917
rect 198549 272912 200284 272914
rect 198549 272856 198554 272912
rect 198610 272856 200284 272912
rect 198549 272854 200284 272856
rect 198549 272851 198615 272854
rect 197445 272370 197511 272373
rect 245929 272370 245995 272373
rect 197445 272368 200284 272370
rect 197445 272312 197450 272368
rect 197506 272312 200284 272368
rect 197445 272310 200284 272312
rect 244076 272368 245995 272370
rect 244076 272312 245934 272368
rect 245990 272312 245995 272368
rect 244076 272310 245995 272312
rect 197445 272307 197511 272310
rect 245929 272307 245995 272310
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 197445 271554 197511 271557
rect 246021 271554 246087 271557
rect 197445 271552 200284 271554
rect 197445 271496 197450 271552
rect 197506 271496 200284 271552
rect 197445 271494 200284 271496
rect 244076 271552 246087 271554
rect 244076 271496 246026 271552
rect 246082 271496 246087 271552
rect 244076 271494 246087 271496
rect 197445 271491 197511 271494
rect 246021 271491 246087 271494
rect 197353 271010 197419 271013
rect 245929 271010 245995 271013
rect 197353 271008 200284 271010
rect 197353 270952 197358 271008
rect 197414 270952 200284 271008
rect 197353 270950 200284 270952
rect 244076 271008 245995 271010
rect 244076 270952 245934 271008
rect 245990 270952 245995 271008
rect 244076 270950 245995 270952
rect 197353 270947 197419 270950
rect 245929 270947 245995 270950
rect 197445 270194 197511 270197
rect 247125 270194 247191 270197
rect 197445 270192 200284 270194
rect 197445 270136 197450 270192
rect 197506 270136 200284 270192
rect 197445 270134 200284 270136
rect 244076 270192 247191 270194
rect 244076 270136 247130 270192
rect 247186 270136 247191 270192
rect 244076 270134 247191 270136
rect 197445 270131 197511 270134
rect 247125 270131 247191 270134
rect 245929 269650 245995 269653
rect 244076 269648 245995 269650
rect 244076 269592 245934 269648
rect 245990 269592 245995 269648
rect 244076 269590 245995 269592
rect 245929 269587 245995 269590
rect 197353 269378 197419 269381
rect 197353 269376 200284 269378
rect 197353 269320 197358 269376
rect 197414 269320 200284 269376
rect 197353 269318 200284 269320
rect 197353 269315 197419 269318
rect 197445 268834 197511 268837
rect 246021 268834 246087 268837
rect 197445 268832 200284 268834
rect 197445 268776 197450 268832
rect 197506 268776 200284 268832
rect 197445 268774 200284 268776
rect 244076 268832 246087 268834
rect 244076 268776 246026 268832
rect 246082 268776 246087 268832
rect 244076 268774 246087 268776
rect 197445 268771 197511 268774
rect 246021 268771 246087 268774
rect 197353 268018 197419 268021
rect 245929 268018 245995 268021
rect 197353 268016 200284 268018
rect 197353 267960 197358 268016
rect 197414 267960 200284 268016
rect 197353 267958 200284 267960
rect 244076 268016 245995 268018
rect 244076 267960 245934 268016
rect 245990 267960 245995 268016
rect 244076 267958 245995 267960
rect 197353 267955 197419 267958
rect 245929 267955 245995 267958
rect 246021 267474 246087 267477
rect 244076 267472 246087 267474
rect 244076 267416 246026 267472
rect 246082 267416 246087 267472
rect 244076 267414 246087 267416
rect 246021 267411 246087 267414
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 197905 267202 197971 267205
rect 197905 267200 200284 267202
rect 197905 267144 197910 267200
rect 197966 267144 200284 267200
rect 197905 267142 200284 267144
rect 197905 267139 197971 267142
rect 197353 266658 197419 266661
rect 246389 266658 246455 266661
rect 197353 266656 200284 266658
rect 197353 266600 197358 266656
rect 197414 266600 200284 266656
rect 197353 266598 200284 266600
rect 244076 266656 246455 266658
rect 244076 266600 246394 266656
rect 246450 266600 246455 266656
rect 244076 266598 246455 266600
rect 197353 266595 197419 266598
rect 246389 266595 246455 266598
rect 197445 265842 197511 265845
rect 245837 265842 245903 265845
rect 197445 265840 200284 265842
rect 197445 265784 197450 265840
rect 197506 265784 200284 265840
rect 197445 265782 200284 265784
rect 244076 265840 245903 265842
rect 244076 265784 245842 265840
rect 245898 265784 245903 265840
rect 244076 265782 245903 265784
rect 197445 265779 197511 265782
rect 245837 265779 245903 265782
rect 198089 265298 198155 265301
rect 245929 265298 245995 265301
rect 198089 265296 200284 265298
rect 198089 265240 198094 265296
rect 198150 265240 200284 265296
rect 198089 265238 200284 265240
rect 244076 265296 245995 265298
rect 244076 265240 245934 265296
rect 245990 265240 245995 265296
rect 244076 265238 245995 265240
rect 198089 265235 198155 265238
rect 245929 265235 245995 265238
rect 197353 264482 197419 264485
rect 245929 264482 245995 264485
rect 197353 264480 200284 264482
rect 197353 264424 197358 264480
rect 197414 264424 200284 264480
rect 197353 264422 200284 264424
rect 244076 264480 245995 264482
rect 244076 264424 245934 264480
rect 245990 264424 245995 264480
rect 244076 264422 245995 264424
rect 197353 264419 197419 264422
rect 245929 264419 245995 264422
rect 245745 263938 245811 263941
rect 244076 263936 245811 263938
rect 244076 263880 245750 263936
rect 245806 263880 245811 263936
rect 244076 263878 245811 263880
rect 245745 263875 245811 263878
rect 197353 263666 197419 263669
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 197353 263603 197419 263606
rect 198641 263122 198707 263125
rect 245653 263122 245719 263125
rect 198641 263120 200284 263122
rect 198641 263064 198646 263120
rect 198702 263064 200284 263120
rect 198641 263062 200284 263064
rect 244076 263120 245719 263122
rect 244076 263064 245658 263120
rect 245714 263064 245719 263120
rect 244076 263062 245719 263064
rect 198641 263059 198707 263062
rect 245653 263059 245719 263062
rect 197445 262306 197511 262309
rect 245929 262306 245995 262309
rect 197445 262304 200284 262306
rect 197445 262248 197450 262304
rect 197506 262248 200284 262304
rect 197445 262246 200284 262248
rect 244076 262304 245995 262306
rect 244076 262248 245934 262304
rect 245990 262248 245995 262304
rect 244076 262246 245995 262248
rect 197445 262243 197511 262246
rect 245929 262243 245995 262246
rect 245837 261762 245903 261765
rect 244076 261760 245903 261762
rect 244076 261704 245842 261760
rect 245898 261704 245903 261760
rect 244076 261702 245903 261704
rect 245837 261699 245903 261702
rect 197353 261490 197419 261493
rect 197353 261488 200284 261490
rect 197353 261432 197358 261488
rect 197414 261432 200284 261488
rect 197353 261430 200284 261432
rect 197353 261427 197419 261430
rect 196985 260946 197051 260949
rect 244273 260946 244339 260949
rect 196985 260944 200284 260946
rect 196985 260888 196990 260944
rect 197046 260888 200284 260944
rect 196985 260886 200284 260888
rect 244076 260944 244339 260946
rect 244076 260888 244278 260944
rect 244334 260888 244339 260944
rect 244076 260886 244339 260888
rect 196985 260883 197051 260886
rect 244273 260883 244339 260886
rect 197353 260130 197419 260133
rect 246113 260130 246179 260133
rect 197353 260128 200284 260130
rect 197353 260072 197358 260128
rect 197414 260072 200284 260128
rect 197353 260070 200284 260072
rect 244076 260128 246179 260130
rect 244076 260072 246118 260128
rect 246174 260072 246179 260128
rect 244076 260070 246179 260072
rect 197353 260067 197419 260070
rect 246113 260067 246179 260070
rect 245929 259586 245995 259589
rect 244076 259584 245995 259586
rect 244076 259528 245934 259584
rect 245990 259528 245995 259584
rect 244076 259526 245995 259528
rect 245929 259523 245995 259526
rect 198549 259450 198615 259453
rect 198774 259450 198780 259452
rect 198549 259448 198780 259450
rect 198549 259392 198554 259448
rect 198610 259392 198780 259448
rect 198549 259390 198780 259392
rect 198549 259387 198615 259390
rect 198774 259388 198780 259390
rect 198844 259388 198850 259452
rect 197445 259314 197511 259317
rect 197445 259312 200284 259314
rect 197445 259256 197450 259312
rect 197506 259256 200284 259312
rect 197445 259254 200284 259256
rect 197445 259251 197511 259254
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 197353 258770 197419 258773
rect 246021 258770 246087 258773
rect 197353 258768 200284 258770
rect 197353 258712 197358 258768
rect 197414 258712 200284 258768
rect 197353 258710 200284 258712
rect 244076 258768 246087 258770
rect 244076 258712 246026 258768
rect 246082 258712 246087 258768
rect 583520 258756 584960 258846
rect 244076 258710 246087 258712
rect 197353 258707 197419 258710
rect 246021 258707 246087 258710
rect 245929 258226 245995 258229
rect 244076 258224 245995 258226
rect 244076 258168 245934 258224
rect 245990 258168 245995 258224
rect 244076 258166 245995 258168
rect 245929 258163 245995 258166
rect 197353 257954 197419 257957
rect 197353 257952 200284 257954
rect 197353 257896 197358 257952
rect 197414 257896 200284 257952
rect 197353 257894 200284 257896
rect 197353 257891 197419 257894
rect 197537 257410 197603 257413
rect 245929 257410 245995 257413
rect 197537 257408 200284 257410
rect 197537 257352 197542 257408
rect 197598 257352 200284 257408
rect 197537 257350 200284 257352
rect 244076 257408 245995 257410
rect 244076 257352 245934 257408
rect 245990 257352 245995 257408
rect 244076 257350 245995 257352
rect 197537 257347 197603 257350
rect 245929 257347 245995 257350
rect 197353 256594 197419 256597
rect 246389 256594 246455 256597
rect 197353 256592 200284 256594
rect 197353 256536 197358 256592
rect 197414 256536 200284 256592
rect 197353 256534 200284 256536
rect 244076 256592 246455 256594
rect 244076 256536 246394 256592
rect 246450 256536 246455 256592
rect 244076 256534 246455 256536
rect 197353 256531 197419 256534
rect 246389 256531 246455 256534
rect 245745 256050 245811 256053
rect 244076 256048 245811 256050
rect 244076 255992 245750 256048
rect 245806 255992 245811 256048
rect 244076 255990 245811 255992
rect 245745 255987 245811 255990
rect 197905 255778 197971 255781
rect 197905 255776 200284 255778
rect 197905 255720 197910 255776
rect 197966 255720 200284 255776
rect 197905 255718 200284 255720
rect 197905 255715 197971 255718
rect 197445 255234 197511 255237
rect 245929 255234 245995 255237
rect 197445 255232 200284 255234
rect 197445 255176 197450 255232
rect 197506 255176 200284 255232
rect 197445 255174 200284 255176
rect 244076 255232 245995 255234
rect 244076 255176 245934 255232
rect 245990 255176 245995 255232
rect 244076 255174 245995 255176
rect 197445 255171 197511 255174
rect 245929 255171 245995 255174
rect 197353 254418 197419 254421
rect 245837 254418 245903 254421
rect 197353 254416 200284 254418
rect 197353 254360 197358 254416
rect 197414 254360 200284 254416
rect 197353 254358 200284 254360
rect 244076 254416 245903 254418
rect 244076 254360 245842 254416
rect 245898 254360 245903 254416
rect 244076 254358 245903 254360
rect 197353 254355 197419 254358
rect 245837 254355 245903 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 245929 253874 245995 253877
rect 244076 253872 245995 253874
rect 244076 253816 245934 253872
rect 245990 253816 245995 253872
rect 244076 253814 245995 253816
rect 245929 253811 245995 253814
rect 197353 253602 197419 253605
rect 197353 253600 200284 253602
rect 197353 253544 197358 253600
rect 197414 253544 200284 253600
rect 197353 253542 200284 253544
rect 197353 253539 197419 253542
rect 198549 253058 198615 253061
rect 245837 253058 245903 253061
rect 198549 253056 200284 253058
rect 198549 253000 198554 253056
rect 198610 253000 200284 253056
rect 198549 252998 200284 253000
rect 244076 253056 245903 253058
rect 244076 253000 245842 253056
rect 245898 253000 245903 253056
rect 244076 252998 245903 253000
rect 198549 252995 198615 252998
rect 245837 252995 245903 252998
rect 197118 252180 197124 252244
rect 197188 252242 197194 252244
rect 245929 252242 245995 252245
rect 197188 252182 200284 252242
rect 244076 252240 245995 252242
rect 244076 252184 245934 252240
rect 245990 252184 245995 252240
rect 244076 252182 245995 252184
rect 197188 252180 197194 252182
rect 245929 252179 245995 252182
rect 198365 251698 198431 251701
rect 245929 251698 245995 251701
rect 198365 251696 200284 251698
rect 198365 251640 198370 251696
rect 198426 251640 200284 251696
rect 198365 251638 200284 251640
rect 244076 251696 245995 251698
rect 244076 251640 245934 251696
rect 245990 251640 245995 251696
rect 244076 251638 245995 251640
rect 198365 251635 198431 251638
rect 245929 251635 245995 251638
rect 197077 250882 197143 250885
rect 244365 250882 244431 250885
rect 197077 250880 200284 250882
rect 197077 250824 197082 250880
rect 197138 250824 200284 250880
rect 197077 250822 200284 250824
rect 244076 250880 244431 250882
rect 244076 250824 244370 250880
rect 244426 250824 244431 250880
rect 244076 250822 244431 250824
rect 197077 250819 197143 250822
rect 244365 250819 244431 250822
rect 245837 250338 245903 250341
rect 244076 250336 245903 250338
rect 244076 250280 245842 250336
rect 245898 250280 245903 250336
rect 244076 250278 245903 250280
rect 245837 250275 245903 250278
rect 197353 250066 197419 250069
rect 197353 250064 200284 250066
rect 197353 250008 197358 250064
rect 197414 250008 200284 250064
rect 197353 250006 200284 250008
rect 197353 250003 197419 250006
rect 197445 249522 197511 249525
rect 245929 249522 245995 249525
rect 197445 249520 200284 249522
rect 197445 249464 197450 249520
rect 197506 249464 200284 249520
rect 197445 249462 200284 249464
rect 244076 249520 245995 249522
rect 244076 249464 245934 249520
rect 245990 249464 245995 249520
rect 244076 249462 245995 249464
rect 197445 249459 197511 249462
rect 245929 249459 245995 249462
rect 197353 248706 197419 248709
rect 248638 248706 248644 248708
rect 197353 248704 200284 248706
rect 197353 248648 197358 248704
rect 197414 248648 200284 248704
rect 197353 248646 200284 248648
rect 244076 248646 248644 248706
rect 197353 248643 197419 248646
rect 248638 248644 248644 248646
rect 248708 248644 248714 248708
rect 245837 248162 245903 248165
rect 244076 248160 245903 248162
rect 244076 248104 245842 248160
rect 245898 248104 245903 248160
rect 244076 248102 245903 248104
rect 245837 248099 245903 248102
rect 197629 247890 197695 247893
rect 197629 247888 200284 247890
rect 197629 247832 197634 247888
rect 197690 247832 200284 247888
rect 197629 247830 200284 247832
rect 197629 247827 197695 247830
rect 197353 247346 197419 247349
rect 245929 247346 245995 247349
rect 197353 247344 200284 247346
rect 197353 247288 197358 247344
rect 197414 247288 200284 247344
rect 197353 247286 200284 247288
rect 244076 247344 245995 247346
rect 244076 247288 245934 247344
rect 245990 247288 245995 247344
rect 244076 247286 245995 247288
rect 197353 247283 197419 247286
rect 245929 247283 245995 247286
rect 198457 246530 198523 246533
rect 246481 246530 246547 246533
rect 198457 246528 200284 246530
rect 198457 246472 198462 246528
rect 198518 246472 200284 246528
rect 198457 246470 200284 246472
rect 244076 246528 246547 246530
rect 244076 246472 246486 246528
rect 246542 246472 246547 246528
rect 244076 246470 246547 246472
rect 198457 246467 198523 246470
rect 246481 246467 246547 246470
rect 243486 246196 243492 246260
rect 243556 246258 243562 246260
rect 542353 246258 542419 246261
rect 243556 246256 542419 246258
rect 243556 246200 542358 246256
rect 542414 246200 542419 246256
rect 243556 246198 542419 246200
rect 243556 246196 243562 246198
rect 542353 246195 542419 246198
rect 197353 245986 197419 245989
rect 245929 245986 245995 245989
rect 197353 245984 200284 245986
rect 197353 245928 197358 245984
rect 197414 245928 200284 245984
rect 197353 245926 200284 245928
rect 244076 245984 245995 245986
rect 244076 245928 245934 245984
rect 245990 245928 245995 245984
rect 244076 245926 245995 245928
rect 197353 245923 197419 245926
rect 245929 245923 245995 245926
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 583520 245428 584960 245518
rect 199745 245170 199811 245173
rect 246021 245170 246087 245173
rect 199745 245168 200284 245170
rect 199745 245112 199750 245168
rect 199806 245112 200284 245168
rect 199745 245110 200284 245112
rect 244076 245168 246087 245170
rect 244076 245112 246026 245168
rect 246082 245112 246087 245168
rect 244076 245110 246087 245112
rect 199745 245107 199811 245110
rect 246021 245107 246087 245110
rect 245929 244626 245995 244629
rect 244076 244624 245995 244626
rect 244076 244568 245934 244624
rect 245990 244568 245995 244624
rect 244076 244566 245995 244568
rect 245929 244563 245995 244566
rect 199837 244354 199903 244357
rect 199837 244352 200284 244354
rect 199837 244296 199842 244352
rect 199898 244296 200284 244352
rect 199837 244294 200284 244296
rect 199837 244291 199903 244294
rect 244181 244220 244247 244221
rect 244181 244218 244228 244220
rect 244136 244216 244228 244218
rect 244136 244160 244186 244216
rect 244136 244158 244228 244160
rect 244181 244156 244228 244158
rect 244292 244156 244298 244220
rect 244181 244155 244247 244156
rect 244222 244020 244228 244084
rect 244292 244082 244298 244084
rect 298185 244082 298251 244085
rect 244292 244080 298251 244082
rect 244292 244024 298190 244080
rect 298246 244024 298251 244080
rect 244292 244022 298251 244024
rect 244292 244020 244298 244022
rect 298185 244019 298251 244022
rect 197353 243810 197419 243813
rect 245837 243810 245903 243813
rect 197353 243808 200284 243810
rect 197353 243752 197358 243808
rect 197414 243752 200284 243808
rect 197353 243750 200284 243752
rect 244076 243808 245903 243810
rect 244076 243752 245842 243808
rect 245898 243752 245903 243808
rect 244076 243750 245903 243752
rect 197353 243747 197419 243750
rect 245837 243747 245903 243750
rect 245878 243476 245884 243540
rect 245948 243538 245954 243540
rect 583201 243538 583267 243541
rect 245948 243536 583267 243538
rect 245948 243480 583206 243536
rect 583262 243480 583267 243536
rect 245948 243478 583267 243480
rect 245948 243476 245954 243478
rect 583201 243475 583267 243478
rect 197445 242994 197511 242997
rect 246297 242994 246363 242997
rect 197445 242992 200284 242994
rect 197445 242936 197450 242992
rect 197506 242936 200284 242992
rect 197445 242934 200284 242936
rect 244076 242992 246363 242994
rect 244076 242936 246302 242992
rect 246358 242936 246363 242992
rect 244076 242934 246363 242936
rect 197445 242931 197511 242934
rect 246297 242931 246363 242934
rect 245837 242450 245903 242453
rect 244076 242448 245903 242450
rect 244076 242392 245842 242448
rect 245898 242392 245903 242448
rect 244076 242390 245903 242392
rect 245837 242387 245903 242390
rect 197445 242178 197511 242181
rect 197445 242176 200284 242178
rect 197445 242120 197450 242176
rect 197506 242120 200284 242176
rect 197445 242118 200284 242120
rect 197445 242115 197511 242118
rect 197353 241634 197419 241637
rect 245745 241634 245811 241637
rect 197353 241632 200284 241634
rect 197353 241576 197358 241632
rect 197414 241576 200284 241632
rect 197353 241574 200284 241576
rect 244076 241632 245811 241634
rect 244076 241576 245750 241632
rect 245806 241576 245811 241632
rect 244076 241574 245811 241576
rect 197353 241571 197419 241574
rect 245745 241571 245811 241574
rect 198774 241436 198780 241500
rect 198844 241498 198850 241500
rect 199101 241498 199167 241501
rect 198844 241496 199167 241498
rect 198844 241440 199106 241496
rect 199162 241440 199167 241496
rect 198844 241438 199167 241440
rect 198844 241436 198850 241438
rect 199101 241435 199167 241438
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 245929 240818 245995 240821
rect 244076 240816 245995 240818
rect 200806 240138 200866 240788
rect 244076 240760 245934 240816
rect 245990 240760 245995 240816
rect 244076 240758 245995 240760
rect 245929 240755 245995 240758
rect 245878 240274 245884 240276
rect 244076 240214 245884 240274
rect 245878 240212 245884 240214
rect 245948 240212 245954 240276
rect 204713 240138 204779 240141
rect 200806 240136 204779 240138
rect 200806 240080 204718 240136
rect 204774 240080 204779 240136
rect 200806 240078 204779 240080
rect 204713 240075 204779 240078
rect 204846 240076 204852 240140
rect 204916 240138 204922 240140
rect 205541 240138 205607 240141
rect 204916 240136 205607 240138
rect 204916 240080 205546 240136
rect 205602 240080 205607 240136
rect 204916 240078 205607 240080
rect 204916 240076 204922 240078
rect 205541 240075 205607 240078
rect 218094 240076 218100 240140
rect 218164 240138 218170 240140
rect 219341 240138 219407 240141
rect 229737 240140 229803 240141
rect 229686 240138 229692 240140
rect 218164 240136 219407 240138
rect 218164 240080 219346 240136
rect 219402 240080 219407 240136
rect 218164 240078 219407 240080
rect 229646 240078 229692 240138
rect 229756 240136 229803 240140
rect 229798 240080 229803 240136
rect 218164 240076 218170 240078
rect 219341 240075 219407 240078
rect 229686 240076 229692 240078
rect 229756 240076 229803 240080
rect 229737 240075 229803 240076
rect 239765 240138 239831 240141
rect 240593 240138 240659 240141
rect 239765 240136 240659 240138
rect 239765 240080 239770 240136
rect 239826 240080 240598 240136
rect 240654 240080 240659 240136
rect 239765 240078 240659 240080
rect 239765 240075 239831 240078
rect 240593 240075 240659 240078
rect 208853 238642 208919 238645
rect 213126 238642 213132 238644
rect 208853 238640 213132 238642
rect 208853 238584 208858 238640
rect 208914 238584 213132 238640
rect 208853 238582 213132 238584
rect 208853 238579 208919 238582
rect 213126 238580 213132 238582
rect 213196 238580 213202 238644
rect 228173 238642 228239 238645
rect 243486 238642 243492 238644
rect 228173 238640 243492 238642
rect 228173 238584 228178 238640
rect 228234 238584 243492 238640
rect 228173 238582 243492 238584
rect 228173 238579 228239 238582
rect 243486 238580 243492 238582
rect 243556 238580 243562 238644
rect 178677 238506 178743 238509
rect 232957 238506 233023 238509
rect 178677 238504 233023 238506
rect 178677 238448 178682 238504
rect 178738 238448 232962 238504
rect 233018 238448 233023 238504
rect 178677 238446 233023 238448
rect 178677 238443 178743 238446
rect 232957 238443 233023 238446
rect 204437 237418 204503 237421
rect 204437 237416 204546 237418
rect 204437 237360 204442 237416
rect 204498 237360 204546 237416
rect 204437 237355 204546 237360
rect 237414 237356 237420 237420
rect 237484 237418 237490 237420
rect 238293 237418 238359 237421
rect 237484 237416 238359 237418
rect 237484 237360 238298 237416
rect 238354 237360 238359 237416
rect 237484 237358 238359 237360
rect 237484 237356 237490 237358
rect 238293 237355 238359 237358
rect 204486 237282 204546 237355
rect 582833 237282 582899 237285
rect 204486 237280 582899 237282
rect 204486 237224 582838 237280
rect 582894 237224 582899 237280
rect 204486 237222 582899 237224
rect 582833 237219 582899 237222
rect 231526 235996 231532 236060
rect 231596 236058 231602 236060
rect 234613 236058 234679 236061
rect 231596 236056 234679 236058
rect 231596 236000 234618 236056
rect 234674 236000 234679 236056
rect 231596 235998 234679 236000
rect 231596 235996 231602 235998
rect 234613 235995 234679 235998
rect 244181 234700 244247 234701
rect 244181 234698 244228 234700
rect 244136 234696 244228 234698
rect 244136 234640 244186 234696
rect 244136 234638 244228 234640
rect 244181 234636 244228 234638
rect 244292 234636 244298 234700
rect 244181 234635 244247 234636
rect 583845 232930 583911 232933
rect 583710 232928 583911 232930
rect 583710 232872 583850 232928
rect 583906 232872 583911 232928
rect 583710 232870 583911 232872
rect 583710 232522 583770 232870
rect 583845 232867 583911 232870
rect 583342 232476 583770 232522
rect 583342 232462 584960 232476
rect 583342 232386 583402 232462
rect 583520 232386 584960 232462
rect 583342 232326 584960 232386
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 198365 225586 198431 225589
rect 284334 225586 284340 225588
rect 198365 225584 284340 225586
rect 198365 225528 198370 225584
rect 198426 225528 284340 225584
rect 198365 225526 284340 225528
rect 198365 225523 198431 225526
rect 284334 225524 284340 225526
rect 284404 225524 284410 225588
rect 212390 224164 212396 224228
rect 212460 224226 212466 224228
rect 309225 224226 309291 224229
rect 212460 224224 309291 224226
rect 212460 224168 309230 224224
rect 309286 224168 309291 224224
rect 212460 224166 309291 224168
rect 212460 224164 212466 224166
rect 309225 224163 309291 224166
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 216581 208994 216647 208997
rect 231894 208994 231900 208996
rect 216581 208992 231900 208994
rect 216581 208936 216586 208992
rect 216642 208936 231900 208992
rect 216581 208934 231900 208936
rect 216581 208931 216647 208934
rect 231894 208932 231900 208934
rect 231964 208932 231970 208996
rect 213729 206274 213795 206277
rect 295374 206274 295380 206276
rect 213729 206272 295380 206274
rect 213729 206216 213734 206272
rect 213790 206216 295380 206272
rect 213729 206214 295380 206216
rect 213729 206211 213795 206214
rect 295374 206212 295380 206214
rect 295444 206212 295450 206276
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 231710 196012 231716 196076
rect 231780 196074 231786 196076
rect 236494 196074 236500 196076
rect 231780 196014 236500 196074
rect 231780 196012 231786 196014
rect 236494 196012 236500 196014
rect 236564 196012 236570 196076
rect 211061 192538 211127 192541
rect 287278 192538 287284 192540
rect 211061 192536 287284 192538
rect 211061 192480 211066 192536
rect 211122 192480 287284 192536
rect 211061 192478 287284 192480
rect 211061 192475 211127 192478
rect 287278 192476 287284 192478
rect 287348 192476 287354 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 194409 191042 194475 191045
rect 281758 191042 281764 191044
rect 194409 191040 281764 191042
rect 194409 190984 194414 191040
rect 194470 190984 281764 191040
rect 194409 190982 281764 190984
rect 194409 190979 194475 190982
rect 281758 190980 281764 190982
rect 281828 190980 281834 191044
rect 187509 189682 187575 189685
rect 274582 189682 274588 189684
rect 187509 189680 274588 189682
rect 187509 189624 187514 189680
rect 187570 189624 274588 189680
rect 187509 189622 274588 189624
rect 187509 189619 187575 189622
rect 274582 189620 274588 189622
rect 274652 189620 274658 189684
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 193121 187098 193187 187101
rect 229686 187098 229692 187100
rect 193121 187096 229692 187098
rect 193121 187040 193126 187096
rect 193182 187040 229692 187096
rect 193121 187038 229692 187040
rect 193121 187035 193187 187038
rect 229686 187036 229692 187038
rect 229756 187036 229762 187100
rect 190361 186962 190427 186965
rect 245694 186962 245700 186964
rect 190361 186960 245700 186962
rect 190361 186904 190366 186960
rect 190422 186904 245700 186960
rect 190361 186902 245700 186904
rect 190361 186899 190427 186902
rect 245694 186900 245700 186902
rect 245764 186900 245770 186964
rect 231761 185738 231827 185741
rect 232078 185738 232084 185740
rect 231761 185736 232084 185738
rect 231761 185680 231766 185736
rect 231822 185680 232084 185736
rect 231761 185678 232084 185680
rect 231761 185675 231827 185678
rect 232078 185676 232084 185678
rect 232148 185676 232154 185740
rect 206737 185602 206803 185605
rect 280286 185602 280292 185604
rect 206737 185600 280292 185602
rect 206737 185544 206742 185600
rect 206798 185544 280292 185600
rect 206737 185542 280292 185544
rect 206737 185539 206803 185542
rect 280286 185540 280292 185542
rect 280356 185540 280362 185604
rect 195881 184242 195947 184245
rect 234654 184242 234660 184244
rect 195881 184240 234660 184242
rect 195881 184184 195886 184240
rect 195942 184184 234660 184240
rect 195881 184182 234660 184184
rect 195881 184179 195947 184182
rect 234654 184180 234660 184182
rect 234724 184180 234730 184244
rect 210734 182956 210740 183020
rect 210804 183018 210810 183020
rect 238845 183018 238911 183021
rect 210804 183016 238911 183018
rect 210804 182960 238850 183016
rect 238906 182960 238911 183016
rect 210804 182958 238911 182960
rect 210804 182956 210810 182958
rect 238845 182955 238911 182958
rect 184841 182882 184907 182885
rect 230422 182882 230428 182884
rect 184841 182880 230428 182882
rect 184841 182824 184846 182880
rect 184902 182824 230428 182880
rect 184841 182822 230428 182824
rect 184841 182819 184907 182822
rect 230422 182820 230428 182822
rect 230492 182820 230498 182884
rect 264237 182882 264303 182885
rect 288566 182882 288572 182884
rect 264237 182880 288572 182882
rect 264237 182824 264242 182880
rect 264298 182824 288572 182880
rect 264237 182822 288572 182824
rect 264237 182819 264303 182822
rect 288566 182820 288572 182822
rect 288636 182820 288642 182884
rect 190269 181522 190335 181525
rect 237598 181522 237604 181524
rect 190269 181520 237604 181522
rect 190269 181464 190274 181520
rect 190330 181464 237604 181520
rect 190269 181462 237604 181464
rect 190269 181459 190335 181462
rect 237598 181460 237604 181462
rect 237668 181460 237674 181524
rect 198549 181386 198615 181389
rect 284518 181386 284524 181388
rect 198549 181384 284524 181386
rect 198549 181328 198554 181384
rect 198610 181328 284524 181384
rect 198549 181326 284524 181328
rect 198549 181323 198615 181326
rect 284518 181324 284524 181326
rect 284588 181324 284594 181388
rect 217542 180100 217548 180164
rect 217612 180162 217618 180164
rect 227621 180162 227687 180165
rect 217612 180160 227687 180162
rect 217612 180104 227626 180160
rect 227682 180104 227687 180160
rect 217612 180102 227687 180104
rect 217612 180100 217618 180102
rect 227621 180099 227687 180102
rect 186221 180026 186287 180029
rect 240358 180026 240364 180028
rect 186221 180024 240364 180026
rect 186221 179968 186226 180024
rect 186282 179968 240364 180024
rect 186221 179966 240364 179968
rect 186221 179963 186287 179966
rect 240358 179964 240364 179966
rect 240428 179964 240434 180028
rect 583661 179482 583727 179485
rect 583526 179480 583727 179482
rect 583526 179424 583666 179480
rect 583722 179424 583727 179480
rect 583526 179422 583727 179424
rect 583526 179346 583586 179422
rect 583661 179419 583727 179422
rect 583342 179300 583586 179346
rect 583342 179286 584960 179300
rect 583342 179210 583402 179286
rect 583520 179210 584960 179286
rect 583342 179150 584960 179210
rect 583520 179060 584960 179150
rect 212441 178802 212507 178805
rect 226374 178802 226380 178804
rect 212441 178800 226380 178802
rect 212441 178744 212446 178800
rect 212502 178744 226380 178800
rect 212441 178742 226380 178744
rect 212441 178739 212507 178742
rect 226374 178740 226380 178742
rect 226444 178740 226450 178804
rect 197261 178666 197327 178669
rect 240225 178666 240291 178669
rect 197261 178664 240291 178666
rect 197261 178608 197266 178664
rect 197322 178608 240230 178664
rect 240286 178608 240291 178664
rect 197261 178606 240291 178608
rect 197261 178603 197327 178606
rect 240225 178603 240291 178606
rect 265617 178666 265683 178669
rect 299749 178666 299815 178669
rect 265617 178664 299815 178666
rect 265617 178608 265622 178664
rect 265678 178608 299754 178664
rect 299810 178608 299815 178664
rect 265617 178606 299815 178608
rect 265617 178603 265683 178606
rect 299749 178603 299815 178606
rect 177297 178122 177363 178125
rect 97030 178120 177363 178122
rect 97030 178064 177302 178120
rect 177358 178064 177363 178120
rect 97030 178062 177363 178064
rect 97030 177988 97090 178062
rect 177297 178059 177363 178062
rect 201350 178060 201356 178124
rect 201420 178122 201426 178124
rect 206277 178122 206343 178125
rect 201420 178120 206343 178122
rect 201420 178064 206282 178120
rect 206338 178064 206343 178120
rect 201420 178062 206343 178064
rect 201420 178060 201426 178062
rect 206277 178059 206343 178062
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 226190 177924 226196 177988
rect 226260 177986 226266 177988
rect 229093 177986 229159 177989
rect 226260 177984 229159 177986
rect 226260 177928 229098 177984
rect 229154 177928 229159 177984
rect 226260 177926 229159 177928
rect 226260 177924 226266 177926
rect 229093 177923 229159 177926
rect 102041 177580 102107 177581
rect 101990 177578 101996 177580
rect 101950 177518 101996 177578
rect 102060 177576 102107 177580
rect 102102 177520 102107 177576
rect 101990 177516 101996 177518
rect 102060 177516 102107 177520
rect 130694 177516 130700 177580
rect 130764 177578 130770 177580
rect 130929 177578 130995 177581
rect 130764 177576 130995 177578
rect 130764 177520 130934 177576
rect 130990 177520 130995 177576
rect 130764 177518 130995 177520
rect 130764 177516 130770 177518
rect 102041 177515 102107 177516
rect 130929 177515 130995 177518
rect 228214 177380 228220 177444
rect 228284 177442 228290 177444
rect 233417 177442 233483 177445
rect 228284 177440 233483 177442
rect 228284 177384 233422 177440
rect 233478 177384 233483 177440
rect 228284 177382 233483 177384
rect 228284 177380 228290 177382
rect 233417 177379 233483 177382
rect 271137 177442 271203 177445
rect 285806 177442 285812 177444
rect 271137 177440 285812 177442
rect 271137 177384 271142 177440
rect 271198 177384 285812 177440
rect 271137 177382 285812 177384
rect 271137 177379 271203 177382
rect 285806 177380 285812 177382
rect 285876 177380 285882 177444
rect 120758 177244 120764 177308
rect 120828 177306 120834 177308
rect 121269 177306 121335 177309
rect 120828 177304 121335 177306
rect 120828 177248 121274 177304
rect 121330 177248 121335 177304
rect 120828 177246 121335 177248
rect 120828 177244 120834 177246
rect 121269 177243 121335 177246
rect 123150 177244 123156 177308
rect 123220 177306 123226 177308
rect 123293 177306 123359 177309
rect 129457 177308 129523 177309
rect 129406 177306 129412 177308
rect 123220 177304 123359 177306
rect 123220 177248 123298 177304
rect 123354 177248 123359 177304
rect 123220 177246 123359 177248
rect 129366 177246 129412 177306
rect 129476 177304 129523 177308
rect 129518 177248 129523 177304
rect 123220 177244 123226 177246
rect 123293 177243 123359 177246
rect 129406 177244 129412 177246
rect 129476 177244 129523 177248
rect 129457 177243 129523 177244
rect 191741 177306 191807 177309
rect 233366 177306 233372 177308
rect 191741 177304 233372 177306
rect 191741 177248 191746 177304
rect 191802 177248 233372 177304
rect 191741 177246 233372 177248
rect 191741 177243 191807 177246
rect 233366 177244 233372 177246
rect 233436 177244 233442 177308
rect 264329 177306 264395 177309
rect 291142 177306 291148 177308
rect 264329 177304 291148 177306
rect 264329 177248 264334 177304
rect 264390 177248 291148 177304
rect 264329 177246 291148 177248
rect 264329 177243 264395 177246
rect 291142 177244 291148 177246
rect 291212 177244 291218 177308
rect 100702 177108 100708 177172
rect 100772 177170 100778 177172
rect 178769 177170 178835 177173
rect 100772 177168 178835 177170
rect 100772 177112 178774 177168
rect 178830 177112 178835 177168
rect 100772 177110 178835 177112
rect 100772 177108 100778 177110
rect 178769 177107 178835 177110
rect 167637 177034 167703 177037
rect 103286 177032 167703 177034
rect 103286 176976 167642 177032
rect 167698 176976 167703 177032
rect 103286 176974 167703 176976
rect 99465 176762 99531 176765
rect 99422 176760 99531 176762
rect 99422 176704 99470 176760
rect 99526 176704 99531 176760
rect 99422 176699 99531 176704
rect 99422 176492 99482 176699
rect 103286 176492 103346 176974
rect 167637 176971 167703 176974
rect 104566 176836 104572 176900
rect 104636 176898 104642 176900
rect 170397 176898 170463 176901
rect 104636 176896 170463 176898
rect 104636 176840 170402 176896
rect 170458 176840 170463 176896
rect 104636 176838 170463 176840
rect 104636 176836 104642 176838
rect 170397 176835 170463 176838
rect 105721 176764 105787 176765
rect 107009 176764 107075 176765
rect 108113 176764 108179 176765
rect 109585 176764 109651 176765
rect 110689 176764 110755 176765
rect 105670 176762 105676 176764
rect 105630 176702 105676 176762
rect 105740 176760 105787 176764
rect 106958 176762 106964 176764
rect 105782 176704 105787 176760
rect 105670 176700 105676 176702
rect 105740 176700 105787 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 108062 176762 108068 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 109534 176762 109540 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109494 176702 109540 176762
rect 109604 176760 109651 176764
rect 110638 176762 110644 176764
rect 109646 176704 109651 176760
rect 109534 176700 109540 176702
rect 109604 176700 109651 176704
rect 110598 176702 110644 176762
rect 110708 176760 110755 176764
rect 110750 176704 110755 176760
rect 110638 176700 110644 176702
rect 110708 176700 110755 176704
rect 112110 176700 112116 176764
rect 112180 176762 112186 176764
rect 112253 176762 112319 176765
rect 112180 176760 112319 176762
rect 112180 176704 112258 176760
rect 112314 176704 112319 176760
rect 112180 176702 112319 176704
rect 112180 176700 112186 176702
rect 105721 176699 105787 176700
rect 107009 176699 107075 176700
rect 108113 176699 108179 176700
rect 109585 176699 109651 176700
rect 110689 176699 110755 176700
rect 112253 176699 112319 176702
rect 113214 176700 113220 176764
rect 113284 176762 113290 176764
rect 114461 176762 114527 176765
rect 116945 176764 117011 176765
rect 119521 176764 119587 176765
rect 116894 176762 116900 176764
rect 113284 176760 114527 176762
rect 113284 176704 114466 176760
rect 114522 176704 114527 176760
rect 113284 176702 114527 176704
rect 116854 176702 116900 176762
rect 116964 176760 117011 176764
rect 119470 176762 119476 176764
rect 117006 176704 117011 176760
rect 113284 176700 113290 176702
rect 114461 176699 114527 176702
rect 116894 176700 116900 176702
rect 116964 176700 117011 176704
rect 119430 176702 119476 176762
rect 119540 176760 119587 176764
rect 119582 176704 119587 176760
rect 119470 176700 119476 176702
rect 119540 176700 119587 176704
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 125961 176762 126027 176765
rect 125796 176760 126027 176762
rect 125796 176704 125966 176760
rect 126022 176704 126027 176760
rect 125796 176702 126027 176704
rect 125796 176700 125802 176702
rect 116945 176699 117011 176700
rect 119521 176699 119587 176700
rect 125961 176699 126027 176702
rect 127014 176700 127020 176764
rect 127084 176762 127090 176764
rect 127157 176762 127223 176765
rect 128169 176762 128235 176765
rect 132401 176764 132467 176765
rect 134425 176764 134491 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 158897 176764 158963 176765
rect 132350 176762 132356 176764
rect 127084 176760 127223 176762
rect 127084 176704 127162 176760
rect 127218 176704 127223 176760
rect 127084 176702 127223 176704
rect 127084 176700 127090 176702
rect 127157 176699 127223 176702
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 132310 176702 132356 176762
rect 132420 176760 132467 176764
rect 134374 176762 134380 176764
rect 132462 176704 132467 176760
rect 132350 176700 132356 176702
rect 132420 176700 132467 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 136030 176762 136036 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 158846 176762 158852 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158806 176702 158852 176762
rect 158916 176760 158963 176764
rect 158958 176704 158963 176760
rect 158846 176700 158852 176702
rect 158916 176700 158963 176704
rect 229134 176700 229140 176764
rect 229204 176762 229210 176764
rect 229737 176762 229803 176765
rect 229204 176760 229803 176762
rect 229204 176704 229742 176760
rect 229798 176704 229803 176760
rect 229204 176702 229803 176704
rect 229204 176700 229210 176702
rect 132401 176699 132467 176700
rect 134425 176699 134491 176700
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 158897 176699 158963 176700
rect 229737 176699 229803 176702
rect 128126 176492 128186 176699
rect 283005 176626 283071 176629
rect 283782 176626 283788 176628
rect 283005 176624 283788 176626
rect 283005 176568 283010 176624
rect 283066 176568 283788 176624
rect 283005 176566 283788 176568
rect 283005 176563 283071 176566
rect 283782 176564 283788 176566
rect 283852 176564 283858 176628
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 241513 176490 241579 176493
rect 241646 176490 241652 176492
rect 241513 176488 241652 176490
rect 241513 176432 241518 176488
rect 241574 176432 241652 176488
rect 241513 176430 241652 176432
rect 241513 176427 241579 176430
rect 241646 176428 241652 176430
rect 241716 176428 241722 176492
rect 228357 176082 228423 176085
rect 238518 176082 238524 176084
rect 228357 176080 238524 176082
rect -960 175796 480 176036
rect 228357 176024 228362 176080
rect 228418 176024 238524 176080
rect 228357 176022 238524 176024
rect 228357 176019 228423 176022
rect 238518 176020 238524 176022
rect 238588 176020 238594 176084
rect 278773 176082 278839 176085
rect 278773 176080 279434 176082
rect 278773 176024 278778 176080
rect 278834 176024 279434 176080
rect 278773 176022 279434 176024
rect 278773 176019 278839 176022
rect 220905 175948 220971 175949
rect 220854 175946 220860 175948
rect 220814 175886 220860 175946
rect 220924 175944 220971 175948
rect 220966 175888 220971 175944
rect 220854 175884 220860 175886
rect 220924 175884 220971 175888
rect 223430 175884 223436 175948
rect 223500 175946 223506 175948
rect 234705 175946 234771 175949
rect 223500 175944 234771 175946
rect 223500 175888 234710 175944
rect 234766 175888 234771 175944
rect 223500 175886 234771 175888
rect 223500 175884 223506 175886
rect 220905 175883 220971 175884
rect 234705 175883 234771 175886
rect 224217 175812 224283 175813
rect 224166 175810 224172 175812
rect 224126 175750 224172 175810
rect 224236 175808 224283 175812
rect 224278 175752 224283 175808
rect 224166 175748 224172 175750
rect 224236 175748 224283 175752
rect 224217 175747 224283 175748
rect 227621 175810 227687 175813
rect 227621 175808 228282 175810
rect 227621 175752 227626 175808
rect 227682 175752 228282 175808
rect 227621 175750 228282 175752
rect 227621 175747 227687 175750
rect 124489 175676 124555 175677
rect 133137 175676 133203 175677
rect 114318 175612 114324 175676
rect 114388 175674 114394 175676
rect 124438 175674 124444 175676
rect 114388 175614 122850 175674
rect 124398 175614 124444 175674
rect 124508 175672 124555 175676
rect 133086 175674 133092 175676
rect 124550 175616 124555 175672
rect 114388 175612 114394 175614
rect 118417 175540 118483 175541
rect 121913 175540 121979 175541
rect 118366 175538 118372 175540
rect 118326 175478 118372 175538
rect 118436 175536 118483 175540
rect 121862 175538 121868 175540
rect 118478 175480 118483 175536
rect 118366 175476 118372 175478
rect 118436 175476 118483 175480
rect 121822 175478 121868 175538
rect 121932 175536 121979 175540
rect 121974 175480 121979 175536
rect 121862 175476 121868 175478
rect 121932 175476 121979 175480
rect 122790 175538 122850 175614
rect 124438 175612 124444 175614
rect 124508 175612 124555 175616
rect 133046 175614 133092 175674
rect 133156 175672 133203 175676
rect 133198 175616 133203 175672
rect 133086 175612 133092 175614
rect 133156 175612 133203 175616
rect 124489 175611 124555 175612
rect 133137 175611 133203 175612
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 228222 175644 228282 175750
rect 274582 175748 274588 175812
rect 274652 175810 274658 175812
rect 279182 175810 279188 175812
rect 274652 175750 279188 175810
rect 274652 175748 274658 175750
rect 279182 175748 279188 175750
rect 279252 175748 279258 175812
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 213913 175614 217212 175616
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 213913 175611 213979 175614
rect 264973 175611 265039 175614
rect 171777 175538 171843 175541
rect 122790 175536 171843 175538
rect 122790 175480 171782 175536
rect 171838 175480 171843 175536
rect 279374 175508 279434 176022
rect 122790 175478 171843 175480
rect 118417 175475 118483 175476
rect 121913 175475 121979 175476
rect 171777 175475 171843 175478
rect 98310 175340 98316 175404
rect 98380 175402 98386 175404
rect 166257 175402 166323 175405
rect 98380 175400 166323 175402
rect 98380 175344 166262 175400
rect 166318 175344 166323 175400
rect 98380 175342 166323 175344
rect 98380 175340 98386 175342
rect 166257 175339 166323 175342
rect 231761 175266 231827 175269
rect 228804 175264 231827 175266
rect 228804 175208 231766 175264
rect 231822 175208 231827 175264
rect 228804 175206 231827 175208
rect 231761 175203 231827 175206
rect 265249 175266 265315 175269
rect 279325 175266 279391 175269
rect 265249 175264 268180 175266
rect 265249 175208 265254 175264
rect 265310 175208 268180 175264
rect 265249 175206 268180 175208
rect 279325 175264 279434 175266
rect 279325 175208 279330 175264
rect 279386 175208 279434 175264
rect 265249 175203 265315 175206
rect 279325 175203 279434 175208
rect 115749 174996 115815 174997
rect 115720 174994 115726 174996
rect 115658 174934 115726 174994
rect 115790 174992 115815 174996
rect 115810 174936 115815 174992
rect 115720 174932 115726 174934
rect 115790 174932 115815 174936
rect 115749 174931 115815 174932
rect 213913 174994 213979 174997
rect 230473 174994 230539 174997
rect 230606 174994 230612 174996
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 230473 174992 230612 174994
rect 230473 174936 230478 174992
rect 230534 174936 230612 174992
rect 230473 174934 230612 174936
rect 213913 174931 213979 174934
rect 230473 174931 230539 174934
rect 230606 174932 230612 174934
rect 230676 174932 230682 174996
rect 264973 174858 265039 174861
rect 264973 174856 268180 174858
rect 264973 174800 264978 174856
rect 265034 174800 268180 174856
rect 264973 174798 268180 174800
rect 264973 174795 265039 174798
rect 231117 174722 231183 174725
rect 228804 174720 231183 174722
rect 228804 174664 231122 174720
rect 231178 174664 231183 174720
rect 279374 174692 279434 175203
rect 228804 174662 231183 174664
rect 231117 174659 231183 174662
rect 265065 174450 265131 174453
rect 265065 174448 268180 174450
rect 265065 174392 265070 174448
rect 265126 174392 268180 174448
rect 265065 174390 268180 174392
rect 265065 174387 265131 174390
rect 214005 174314 214071 174317
rect 230657 174314 230723 174317
rect 214005 174312 217212 174314
rect 214005 174256 214010 174312
rect 214066 174256 217212 174312
rect 214005 174254 217212 174256
rect 228804 174312 230723 174314
rect 228804 174256 230662 174312
rect 230718 174256 230723 174312
rect 228804 174254 230723 174256
rect 214005 174251 214071 174254
rect 230657 174251 230723 174254
rect 265157 174042 265223 174045
rect 281758 174042 281764 174044
rect 265157 174040 268180 174042
rect 265157 173984 265162 174040
rect 265218 173984 268180 174040
rect 265157 173982 268180 173984
rect 279956 173982 281764 174042
rect 265157 173979 265223 173982
rect 281758 173980 281764 173982
rect 281828 173980 281834 174044
rect 229185 173770 229251 173773
rect 228804 173768 229251 173770
rect 228804 173712 229190 173768
rect 229246 173712 229251 173768
rect 228804 173710 229251 173712
rect 229185 173707 229251 173710
rect 213913 173634 213979 173637
rect 264973 173634 265039 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 264973 173632 268180 173634
rect 264973 173576 264978 173632
rect 265034 173576 268180 173632
rect 264973 173574 268180 173576
rect 213913 173571 213979 173574
rect 264973 173571 265039 173574
rect 229093 173362 229159 173365
rect 228804 173360 229159 173362
rect 228804 173304 229098 173360
rect 229154 173304 229159 173360
rect 228804 173302 229159 173304
rect 229093 173299 229159 173302
rect 281717 173226 281783 173229
rect 279956 173224 281783 173226
rect 279956 173168 281722 173224
rect 281778 173168 281783 173224
rect 279956 173166 281783 173168
rect 281717 173163 281783 173166
rect 265065 173090 265131 173093
rect 265065 173088 268180 173090
rect 265065 173032 265070 173088
rect 265126 173032 268180 173088
rect 265065 173030 268180 173032
rect 265065 173027 265131 173030
rect 214005 172954 214071 172957
rect 214005 172952 217212 172954
rect 214005 172896 214010 172952
rect 214066 172896 217212 172952
rect 214005 172894 217212 172896
rect 214005 172891 214071 172894
rect 231577 172818 231643 172821
rect 228804 172816 231643 172818
rect 228804 172760 231582 172816
rect 231638 172760 231643 172816
rect 228804 172758 231643 172760
rect 231577 172755 231643 172758
rect 264513 172682 264579 172685
rect 264513 172680 268180 172682
rect 264513 172624 264518 172680
rect 264574 172624 268180 172680
rect 264513 172622 268180 172624
rect 264513 172619 264579 172622
rect 231761 172410 231827 172413
rect 282637 172410 282703 172413
rect 228804 172408 231827 172410
rect 228804 172352 231766 172408
rect 231822 172352 231827 172408
rect 228804 172350 231827 172352
rect 279956 172408 282703 172410
rect 279956 172352 282642 172408
rect 282698 172352 282703 172408
rect 279956 172350 282703 172352
rect 231761 172347 231827 172350
rect 282637 172347 282703 172350
rect 213913 172274 213979 172277
rect 264973 172274 265039 172277
rect 213913 172272 217212 172274
rect 213913 172216 213918 172272
rect 213974 172216 217212 172272
rect 213913 172214 217212 172216
rect 264973 172272 268180 172274
rect 264973 172216 264978 172272
rect 265034 172216 268180 172272
rect 264973 172214 268180 172216
rect 213913 172211 213979 172214
rect 264973 172211 265039 172214
rect 279366 172076 279372 172140
rect 279436 172076 279442 172140
rect 231669 171866 231735 171869
rect 228804 171864 231735 171866
rect 228804 171808 231674 171864
rect 231730 171808 231735 171864
rect 228804 171806 231735 171808
rect 231669 171803 231735 171806
rect 265065 171866 265131 171869
rect 265065 171864 268180 171866
rect 265065 171808 265070 171864
rect 265126 171808 268180 171864
rect 265065 171806 268180 171808
rect 265065 171803 265131 171806
rect 279374 171700 279434 172076
rect 164724 171594 165354 171600
rect 167913 171594 167979 171597
rect 164724 171592 167979 171594
rect 164724 171540 167918 171592
rect 165294 171536 167918 171540
rect 167974 171536 167979 171592
rect 165294 171534 167979 171536
rect 167913 171531 167979 171534
rect 214005 171594 214071 171597
rect 214005 171592 217212 171594
rect 214005 171536 214010 171592
rect 214066 171536 217212 171592
rect 214005 171534 217212 171536
rect 214005 171531 214071 171534
rect 231485 171458 231551 171461
rect 228804 171456 231551 171458
rect 228804 171400 231490 171456
rect 231546 171400 231551 171456
rect 228804 171398 231551 171400
rect 231485 171395 231551 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 213913 171050 213979 171053
rect 265065 171050 265131 171053
rect 213913 171048 217212 171050
rect 213913 170992 213918 171048
rect 213974 170992 217212 171048
rect 213913 170990 217212 170992
rect 265065 171048 268180 171050
rect 265065 170992 265070 171048
rect 265126 170992 268180 171048
rect 265065 170990 268180 170992
rect 213913 170987 213979 170990
rect 265065 170987 265131 170990
rect 231761 170914 231827 170917
rect 280429 170914 280495 170917
rect 228804 170912 231827 170914
rect 228804 170856 231766 170912
rect 231822 170856 231827 170912
rect 228804 170854 231827 170856
rect 279956 170912 280495 170914
rect 279956 170856 280434 170912
rect 280490 170856 280495 170912
rect 279956 170854 280495 170856
rect 231761 170851 231827 170854
rect 280429 170851 280495 170854
rect 231209 170506 231275 170509
rect 228804 170504 231275 170506
rect 228804 170448 231214 170504
rect 231270 170448 231275 170504
rect 228804 170446 231275 170448
rect 231209 170443 231275 170446
rect 265157 170506 265223 170509
rect 265157 170504 268180 170506
rect 265157 170448 265162 170504
rect 265218 170448 268180 170504
rect 265157 170446 268180 170448
rect 265157 170443 265223 170446
rect 214005 170370 214071 170373
rect 214005 170368 217212 170370
rect 214005 170312 214010 170368
rect 214066 170312 217212 170368
rect 214005 170310 217212 170312
rect 214005 170307 214071 170310
rect 264973 170098 265039 170101
rect 281717 170098 281783 170101
rect 264973 170096 268180 170098
rect 264973 170040 264978 170096
rect 265034 170040 268180 170096
rect 264973 170038 268180 170040
rect 279956 170096 281783 170098
rect 279956 170040 281722 170096
rect 281778 170040 281783 170096
rect 279956 170038 281783 170040
rect 264973 170035 265039 170038
rect 281717 170035 281783 170038
rect 231485 169962 231551 169965
rect 228804 169960 231551 169962
rect 228804 169904 231490 169960
rect 231546 169904 231551 169960
rect 228804 169902 231551 169904
rect 231485 169899 231551 169902
rect 213913 169690 213979 169693
rect 265065 169690 265131 169693
rect 213913 169688 217212 169690
rect 213913 169632 213918 169688
rect 213974 169632 217212 169688
rect 213913 169630 217212 169632
rect 265065 169688 268180 169690
rect 265065 169632 265070 169688
rect 265126 169632 268180 169688
rect 265065 169630 268180 169632
rect 213913 169627 213979 169630
rect 265065 169627 265131 169630
rect 231669 169554 231735 169557
rect 228804 169552 231735 169554
rect 228804 169496 231674 169552
rect 231730 169496 231735 169552
rect 228804 169494 231735 169496
rect 231669 169491 231735 169494
rect 282729 169418 282795 169421
rect 279956 169416 282795 169418
rect 279956 169360 282734 169416
rect 282790 169360 282795 169416
rect 279956 169358 282795 169360
rect 282729 169355 282795 169358
rect 264973 169282 265039 169285
rect 264973 169280 268180 169282
rect 264973 169224 264978 169280
rect 265034 169224 268180 169280
rect 264973 169222 268180 169224
rect 264973 169219 265039 169222
rect 214005 169010 214071 169013
rect 231761 169010 231827 169013
rect 214005 169008 217212 169010
rect 214005 168952 214010 169008
rect 214066 168952 217212 169008
rect 214005 168950 217212 168952
rect 228804 169008 231827 169010
rect 228804 168952 231766 169008
rect 231822 168952 231827 169008
rect 228804 168950 231827 168952
rect 214005 168947 214071 168950
rect 231761 168947 231827 168950
rect 265157 168874 265223 168877
rect 265157 168872 268180 168874
rect 265157 168816 265162 168872
rect 265218 168816 268180 168872
rect 265157 168814 268180 168816
rect 265157 168811 265223 168814
rect 231117 168602 231183 168605
rect 282821 168602 282887 168605
rect 228804 168600 231183 168602
rect 228804 168544 231122 168600
rect 231178 168544 231183 168600
rect 228804 168542 231183 168544
rect 279956 168600 282887 168602
rect 279956 168544 282826 168600
rect 282882 168544 282887 168600
rect 279956 168542 282887 168544
rect 231117 168539 231183 168542
rect 282821 168539 282887 168542
rect 265249 168466 265315 168469
rect 265249 168464 268180 168466
rect 265249 168408 265254 168464
rect 265310 168408 268180 168464
rect 265249 168406 268180 168408
rect 265249 168403 265315 168406
rect 213913 168330 213979 168333
rect 213913 168328 217212 168330
rect 213913 168272 213918 168328
rect 213974 168272 217212 168328
rect 213913 168270 217212 168272
rect 213913 168267 213979 168270
rect 231669 168058 231735 168061
rect 228804 168056 231735 168058
rect 228804 168000 231674 168056
rect 231730 168000 231735 168056
rect 228804 167998 231735 168000
rect 231669 167995 231735 167998
rect 265157 167922 265223 167925
rect 265157 167920 268180 167922
rect 265157 167864 265162 167920
rect 265218 167864 268180 167920
rect 265157 167862 268180 167864
rect 265157 167859 265223 167862
rect 282821 167786 282887 167789
rect 279956 167784 282887 167786
rect 279956 167728 282826 167784
rect 282882 167728 282887 167784
rect 279956 167726 282887 167728
rect 282821 167723 282887 167726
rect 214005 167650 214071 167653
rect 231393 167650 231459 167653
rect 214005 167648 217212 167650
rect 214005 167592 214010 167648
rect 214066 167592 217212 167648
rect 214005 167590 217212 167592
rect 228804 167648 231459 167650
rect 228804 167592 231398 167648
rect 231454 167592 231459 167648
rect 228804 167590 231459 167592
rect 214005 167587 214071 167590
rect 231393 167587 231459 167590
rect 264973 167514 265039 167517
rect 264973 167512 268180 167514
rect 264973 167456 264978 167512
rect 265034 167456 268180 167512
rect 264973 167454 268180 167456
rect 264973 167451 265039 167454
rect 231761 167106 231827 167109
rect 228804 167104 231827 167106
rect 228804 167048 231766 167104
rect 231822 167048 231827 167104
rect 228804 167046 231827 167048
rect 231761 167043 231827 167046
rect 265065 167106 265131 167109
rect 282729 167106 282795 167109
rect 265065 167104 268180 167106
rect 265065 167048 265070 167104
rect 265126 167048 268180 167104
rect 265065 167046 268180 167048
rect 279956 167104 282795 167106
rect 279956 167048 282734 167104
rect 282790 167048 282795 167104
rect 279956 167046 282795 167048
rect 265065 167043 265131 167046
rect 282729 167043 282795 167046
rect 213913 166970 213979 166973
rect 213913 166968 217212 166970
rect 213913 166912 213918 166968
rect 213974 166912 217212 166968
rect 213913 166910 217212 166912
rect 213913 166907 213979 166910
rect 279366 166772 279372 166836
rect 279436 166772 279442 166836
rect 231025 166698 231091 166701
rect 228804 166696 231091 166698
rect 228804 166640 231030 166696
rect 231086 166640 231091 166696
rect 228804 166638 231091 166640
rect 231025 166635 231091 166638
rect 265157 166698 265223 166701
rect 265157 166696 268180 166698
rect 265157 166640 265162 166696
rect 265218 166640 268180 166696
rect 265157 166638 268180 166640
rect 265157 166635 265223 166638
rect 214097 166426 214163 166429
rect 214097 166424 217212 166426
rect 214097 166368 214102 166424
rect 214158 166368 217212 166424
rect 214097 166366 217212 166368
rect 214097 166363 214163 166366
rect 265065 166290 265131 166293
rect 265065 166288 268180 166290
rect 265065 166232 265070 166288
rect 265126 166232 268180 166288
rect 279374 166260 279434 166772
rect 265065 166230 268180 166232
rect 265065 166227 265131 166230
rect 231301 166154 231367 166157
rect 228804 166152 231367 166154
rect 228804 166096 231306 166152
rect 231362 166096 231367 166152
rect 228804 166094 231367 166096
rect 231301 166091 231367 166094
rect 264973 165882 265039 165885
rect 583385 165882 583451 165885
rect 583520 165882 584960 165972
rect 264973 165880 268180 165882
rect 264973 165824 264978 165880
rect 265034 165824 268180 165880
rect 264973 165822 268180 165824
rect 583385 165880 584960 165882
rect 583385 165824 583390 165880
rect 583446 165824 584960 165880
rect 583385 165822 584960 165824
rect 264973 165819 265039 165822
rect 583385 165819 583451 165822
rect 214005 165746 214071 165749
rect 230473 165746 230539 165749
rect 214005 165744 217212 165746
rect 214005 165688 214010 165744
rect 214066 165688 217212 165744
rect 214005 165686 217212 165688
rect 228804 165744 230539 165746
rect 228804 165688 230478 165744
rect 230534 165688 230539 165744
rect 583520 165732 584960 165822
rect 228804 165686 230539 165688
rect 214005 165683 214071 165686
rect 230473 165683 230539 165686
rect 282821 165474 282887 165477
rect 279956 165472 282887 165474
rect 279956 165416 282826 165472
rect 282882 165416 282887 165472
rect 279956 165414 282887 165416
rect 282821 165411 282887 165414
rect 264973 165338 265039 165341
rect 264973 165336 268180 165338
rect 264973 165280 264978 165336
rect 265034 165280 268180 165336
rect 264973 165278 268180 165280
rect 264973 165275 265039 165278
rect 231393 165202 231459 165205
rect 228804 165200 231459 165202
rect 228804 165144 231398 165200
rect 231454 165144 231459 165200
rect 228804 165142 231459 165144
rect 231393 165139 231459 165142
rect 213913 165066 213979 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 213913 165003 213979 165006
rect 265065 164930 265131 164933
rect 265065 164928 268180 164930
rect 265065 164872 265070 164928
rect 265126 164872 268180 164928
rect 265065 164870 268180 164872
rect 265065 164867 265131 164870
rect 230933 164794 230999 164797
rect 281993 164794 282059 164797
rect 228804 164792 230999 164794
rect 228804 164736 230938 164792
rect 230994 164736 230999 164792
rect 228804 164734 230999 164736
rect 279956 164792 282059 164794
rect 279956 164736 281998 164792
rect 282054 164736 282059 164792
rect 279956 164734 282059 164736
rect 230933 164731 230999 164734
rect 281993 164731 282059 164734
rect 265617 164522 265683 164525
rect 265617 164520 268180 164522
rect 265617 164464 265622 164520
rect 265678 164464 268180 164520
rect 265617 164462 268180 164464
rect 265617 164459 265683 164462
rect 214005 164386 214071 164389
rect 231301 164386 231367 164389
rect 214005 164384 217212 164386
rect 214005 164328 214010 164384
rect 214066 164328 217212 164384
rect 214005 164326 217212 164328
rect 228804 164384 231367 164386
rect 228804 164328 231306 164384
rect 231362 164328 231367 164384
rect 228804 164326 231367 164328
rect 214005 164323 214071 164326
rect 231301 164323 231367 164326
rect 265157 164114 265223 164117
rect 265157 164112 268180 164114
rect 265157 164056 265162 164112
rect 265218 164056 268180 164112
rect 265157 164054 268180 164056
rect 265157 164051 265223 164054
rect 280337 163978 280403 163981
rect 279956 163976 280403 163978
rect 279956 163920 280342 163976
rect 280398 163920 280403 163976
rect 279956 163918 280403 163920
rect 280337 163915 280403 163918
rect 231393 163842 231459 163845
rect 228804 163840 231459 163842
rect 228804 163784 231398 163840
rect 231454 163784 231459 163840
rect 228804 163782 231459 163784
rect 231393 163779 231459 163782
rect 214557 163706 214623 163709
rect 265065 163706 265131 163709
rect 214557 163704 217212 163706
rect 214557 163648 214562 163704
rect 214618 163648 217212 163704
rect 214557 163646 217212 163648
rect 265065 163704 268180 163706
rect 265065 163648 265070 163704
rect 265126 163648 268180 163704
rect 265065 163646 268180 163648
rect 214557 163643 214623 163646
rect 265065 163643 265131 163646
rect 230606 163434 230612 163436
rect 228804 163374 230612 163434
rect 230606 163372 230612 163374
rect 230676 163372 230682 163436
rect 264973 163298 265039 163301
rect 264973 163296 268180 163298
rect 264973 163240 264978 163296
rect 265034 163240 268180 163296
rect 264973 163238 268180 163240
rect 264973 163235 265039 163238
rect 283782 163162 283788 163164
rect 279956 163102 283788 163162
rect 283782 163100 283788 163102
rect 283852 163100 283858 163164
rect 213913 163026 213979 163029
rect 213913 163024 217212 163026
rect -960 162890 480 162980
rect 213913 162968 213918 163024
rect 213974 162968 217212 163024
rect 213913 162966 217212 162968
rect 213913 162963 213979 162966
rect 3233 162890 3299 162893
rect 231117 162890 231183 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 228804 162888 231183 162890
rect 228804 162832 231122 162888
rect 231178 162832 231183 162888
rect 228804 162830 231183 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 231117 162827 231183 162830
rect 264237 162890 264303 162893
rect 264237 162888 268180 162890
rect 264237 162832 264242 162888
rect 264298 162832 268180 162888
rect 264237 162830 268180 162832
rect 264237 162827 264303 162830
rect 231393 162482 231459 162485
rect 282085 162482 282151 162485
rect 228804 162480 231459 162482
rect 228804 162424 231398 162480
rect 231454 162424 231459 162480
rect 228804 162422 231459 162424
rect 279956 162480 282151 162482
rect 279956 162424 282090 162480
rect 282146 162424 282151 162480
rect 279956 162422 282151 162424
rect 231393 162419 231459 162422
rect 282085 162419 282151 162422
rect 213913 162346 213979 162349
rect 265157 162346 265223 162349
rect 213913 162344 217212 162346
rect 213913 162288 213918 162344
rect 213974 162288 217212 162344
rect 213913 162286 217212 162288
rect 265157 162344 268180 162346
rect 265157 162288 265162 162344
rect 265218 162288 268180 162344
rect 265157 162286 268180 162288
rect 213913 162283 213979 162286
rect 265157 162283 265223 162286
rect 279325 162210 279391 162213
rect 279325 162208 279434 162210
rect 279325 162152 279330 162208
rect 279386 162152 279434 162208
rect 279325 162147 279434 162152
rect 230933 161938 230999 161941
rect 228804 161936 230999 161938
rect 228804 161880 230938 161936
rect 230994 161880 230999 161936
rect 228804 161878 230999 161880
rect 230933 161875 230999 161878
rect 264973 161938 265039 161941
rect 264973 161936 268180 161938
rect 264973 161880 264978 161936
rect 265034 161880 268180 161936
rect 264973 161878 268180 161880
rect 264973 161875 265039 161878
rect 214005 161802 214071 161805
rect 214005 161800 217212 161802
rect 214005 161744 214010 161800
rect 214066 161744 217212 161800
rect 214005 161742 217212 161744
rect 214005 161739 214071 161742
rect 229686 161604 229692 161668
rect 229756 161666 229762 161668
rect 230473 161666 230539 161669
rect 229756 161664 230539 161666
rect 229756 161608 230478 161664
rect 230534 161608 230539 161664
rect 279374 161636 279434 162147
rect 229756 161606 230539 161608
rect 229756 161604 229762 161606
rect 230473 161603 230539 161606
rect 231393 161530 231459 161533
rect 228804 161528 231459 161530
rect 228804 161472 231398 161528
rect 231454 161472 231459 161528
rect 228804 161470 231459 161472
rect 231393 161467 231459 161470
rect 265065 161530 265131 161533
rect 265065 161528 268180 161530
rect 265065 161472 265070 161528
rect 265126 161472 268180 161528
rect 265065 161470 268180 161472
rect 265065 161467 265131 161470
rect 213913 161122 213979 161125
rect 265065 161122 265131 161125
rect 213913 161120 217212 161122
rect 213913 161064 213918 161120
rect 213974 161064 217212 161120
rect 213913 161062 217212 161064
rect 265065 161120 268180 161122
rect 265065 161064 265070 161120
rect 265126 161064 268180 161120
rect 265065 161062 268180 161064
rect 213913 161059 213979 161062
rect 265065 161059 265131 161062
rect 231393 160986 231459 160989
rect 228804 160984 231459 160986
rect 228804 160928 231398 160984
rect 231454 160928 231459 160984
rect 228804 160926 231459 160928
rect 231393 160923 231459 160926
rect 282821 160850 282887 160853
rect 279956 160848 282887 160850
rect 279956 160792 282826 160848
rect 282882 160792 282887 160848
rect 279956 160790 282887 160792
rect 282821 160787 282887 160790
rect 265157 160714 265223 160717
rect 265157 160712 268180 160714
rect 265157 160656 265162 160712
rect 265218 160656 268180 160712
rect 265157 160654 268180 160656
rect 265157 160651 265223 160654
rect 230933 160578 230999 160581
rect 228804 160576 230999 160578
rect 228804 160520 230938 160576
rect 230994 160520 230999 160576
rect 228804 160518 230999 160520
rect 230933 160515 230999 160518
rect 214005 160442 214071 160445
rect 214005 160440 217212 160442
rect 214005 160384 214010 160440
rect 214066 160384 217212 160440
rect 214005 160382 217212 160384
rect 214005 160379 214071 160382
rect 264973 160306 265039 160309
rect 264973 160304 268180 160306
rect 264973 160248 264978 160304
rect 265034 160248 268180 160304
rect 264973 160246 268180 160248
rect 264973 160243 265039 160246
rect 282453 160170 282519 160173
rect 279956 160168 282519 160170
rect 279956 160112 282458 160168
rect 282514 160112 282519 160168
rect 279956 160110 282519 160112
rect 282453 160107 282519 160110
rect 231393 160034 231459 160037
rect 228804 160032 231459 160034
rect 228804 159976 231398 160032
rect 231454 159976 231459 160032
rect 228804 159974 231459 159976
rect 231393 159971 231459 159974
rect 213913 159762 213979 159765
rect 265065 159762 265131 159765
rect 213913 159760 217212 159762
rect 213913 159704 213918 159760
rect 213974 159704 217212 159760
rect 213913 159702 217212 159704
rect 265065 159760 268180 159762
rect 265065 159704 265070 159760
rect 265126 159704 268180 159760
rect 265065 159702 268180 159704
rect 213913 159699 213979 159702
rect 265065 159699 265131 159702
rect 238518 159626 238524 159628
rect 228804 159566 238524 159626
rect 238518 159564 238524 159566
rect 238588 159564 238594 159628
rect 264973 159354 265039 159357
rect 282085 159354 282151 159357
rect 264973 159352 268180 159354
rect 264973 159296 264978 159352
rect 265034 159296 268180 159352
rect 264973 159294 268180 159296
rect 279956 159352 282151 159354
rect 279956 159296 282090 159352
rect 282146 159296 282151 159352
rect 279956 159294 282151 159296
rect 264973 159291 265039 159294
rect 282085 159291 282151 159294
rect 214005 159082 214071 159085
rect 230933 159082 230999 159085
rect 214005 159080 217212 159082
rect 214005 159024 214010 159080
rect 214066 159024 217212 159080
rect 214005 159022 217212 159024
rect 228804 159080 230999 159082
rect 228804 159024 230938 159080
rect 230994 159024 230999 159080
rect 228804 159022 230999 159024
rect 214005 159019 214071 159022
rect 230933 159019 230999 159022
rect 265157 158946 265223 158949
rect 265157 158944 268180 158946
rect 265157 158888 265162 158944
rect 265218 158888 268180 158944
rect 265157 158886 268180 158888
rect 265157 158883 265223 158886
rect 230473 158674 230539 158677
rect 228804 158672 230539 158674
rect 228804 158616 230478 158672
rect 230534 158616 230539 158672
rect 228804 158614 230539 158616
rect 230473 158611 230539 158614
rect 265157 158538 265223 158541
rect 282821 158538 282887 158541
rect 265157 158536 268180 158538
rect 265157 158480 265162 158536
rect 265218 158480 268180 158536
rect 265157 158478 268180 158480
rect 279956 158536 282887 158538
rect 279956 158480 282826 158536
rect 282882 158480 282887 158536
rect 279956 158478 282887 158480
rect 265157 158475 265223 158478
rect 282821 158475 282887 158478
rect 213913 158402 213979 158405
rect 213913 158400 217212 158402
rect 213913 158344 213918 158400
rect 213974 158344 217212 158400
rect 213913 158342 217212 158344
rect 213913 158339 213979 158342
rect 229277 158130 229343 158133
rect 228804 158128 229343 158130
rect 228804 158072 229282 158128
rect 229338 158072 229343 158128
rect 228804 158070 229343 158072
rect 229277 158067 229343 158070
rect 265065 158130 265131 158133
rect 265065 158128 268180 158130
rect 265065 158072 265070 158128
rect 265126 158072 268180 158128
rect 265065 158070 268180 158072
rect 265065 158067 265131 158070
rect 281574 157858 281580 157860
rect 279956 157798 281580 157858
rect 281574 157796 281580 157798
rect 281644 157796 281650 157860
rect 214005 157722 214071 157725
rect 230565 157722 230631 157725
rect 214005 157720 217212 157722
rect 214005 157664 214010 157720
rect 214066 157664 217212 157720
rect 214005 157662 217212 157664
rect 228804 157720 230631 157722
rect 228804 157664 230570 157720
rect 230626 157664 230631 157720
rect 228804 157662 230631 157664
rect 214005 157659 214071 157662
rect 230565 157659 230631 157662
rect 264973 157722 265039 157725
rect 264973 157720 268180 157722
rect 264973 157664 264978 157720
rect 265034 157664 268180 157720
rect 264973 157662 268180 157664
rect 264973 157659 265039 157662
rect 214925 157178 214991 157181
rect 231761 157178 231827 157181
rect 214925 157176 217212 157178
rect 214925 157120 214930 157176
rect 214986 157120 217212 157176
rect 214925 157118 217212 157120
rect 228804 157176 231827 157178
rect 228804 157120 231766 157176
rect 231822 157120 231827 157176
rect 228804 157118 231827 157120
rect 214925 157115 214991 157118
rect 231761 157115 231827 157118
rect 265157 157178 265223 157181
rect 265157 157176 268180 157178
rect 265157 157120 265162 157176
rect 265218 157120 268180 157176
rect 265157 157118 268180 157120
rect 265157 157115 265223 157118
rect 281533 157042 281599 157045
rect 279956 157040 281599 157042
rect 279956 156984 281538 157040
rect 281594 156984 281599 157040
rect 279956 156982 281599 156984
rect 281533 156979 281599 156982
rect 231117 156770 231183 156773
rect 228804 156768 231183 156770
rect 228804 156712 231122 156768
rect 231178 156712 231183 156768
rect 228804 156710 231183 156712
rect 231117 156707 231183 156710
rect 265065 156770 265131 156773
rect 265065 156768 268180 156770
rect 265065 156712 265070 156768
rect 265126 156712 268180 156768
rect 265065 156710 268180 156712
rect 265065 156707 265131 156710
rect 213913 156498 213979 156501
rect 213913 156496 217212 156498
rect 213913 156440 213918 156496
rect 213974 156440 217212 156496
rect 213913 156438 217212 156440
rect 213913 156435 213979 156438
rect 264973 156362 265039 156365
rect 280245 156362 280311 156365
rect 264973 156360 268180 156362
rect 264973 156304 264978 156360
rect 265034 156304 268180 156360
rect 264973 156302 268180 156304
rect 279956 156360 280311 156362
rect 279956 156304 280250 156360
rect 280306 156304 280311 156360
rect 279956 156302 280311 156304
rect 264973 156299 265039 156302
rect 280245 156299 280311 156302
rect 230422 156226 230428 156228
rect 228804 156166 230428 156226
rect 230422 156164 230428 156166
rect 230492 156164 230498 156228
rect 265065 155954 265131 155957
rect 265065 155952 268180 155954
rect 265065 155896 265070 155952
rect 265126 155896 268180 155952
rect 265065 155894 268180 155896
rect 265065 155891 265131 155894
rect 213913 155818 213979 155821
rect 229185 155818 229251 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 228804 155816 229251 155818
rect 228804 155760 229190 155816
rect 229246 155760 229251 155816
rect 228804 155758 229251 155760
rect 213913 155755 213979 155758
rect 229185 155755 229251 155758
rect 264973 155546 265039 155549
rect 281717 155546 281783 155549
rect 264973 155544 268180 155546
rect 264973 155488 264978 155544
rect 265034 155488 268180 155544
rect 264973 155486 268180 155488
rect 279956 155544 281783 155546
rect 279956 155488 281722 155544
rect 281778 155488 281783 155544
rect 279956 155486 281783 155488
rect 264973 155483 265039 155486
rect 281717 155483 281783 155486
rect 229093 155274 229159 155277
rect 228804 155272 229159 155274
rect 228804 155216 229098 155272
rect 229154 155216 229159 155272
rect 228804 155214 229159 155216
rect 229093 155211 229159 155214
rect 279325 155274 279391 155277
rect 279325 155272 279434 155274
rect 279325 155216 279330 155272
rect 279386 155216 279434 155272
rect 279325 155211 279434 155216
rect 214005 155138 214071 155141
rect 265157 155138 265223 155141
rect 214005 155136 217212 155138
rect 214005 155080 214010 155136
rect 214066 155080 217212 155136
rect 214005 155078 217212 155080
rect 265157 155136 268180 155138
rect 265157 155080 265162 155136
rect 265218 155080 268180 155136
rect 265157 155078 268180 155080
rect 214005 155075 214071 155078
rect 265157 155075 265223 155078
rect 230933 154866 230999 154869
rect 228804 154864 230999 154866
rect 228804 154808 230938 154864
rect 230994 154808 230999 154864
rect 228804 154806 230999 154808
rect 230933 154803 230999 154806
rect 279374 154700 279434 155211
rect 265341 154594 265407 154597
rect 265341 154592 268180 154594
rect 265341 154536 265346 154592
rect 265402 154536 268180 154592
rect 265341 154534 268180 154536
rect 265341 154531 265407 154534
rect 214005 154458 214071 154461
rect 214005 154456 217212 154458
rect 214005 154400 214010 154456
rect 214066 154400 217212 154456
rect 214005 154398 217212 154400
rect 214005 154395 214071 154398
rect 231761 154322 231827 154325
rect 228804 154320 231827 154322
rect 228804 154264 231766 154320
rect 231822 154264 231827 154320
rect 228804 154262 231827 154264
rect 231761 154259 231827 154262
rect 265065 154186 265131 154189
rect 265065 154184 268180 154186
rect 265065 154128 265070 154184
rect 265126 154128 268180 154184
rect 265065 154126 268180 154128
rect 265065 154123 265131 154126
rect 281717 154050 281783 154053
rect 279956 154048 281783 154050
rect 279956 153992 281722 154048
rect 281778 153992 281783 154048
rect 279956 153990 281783 153992
rect 281717 153987 281783 153990
rect 240358 153914 240364 153916
rect 228804 153854 240364 153914
rect 240358 153852 240364 153854
rect 240428 153852 240434 153916
rect 213913 153778 213979 153781
rect 231669 153778 231735 153781
rect 244222 153778 244228 153780
rect 213913 153776 217212 153778
rect 213913 153720 213918 153776
rect 213974 153720 217212 153776
rect 213913 153718 217212 153720
rect 231669 153776 244228 153778
rect 231669 153720 231674 153776
rect 231730 153720 244228 153776
rect 231669 153718 244228 153720
rect 213913 153715 213979 153718
rect 231669 153715 231735 153718
rect 244222 153716 244228 153718
rect 244292 153716 244298 153780
rect 265157 153778 265223 153781
rect 279417 153778 279483 153781
rect 265157 153776 268180 153778
rect 265157 153720 265162 153776
rect 265218 153720 268180 153776
rect 265157 153718 268180 153720
rect 279374 153776 279483 153778
rect 279374 153720 279422 153776
rect 279478 153720 279483 153776
rect 265157 153715 265223 153718
rect 279374 153715 279483 153720
rect 231485 153370 231551 153373
rect 228804 153368 231551 153370
rect 228804 153312 231490 153368
rect 231546 153312 231551 153368
rect 228804 153310 231551 153312
rect 231485 153307 231551 153310
rect 264973 153370 265039 153373
rect 264973 153368 268180 153370
rect 264973 153312 264978 153368
rect 265034 153312 268180 153368
rect 264973 153310 268180 153312
rect 264973 153307 265039 153310
rect 279374 153204 279434 153715
rect 214005 153098 214071 153101
rect 214005 153096 217212 153098
rect 214005 153040 214010 153096
rect 214066 153040 217212 153096
rect 214005 153038 217212 153040
rect 214005 153035 214071 153038
rect 231669 152962 231735 152965
rect 228804 152960 231735 152962
rect 228804 152904 231674 152960
rect 231730 152904 231735 152960
rect 228804 152902 231735 152904
rect 231669 152899 231735 152902
rect 265065 152962 265131 152965
rect 265065 152960 268180 152962
rect 265065 152904 265070 152960
rect 265126 152904 268180 152960
rect 265065 152902 268180 152904
rect 265065 152899 265131 152902
rect 583385 152690 583451 152693
rect 583520 152690 584960 152780
rect 583385 152688 584960 152690
rect 583385 152632 583390 152688
rect 583446 152632 584960 152688
rect 583385 152630 584960 152632
rect 583385 152627 583451 152630
rect 213913 152554 213979 152557
rect 231761 152554 231827 152557
rect 213913 152552 217212 152554
rect 213913 152496 213918 152552
rect 213974 152496 217212 152552
rect 213913 152494 217212 152496
rect 228804 152552 231827 152554
rect 228804 152496 231766 152552
rect 231822 152496 231827 152552
rect 228804 152494 231827 152496
rect 213913 152491 213979 152494
rect 231761 152491 231827 152494
rect 265249 152554 265315 152557
rect 265249 152552 268180 152554
rect 265249 152496 265254 152552
rect 265310 152496 268180 152552
rect 583520 152540 584960 152630
rect 265249 152494 268180 152496
rect 265249 152491 265315 152494
rect 281625 152418 281691 152421
rect 279956 152416 281691 152418
rect 279956 152360 281630 152416
rect 281686 152360 281691 152416
rect 279956 152358 281691 152360
rect 281625 152355 281691 152358
rect 231393 152010 231459 152013
rect 228804 152008 231459 152010
rect 228804 151952 231398 152008
rect 231454 151952 231459 152008
rect 228804 151950 231459 151952
rect 231393 151947 231459 151950
rect 264973 152010 265039 152013
rect 264973 152008 268180 152010
rect 264973 151952 264978 152008
rect 265034 151952 268180 152008
rect 264973 151950 268180 151952
rect 264973 151947 265039 151950
rect 214465 151874 214531 151877
rect 214465 151872 217212 151874
rect 214465 151816 214470 151872
rect 214526 151816 217212 151872
rect 214465 151814 217212 151816
rect 214465 151811 214531 151814
rect 282821 151738 282887 151741
rect 279956 151736 282887 151738
rect 279956 151680 282826 151736
rect 282882 151680 282887 151736
rect 279956 151678 282887 151680
rect 282821 151675 282887 151678
rect 231209 151602 231275 151605
rect 228804 151600 231275 151602
rect 228804 151544 231214 151600
rect 231270 151544 231275 151600
rect 228804 151542 231275 151544
rect 231209 151539 231275 151542
rect 266077 151602 266143 151605
rect 266077 151600 268180 151602
rect 266077 151544 266082 151600
rect 266138 151544 268180 151600
rect 266077 151542 268180 151544
rect 266077 151539 266143 151542
rect 215201 151194 215267 151197
rect 265341 151194 265407 151197
rect 215201 151192 217212 151194
rect 215201 151136 215206 151192
rect 215262 151136 217212 151192
rect 215201 151134 217212 151136
rect 265341 151192 268180 151194
rect 265341 151136 265346 151192
rect 265402 151136 268180 151192
rect 265341 151134 268180 151136
rect 215201 151131 215267 151134
rect 265341 151131 265407 151134
rect 231894 151058 231900 151060
rect 228804 150998 231900 151058
rect 231894 150996 231900 150998
rect 231964 150996 231970 151060
rect 282637 150922 282703 150925
rect 279956 150920 282703 150922
rect 279956 150864 282642 150920
rect 282698 150864 282703 150920
rect 279956 150862 282703 150864
rect 282637 150859 282703 150862
rect 264973 150786 265039 150789
rect 264973 150784 268180 150786
rect 264973 150728 264978 150784
rect 265034 150728 268180 150784
rect 264973 150726 268180 150728
rect 264973 150723 265039 150726
rect 232037 150650 232103 150653
rect 228804 150648 232103 150650
rect 228804 150592 232042 150648
rect 232098 150592 232103 150648
rect 228804 150590 232103 150592
rect 232037 150587 232103 150590
rect 213913 150514 213979 150517
rect 213913 150512 217212 150514
rect 213913 150456 213918 150512
rect 213974 150456 217212 150512
rect 213913 150454 217212 150456
rect 213913 150451 213979 150454
rect 265065 150378 265131 150381
rect 265065 150376 268180 150378
rect 265065 150320 265070 150376
rect 265126 150320 268180 150376
rect 265065 150318 268180 150320
rect 265065 150315 265131 150318
rect 230933 150106 230999 150109
rect 282821 150106 282887 150109
rect 228804 150104 230999 150106
rect 228804 150048 230938 150104
rect 230994 150048 230999 150104
rect 228804 150046 230999 150048
rect 279956 150104 282887 150106
rect 279956 150048 282826 150104
rect 282882 150048 282887 150104
rect 279956 150046 282887 150048
rect 230933 150043 230999 150046
rect 282821 150043 282887 150046
rect 265433 149970 265499 149973
rect 265433 149968 268180 149970
rect -960 149834 480 149924
rect 265433 149912 265438 149968
rect 265494 149912 268180 149968
rect 265433 149910 268180 149912
rect 265433 149907 265499 149910
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 213913 149834 213979 149837
rect 213913 149832 217212 149834
rect 213913 149776 213918 149832
rect 213974 149776 217212 149832
rect 213913 149774 217212 149776
rect 213913 149771 213979 149774
rect 230749 149698 230815 149701
rect 228804 149696 230815 149698
rect 228804 149640 230754 149696
rect 230810 149640 230815 149696
rect 228804 149638 230815 149640
rect 230749 149635 230815 149638
rect 264973 149562 265039 149565
rect 264973 149560 268180 149562
rect 264973 149504 264978 149560
rect 265034 149504 268180 149560
rect 264973 149502 268180 149504
rect 264973 149499 265039 149502
rect 281717 149426 281783 149429
rect 279956 149424 281783 149426
rect 279956 149368 281722 149424
rect 281778 149368 281783 149424
rect 279956 149366 281783 149368
rect 281717 149363 281783 149366
rect 214005 149154 214071 149157
rect 230841 149154 230907 149157
rect 214005 149152 217212 149154
rect 214005 149096 214010 149152
rect 214066 149096 217212 149152
rect 214005 149094 217212 149096
rect 228804 149152 230907 149154
rect 228804 149096 230846 149152
rect 230902 149096 230907 149152
rect 228804 149094 230907 149096
rect 214005 149091 214071 149094
rect 230841 149091 230907 149094
rect 265065 149018 265131 149021
rect 265065 149016 268180 149018
rect 265065 148960 265070 149016
rect 265126 148960 268180 149016
rect 265065 148958 268180 148960
rect 265065 148955 265131 148958
rect 231761 148746 231827 148749
rect 228804 148744 231827 148746
rect 228804 148688 231766 148744
rect 231822 148688 231827 148744
rect 228804 148686 231827 148688
rect 231761 148683 231827 148686
rect 265157 148610 265223 148613
rect 282821 148610 282887 148613
rect 265157 148608 268180 148610
rect 265157 148552 265162 148608
rect 265218 148552 268180 148608
rect 265157 148550 268180 148552
rect 279956 148608 282887 148610
rect 279956 148552 282826 148608
rect 282882 148552 282887 148608
rect 279956 148550 282887 148552
rect 265157 148547 265223 148550
rect 282821 148547 282887 148550
rect 213913 148474 213979 148477
rect 213913 148472 217212 148474
rect 213913 148416 213918 148472
rect 213974 148416 217212 148472
rect 213913 148414 217212 148416
rect 213913 148411 213979 148414
rect 231117 148202 231183 148205
rect 228804 148200 231183 148202
rect 228804 148144 231122 148200
rect 231178 148144 231183 148200
rect 228804 148142 231183 148144
rect 231117 148139 231183 148142
rect 264973 148202 265039 148205
rect 264973 148200 268180 148202
rect 264973 148144 264978 148200
rect 265034 148144 268180 148200
rect 264973 148142 268180 148144
rect 264973 148139 265039 148142
rect 213913 147930 213979 147933
rect 213913 147928 217212 147930
rect 213913 147872 213918 147928
rect 213974 147872 217212 147928
rect 213913 147870 217212 147872
rect 213913 147867 213979 147870
rect 245694 147794 245700 147796
rect 228804 147734 245700 147794
rect 245694 147732 245700 147734
rect 245764 147732 245770 147796
rect 265801 147794 265867 147797
rect 282729 147794 282795 147797
rect 265801 147792 268180 147794
rect 265801 147736 265806 147792
rect 265862 147736 268180 147792
rect 265801 147734 268180 147736
rect 279956 147792 282795 147794
rect 279956 147736 282734 147792
rect 282790 147736 282795 147792
rect 279956 147734 282795 147736
rect 265801 147731 265867 147734
rect 282729 147731 282795 147734
rect 265065 147386 265131 147389
rect 265065 147384 268180 147386
rect 265065 147328 265070 147384
rect 265126 147328 268180 147384
rect 265065 147326 268180 147328
rect 265065 147323 265131 147326
rect 214005 147250 214071 147253
rect 233182 147250 233188 147252
rect 214005 147248 217212 147250
rect 214005 147192 214010 147248
rect 214066 147192 217212 147248
rect 214005 147190 217212 147192
rect 228804 147190 233188 147250
rect 214005 147187 214071 147190
rect 233182 147188 233188 147190
rect 233252 147188 233258 147252
rect 265249 146978 265315 146981
rect 265249 146976 268180 146978
rect 265249 146920 265254 146976
rect 265310 146920 268180 146976
rect 265249 146918 268180 146920
rect 265249 146915 265315 146918
rect 231761 146842 231827 146845
rect 228804 146840 231827 146842
rect 228804 146784 231766 146840
rect 231822 146784 231827 146840
rect 228804 146782 231827 146784
rect 231761 146779 231827 146782
rect 213913 146570 213979 146573
rect 213913 146568 217212 146570
rect 213913 146512 213918 146568
rect 213974 146512 217212 146568
rect 213913 146510 217212 146512
rect 213913 146507 213979 146510
rect 264973 146434 265039 146437
rect 279926 146434 279986 147084
rect 291142 146434 291148 146436
rect 264973 146432 268180 146434
rect 264973 146376 264978 146432
rect 265034 146376 268180 146432
rect 264973 146374 268180 146376
rect 279926 146374 291148 146434
rect 264973 146371 265039 146374
rect 291142 146372 291148 146374
rect 291212 146372 291218 146436
rect 229829 146298 229895 146301
rect 282821 146298 282887 146301
rect 228804 146296 229895 146298
rect 228804 146240 229834 146296
rect 229890 146240 229895 146296
rect 228804 146238 229895 146240
rect 279956 146296 282887 146298
rect 279956 146240 282826 146296
rect 282882 146240 282887 146296
rect 279956 146238 282887 146240
rect 229829 146235 229895 146238
rect 282821 146235 282887 146238
rect 265157 146026 265223 146029
rect 265157 146024 268180 146026
rect 265157 145968 265162 146024
rect 265218 145968 268180 146024
rect 265157 145966 268180 145968
rect 265157 145963 265223 145966
rect 214005 145890 214071 145893
rect 231761 145890 231827 145893
rect 214005 145888 217212 145890
rect 214005 145832 214010 145888
rect 214066 145832 217212 145888
rect 214005 145830 217212 145832
rect 228804 145888 231827 145890
rect 228804 145832 231766 145888
rect 231822 145832 231827 145888
rect 228804 145830 231827 145832
rect 214005 145827 214071 145830
rect 231761 145827 231827 145830
rect 230933 145618 230999 145621
rect 249742 145618 249748 145620
rect 230933 145616 249748 145618
rect 230933 145560 230938 145616
rect 230994 145560 249748 145616
rect 230933 145558 249748 145560
rect 230933 145555 230999 145558
rect 249742 145556 249748 145558
rect 249812 145556 249818 145620
rect 265065 145618 265131 145621
rect 265065 145616 268180 145618
rect 265065 145560 265070 145616
rect 265126 145560 268180 145616
rect 265065 145558 268180 145560
rect 265065 145555 265131 145558
rect 281993 145482 282059 145485
rect 279956 145480 282059 145482
rect 279956 145424 281998 145480
rect 282054 145424 282059 145480
rect 279956 145422 282059 145424
rect 281993 145419 282059 145422
rect 233366 145346 233372 145348
rect 228804 145286 233372 145346
rect 233366 145284 233372 145286
rect 233436 145284 233442 145348
rect 213913 145210 213979 145213
rect 264973 145210 265039 145213
rect 213913 145208 217212 145210
rect 213913 145152 213918 145208
rect 213974 145152 217212 145208
rect 213913 145150 217212 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 213913 145147 213979 145150
rect 264973 145147 265039 145150
rect 231669 144938 231735 144941
rect 228804 144936 231735 144938
rect 228804 144880 231674 144936
rect 231730 144880 231735 144936
rect 228804 144878 231735 144880
rect 231669 144875 231735 144878
rect 230422 144740 230428 144804
rect 230492 144802 230498 144804
rect 234654 144802 234660 144804
rect 230492 144742 234660 144802
rect 230492 144740 230498 144742
rect 234654 144740 234660 144742
rect 234724 144740 234730 144804
rect 265065 144802 265131 144805
rect 284334 144802 284340 144804
rect 265065 144800 268180 144802
rect 265065 144744 265070 144800
rect 265126 144744 268180 144800
rect 265065 144742 268180 144744
rect 279956 144742 284340 144802
rect 265065 144739 265131 144742
rect 284334 144740 284340 144742
rect 284404 144740 284410 144804
rect 214005 144530 214071 144533
rect 214005 144528 217212 144530
rect 214005 144472 214010 144528
rect 214066 144472 217212 144528
rect 214005 144470 217212 144472
rect 214005 144467 214071 144470
rect 231301 144394 231367 144397
rect 228804 144392 231367 144394
rect 228804 144336 231306 144392
rect 231362 144336 231367 144392
rect 228804 144334 231367 144336
rect 231301 144331 231367 144334
rect 264973 144394 265039 144397
rect 264973 144392 268180 144394
rect 264973 144336 264978 144392
rect 265034 144336 268180 144392
rect 264973 144334 268180 144336
rect 264973 144331 265039 144334
rect 231485 143986 231551 143989
rect 282821 143986 282887 143989
rect 228804 143984 231551 143986
rect 228804 143928 231490 143984
rect 231546 143928 231551 143984
rect 228804 143926 231551 143928
rect 279956 143984 282887 143986
rect 279956 143928 282826 143984
rect 282882 143928 282887 143984
rect 279956 143926 282887 143928
rect 231485 143923 231551 143926
rect 282821 143923 282887 143926
rect 213913 143850 213979 143853
rect 265709 143850 265775 143853
rect 213913 143848 217212 143850
rect 213913 143792 213918 143848
rect 213974 143792 217212 143848
rect 213913 143790 217212 143792
rect 265709 143848 268180 143850
rect 265709 143792 265714 143848
rect 265770 143792 268180 143848
rect 265709 143790 268180 143792
rect 213913 143787 213979 143790
rect 265709 143787 265775 143790
rect 248638 143442 248644 143444
rect 228804 143382 248644 143442
rect 248638 143380 248644 143382
rect 248708 143380 248714 143444
rect 265157 143442 265223 143445
rect 265157 143440 268180 143442
rect 265157 143384 265162 143440
rect 265218 143384 268180 143440
rect 265157 143382 268180 143384
rect 265157 143379 265223 143382
rect 213913 143306 213979 143309
rect 213913 143304 217212 143306
rect 213913 143248 213918 143304
rect 213974 143248 217212 143304
rect 213913 143246 217212 143248
rect 213913 143243 213979 143246
rect 285622 143170 285628 143172
rect 279956 143110 285628 143170
rect 285622 143108 285628 143110
rect 285692 143108 285698 143172
rect 230933 143034 230999 143037
rect 228804 143032 230999 143034
rect 228804 142976 230938 143032
rect 230994 142976 230999 143032
rect 228804 142974 230999 142976
rect 230933 142971 230999 142974
rect 264973 143034 265039 143037
rect 264973 143032 268180 143034
rect 264973 142976 264978 143032
rect 265034 142976 268180 143032
rect 264973 142974 268180 142976
rect 264973 142971 265039 142974
rect 214925 142626 214991 142629
rect 265065 142626 265131 142629
rect 214925 142624 217212 142626
rect 214925 142568 214930 142624
rect 214986 142568 217212 142624
rect 214925 142566 217212 142568
rect 265065 142624 268180 142626
rect 265065 142568 265070 142624
rect 265126 142568 268180 142624
rect 265065 142566 268180 142568
rect 214925 142563 214991 142566
rect 265065 142563 265131 142566
rect 231301 142490 231367 142493
rect 281625 142490 281691 142493
rect 228804 142488 231367 142490
rect 228804 142432 231306 142488
rect 231362 142432 231367 142488
rect 228804 142430 231367 142432
rect 279956 142488 281691 142490
rect 279956 142432 281630 142488
rect 281686 142432 281691 142488
rect 279956 142430 281691 142432
rect 231301 142427 231367 142430
rect 281625 142427 281691 142430
rect 265893 142218 265959 142221
rect 265893 142216 268180 142218
rect 265893 142160 265898 142216
rect 265954 142160 268180 142216
rect 265893 142158 268180 142160
rect 265893 142155 265959 142158
rect 248454 142082 248460 142084
rect 228804 142022 248460 142082
rect 248454 142020 248460 142022
rect 248524 142020 248530 142084
rect 214005 141946 214071 141949
rect 214005 141944 217212 141946
rect 214005 141888 214010 141944
rect 214066 141888 217212 141944
rect 214005 141886 217212 141888
rect 214005 141883 214071 141886
rect 265065 141810 265131 141813
rect 265065 141808 268180 141810
rect 265065 141752 265070 141808
rect 265126 141752 268180 141808
rect 265065 141750 268180 141752
rect 265065 141747 265131 141750
rect 230422 141674 230428 141676
rect 228804 141614 230428 141674
rect 230422 141612 230428 141614
rect 230492 141612 230498 141676
rect 282821 141674 282887 141677
rect 279956 141672 282887 141674
rect 279956 141616 282826 141672
rect 282882 141616 282887 141672
rect 279956 141614 282887 141616
rect 282821 141611 282887 141614
rect 230974 141340 230980 141404
rect 231044 141402 231050 141404
rect 241145 141402 241211 141405
rect 231044 141400 241211 141402
rect 231044 141344 241150 141400
rect 241206 141344 241211 141400
rect 231044 141342 241211 141344
rect 231044 141340 231050 141342
rect 241145 141339 241211 141342
rect 213913 141266 213979 141269
rect 265157 141266 265223 141269
rect 213913 141264 217212 141266
rect 213913 141208 213918 141264
rect 213974 141208 217212 141264
rect 213913 141206 217212 141208
rect 265157 141264 268180 141266
rect 265157 141208 265162 141264
rect 265218 141208 268180 141264
rect 265157 141206 268180 141208
rect 213913 141203 213979 141206
rect 265157 141203 265223 141206
rect 231761 141130 231827 141133
rect 228804 141128 231827 141130
rect 228804 141072 231766 141128
rect 231822 141072 231827 141128
rect 228804 141070 231827 141072
rect 231761 141067 231827 141070
rect 264973 140858 265039 140861
rect 282729 140858 282795 140861
rect 264973 140856 268180 140858
rect 264973 140800 264978 140856
rect 265034 140800 268180 140856
rect 264973 140798 268180 140800
rect 279956 140856 282795 140858
rect 279956 140800 282734 140856
rect 282790 140800 282795 140856
rect 279956 140798 282795 140800
rect 264973 140795 265039 140798
rect 282729 140795 282795 140798
rect 231761 140722 231827 140725
rect 228804 140720 231827 140722
rect 228804 140664 231766 140720
rect 231822 140664 231827 140720
rect 228804 140662 231827 140664
rect 231761 140659 231827 140662
rect 214005 140586 214071 140589
rect 214005 140584 217212 140586
rect 214005 140528 214010 140584
rect 214066 140528 217212 140584
rect 214005 140526 217212 140528
rect 214005 140523 214071 140526
rect 231669 140178 231735 140181
rect 268150 140178 268210 140420
rect 281901 140178 281967 140181
rect 228804 140176 231735 140178
rect 228804 140120 231674 140176
rect 231730 140120 231735 140176
rect 228804 140118 231735 140120
rect 231669 140115 231735 140118
rect 238710 140118 268210 140178
rect 279956 140176 281967 140178
rect 279956 140120 281906 140176
rect 281962 140120 281967 140176
rect 279956 140118 281967 140120
rect 229686 139980 229692 140044
rect 229756 140042 229762 140044
rect 238710 140042 238770 140118
rect 281901 140115 281967 140118
rect 229756 139982 238770 140042
rect 264973 140042 265039 140045
rect 264973 140040 268180 140042
rect 264973 139984 264978 140040
rect 265034 139984 268180 140040
rect 264973 139982 268180 139984
rect 229756 139980 229762 139982
rect 264973 139979 265039 139982
rect 213913 139906 213979 139909
rect 213913 139904 217212 139906
rect 213913 139848 213918 139904
rect 213974 139848 217212 139904
rect 213913 139846 217212 139848
rect 213913 139843 213979 139846
rect 236494 139770 236500 139772
rect 228804 139710 236500 139770
rect 236494 139708 236500 139710
rect 236564 139708 236570 139772
rect 246246 139572 246252 139636
rect 246316 139634 246322 139636
rect 246316 139574 268180 139634
rect 246316 139572 246322 139574
rect 282821 139362 282887 139365
rect 279956 139360 282887 139362
rect 279956 139304 282826 139360
rect 282882 139304 282887 139360
rect 279956 139302 282887 139304
rect 282821 139299 282887 139302
rect 583385 139362 583451 139365
rect 583520 139362 584960 139452
rect 583385 139360 584960 139362
rect 583385 139304 583390 139360
rect 583446 139304 584960 139360
rect 583385 139302 584960 139304
rect 583385 139299 583451 139302
rect 214005 139226 214071 139229
rect 232078 139226 232084 139228
rect 214005 139224 217212 139226
rect 214005 139168 214010 139224
rect 214066 139168 217212 139224
rect 214005 139166 217212 139168
rect 228804 139166 232084 139226
rect 214005 139163 214071 139166
rect 232078 139164 232084 139166
rect 232148 139164 232154 139228
rect 265065 139226 265131 139229
rect 265065 139224 268180 139226
rect 265065 139168 265070 139224
rect 265126 139168 268180 139224
rect 583520 139212 584960 139302
rect 265065 139166 268180 139168
rect 265065 139163 265131 139166
rect 237598 138818 237604 138820
rect 228804 138758 237604 138818
rect 237598 138756 237604 138758
rect 237668 138756 237674 138820
rect 214557 138682 214623 138685
rect 267273 138682 267339 138685
rect 214557 138680 217212 138682
rect 214557 138624 214562 138680
rect 214618 138624 217212 138680
rect 214557 138622 217212 138624
rect 267273 138680 268180 138682
rect 267273 138624 267278 138680
rect 267334 138624 268180 138680
rect 267273 138622 268180 138624
rect 214557 138619 214623 138622
rect 267273 138619 267339 138622
rect 284518 138546 284524 138548
rect 279956 138486 284524 138546
rect 284518 138484 284524 138486
rect 284588 138484 284594 138548
rect 231761 138274 231827 138277
rect 228804 138272 231827 138274
rect 228804 138216 231766 138272
rect 231822 138216 231827 138272
rect 228804 138214 231827 138216
rect 231761 138211 231827 138214
rect 264973 138274 265039 138277
rect 264973 138272 268180 138274
rect 264973 138216 264978 138272
rect 265034 138216 268180 138272
rect 264973 138214 268180 138216
rect 264973 138211 265039 138214
rect 213913 138002 213979 138005
rect 213913 138000 217212 138002
rect 213913 137944 213918 138000
rect 213974 137944 217212 138000
rect 213913 137942 217212 137944
rect 213913 137939 213979 137942
rect 231669 137866 231735 137869
rect 228804 137864 231735 137866
rect 228804 137808 231674 137864
rect 231730 137808 231735 137864
rect 228804 137806 231735 137808
rect 231669 137803 231735 137806
rect 265249 137866 265315 137869
rect 282821 137866 282887 137869
rect 265249 137864 268180 137866
rect 265249 137808 265254 137864
rect 265310 137808 268180 137864
rect 265249 137806 268180 137808
rect 279956 137864 282887 137866
rect 279956 137808 282826 137864
rect 282882 137808 282887 137864
rect 279956 137806 282887 137808
rect 265249 137803 265315 137806
rect 282821 137803 282887 137806
rect 265065 137458 265131 137461
rect 265065 137456 268180 137458
rect 265065 137400 265070 137456
rect 265126 137400 268180 137456
rect 265065 137398 268180 137400
rect 265065 137395 265131 137398
rect 214097 137322 214163 137325
rect 229134 137322 229140 137324
rect 214097 137320 217212 137322
rect 214097 137264 214102 137320
rect 214158 137264 217212 137320
rect 214097 137262 217212 137264
rect 228804 137262 229140 137322
rect 214097 137259 214163 137262
rect 229134 137260 229140 137262
rect 229204 137260 229210 137324
rect 231158 137260 231164 137324
rect 231228 137322 231234 137324
rect 241237 137322 241303 137325
rect 231228 137320 241303 137322
rect 231228 137264 241242 137320
rect 241298 137264 241303 137320
rect 231228 137262 241303 137264
rect 231228 137260 231234 137262
rect 241237 137259 241303 137262
rect 264973 137050 265039 137053
rect 280153 137050 280219 137053
rect 264973 137048 268180 137050
rect 264973 136992 264978 137048
rect 265034 136992 268180 137048
rect 264973 136990 268180 136992
rect 279956 137048 280219 137050
rect 279956 136992 280158 137048
rect 280214 136992 280219 137048
rect 279956 136990 280219 136992
rect 264973 136987 265039 136990
rect 280153 136987 280219 136990
rect 229737 136914 229803 136917
rect 228804 136912 229803 136914
rect -960 136778 480 136868
rect 228804 136856 229742 136912
rect 229798 136856 229803 136912
rect 228804 136854 229803 136856
rect 229737 136851 229803 136854
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 214005 136642 214071 136645
rect 265157 136642 265223 136645
rect 214005 136640 217212 136642
rect 214005 136584 214010 136640
rect 214066 136584 217212 136640
rect 214005 136582 217212 136584
rect 265157 136640 268180 136642
rect 265157 136584 265162 136640
rect 265218 136584 268180 136640
rect 265157 136582 268180 136584
rect 214005 136579 214071 136582
rect 265157 136579 265223 136582
rect 241646 136370 241652 136372
rect 228804 136310 241652 136370
rect 241646 136308 241652 136310
rect 241716 136308 241722 136372
rect 282545 136370 282611 136373
rect 279956 136368 282611 136370
rect 279956 136312 282550 136368
rect 282606 136312 282611 136368
rect 279956 136310 282611 136312
rect 282545 136307 282611 136310
rect 265065 136234 265131 136237
rect 265065 136232 268180 136234
rect 265065 136176 265070 136232
rect 265126 136176 268180 136232
rect 265065 136174 268180 136176
rect 265065 136171 265131 136174
rect 216029 135962 216095 135965
rect 231209 135962 231275 135965
rect 216029 135960 217212 135962
rect 216029 135904 216034 135960
rect 216090 135904 217212 135960
rect 216029 135902 217212 135904
rect 228804 135960 231275 135962
rect 228804 135904 231214 135960
rect 231270 135904 231275 135960
rect 228804 135902 231275 135904
rect 216029 135899 216095 135902
rect 231209 135899 231275 135902
rect 264973 135690 265039 135693
rect 264973 135688 268180 135690
rect 264973 135632 264978 135688
rect 265034 135632 268180 135688
rect 264973 135630 268180 135632
rect 264973 135627 265039 135630
rect 282361 135554 282427 135557
rect 279956 135552 282427 135554
rect 279956 135496 282366 135552
rect 282422 135496 282427 135552
rect 279956 135494 282427 135496
rect 282361 135491 282427 135494
rect 231393 135418 231459 135421
rect 228804 135416 231459 135418
rect 228804 135360 231398 135416
rect 231454 135360 231459 135416
rect 228804 135358 231459 135360
rect 231393 135355 231459 135358
rect 213913 135282 213979 135285
rect 264329 135282 264395 135285
rect 213913 135280 217212 135282
rect 213913 135224 213918 135280
rect 213974 135224 217212 135280
rect 213913 135222 217212 135224
rect 264329 135280 268180 135282
rect 264329 135224 264334 135280
rect 264390 135224 268180 135280
rect 264329 135222 268180 135224
rect 213913 135219 213979 135222
rect 264329 135219 264395 135222
rect 231761 135010 231827 135013
rect 228804 135008 231827 135010
rect 228804 134952 231766 135008
rect 231822 134952 231827 135008
rect 228804 134950 231827 134952
rect 231761 134947 231827 134950
rect 265157 134874 265223 134877
rect 265157 134872 268180 134874
rect 265157 134816 265162 134872
rect 265218 134816 268180 134872
rect 265157 134814 268180 134816
rect 265157 134811 265223 134814
rect 213913 134602 213979 134605
rect 213913 134600 217212 134602
rect 213913 134544 213918 134600
rect 213974 134544 217212 134600
rect 213913 134542 217212 134544
rect 213913 134539 213979 134542
rect 231669 134466 231735 134469
rect 228804 134464 231735 134466
rect 228804 134408 231674 134464
rect 231730 134408 231735 134464
rect 228804 134406 231735 134408
rect 231669 134403 231735 134406
rect 265065 134466 265131 134469
rect 265065 134464 268180 134466
rect 265065 134408 265070 134464
rect 265126 134408 268180 134464
rect 265065 134406 268180 134408
rect 265065 134403 265131 134406
rect 279926 134194 279986 134708
rect 288566 134194 288572 134196
rect 279926 134134 288572 134194
rect 288566 134132 288572 134134
rect 288636 134132 288642 134196
rect 231025 134058 231091 134061
rect 228804 134056 231091 134058
rect 228804 134000 231030 134056
rect 231086 134000 231091 134056
rect 228804 133998 231091 134000
rect 231025 133995 231091 133998
rect 264973 134058 265039 134061
rect 280102 134058 280108 134060
rect 264973 134056 268180 134058
rect 264973 134000 264978 134056
rect 265034 134000 268180 134056
rect 264973 133998 268180 134000
rect 279956 133998 280108 134058
rect 264973 133995 265039 133998
rect 280102 133996 280108 133998
rect 280172 133996 280178 134060
rect 213361 133922 213427 133925
rect 213361 133920 217212 133922
rect 213361 133864 213366 133920
rect 213422 133864 217212 133920
rect 213361 133862 217212 133864
rect 213361 133859 213427 133862
rect 264973 133650 265039 133653
rect 264973 133648 268180 133650
rect 264973 133592 264978 133648
rect 265034 133592 268180 133648
rect 264973 133590 268180 133592
rect 264973 133587 265039 133590
rect 231761 133514 231827 133517
rect 228804 133512 231827 133514
rect 228804 133456 231766 133512
rect 231822 133456 231827 133512
rect 228804 133454 231827 133456
rect 231761 133451 231827 133454
rect 214005 133378 214071 133381
rect 214005 133376 217212 133378
rect 214005 133320 214010 133376
rect 214066 133320 217212 133376
rect 214005 133318 217212 133320
rect 214005 133315 214071 133318
rect 283097 133242 283163 133245
rect 279956 133240 283163 133242
rect 279956 133184 283102 133240
rect 283158 133184 283163 133240
rect 279956 133182 283163 133184
rect 283097 133179 283163 133182
rect 231117 133106 231183 133109
rect 228804 133104 231183 133106
rect 228804 133048 231122 133104
rect 231178 133048 231183 133104
rect 228804 133046 231183 133048
rect 231117 133043 231183 133046
rect 265065 133106 265131 133109
rect 265065 133104 268180 133106
rect 265065 133048 265070 133104
rect 265126 133048 268180 133104
rect 265065 133046 268180 133048
rect 265065 133043 265131 133046
rect 213913 132698 213979 132701
rect 265617 132698 265683 132701
rect 213913 132696 217212 132698
rect 213913 132640 213918 132696
rect 213974 132640 217212 132696
rect 213913 132638 217212 132640
rect 265617 132696 268180 132698
rect 265617 132640 265622 132696
rect 265678 132640 268180 132696
rect 265617 132638 268180 132640
rect 213913 132635 213979 132638
rect 265617 132635 265683 132638
rect 231669 132562 231735 132565
rect 228804 132560 231735 132562
rect 228804 132504 231674 132560
rect 231730 132504 231735 132560
rect 228804 132502 231735 132504
rect 231669 132499 231735 132502
rect 282821 132426 282887 132429
rect 279956 132424 282887 132426
rect 279956 132368 282826 132424
rect 282882 132368 282887 132424
rect 279956 132366 282887 132368
rect 282821 132363 282887 132366
rect 231761 132154 231827 132157
rect 228804 132152 231827 132154
rect 228804 132096 231766 132152
rect 231822 132096 231827 132152
rect 228804 132094 231827 132096
rect 231761 132091 231827 132094
rect 214649 132018 214715 132021
rect 214649 132016 217212 132018
rect 214649 131960 214654 132016
rect 214710 131960 217212 132016
rect 214649 131958 217212 131960
rect 214649 131955 214715 131958
rect 244774 131956 244780 132020
rect 244844 132018 244850 132020
rect 268150 132018 268210 132260
rect 244844 131958 268210 132018
rect 244844 131956 244850 131958
rect 231669 131610 231735 131613
rect 228804 131608 231735 131610
rect 228804 131552 231674 131608
rect 231730 131552 231735 131608
rect 228804 131550 231735 131552
rect 231669 131547 231735 131550
rect 232446 131548 232452 131612
rect 232516 131610 232522 131612
rect 268150 131610 268210 131852
rect 282729 131746 282795 131749
rect 279956 131744 282795 131746
rect 279956 131688 282734 131744
rect 282790 131688 282795 131744
rect 279956 131686 282795 131688
rect 282729 131683 282795 131686
rect 232516 131550 268210 131610
rect 232516 131548 232522 131550
rect 267089 131474 267155 131477
rect 267089 131472 268180 131474
rect 267089 131416 267094 131472
rect 267150 131416 268180 131472
rect 267089 131414 268180 131416
rect 267089 131411 267155 131414
rect 213913 131338 213979 131341
rect 213913 131336 217212 131338
rect 213913 131280 213918 131336
rect 213974 131280 217212 131336
rect 213913 131278 217212 131280
rect 213913 131275 213979 131278
rect 231301 131202 231367 131205
rect 228804 131200 231367 131202
rect 228804 131144 231306 131200
rect 231362 131144 231367 131200
rect 228804 131142 231367 131144
rect 231301 131139 231367 131142
rect 267181 131066 267247 131069
rect 267181 131064 268180 131066
rect 267181 131008 267186 131064
rect 267242 131008 268180 131064
rect 267181 131006 268180 131008
rect 267181 131003 267247 131006
rect 282821 130930 282887 130933
rect 279956 130928 282887 130930
rect 279956 130872 282826 130928
rect 282882 130872 282887 130928
rect 279956 130870 282887 130872
rect 282821 130867 282887 130870
rect 213913 130658 213979 130661
rect 231761 130658 231827 130661
rect 213913 130656 217212 130658
rect 213913 130600 213918 130656
rect 213974 130600 217212 130656
rect 213913 130598 217212 130600
rect 228804 130656 231827 130658
rect 228804 130600 231766 130656
rect 231822 130600 231827 130656
rect 228804 130598 231827 130600
rect 213913 130595 213979 130598
rect 231761 130595 231827 130598
rect 265065 130522 265131 130525
rect 265065 130520 268180 130522
rect 265065 130464 265070 130520
rect 265126 130464 268180 130520
rect 265065 130462 268180 130464
rect 265065 130459 265131 130462
rect 231669 130250 231735 130253
rect 228804 130248 231735 130250
rect 228804 130192 231674 130248
rect 231730 130192 231735 130248
rect 228804 130190 231735 130192
rect 231669 130187 231735 130190
rect 264973 130114 265039 130117
rect 282177 130114 282243 130117
rect 264973 130112 268180 130114
rect 264973 130056 264978 130112
rect 265034 130056 268180 130112
rect 264973 130054 268180 130056
rect 279956 130112 282243 130114
rect 279956 130056 282182 130112
rect 282238 130056 282243 130112
rect 279956 130054 282243 130056
rect 264973 130051 265039 130054
rect 282177 130051 282243 130054
rect 214005 129978 214071 129981
rect 214005 129976 217212 129978
rect 214005 129920 214010 129976
rect 214066 129920 217212 129976
rect 214005 129918 217212 129920
rect 214005 129915 214071 129918
rect 231577 129842 231643 129845
rect 228804 129840 231643 129842
rect 228804 129784 231582 129840
rect 231638 129784 231643 129840
rect 228804 129782 231643 129784
rect 231577 129779 231643 129782
rect 265065 129706 265131 129709
rect 265065 129704 268180 129706
rect 265065 129648 265070 129704
rect 265126 129648 268180 129704
rect 265065 129646 268180 129648
rect 265065 129643 265131 129646
rect 280470 129434 280476 129436
rect 279956 129374 280476 129434
rect 280470 129372 280476 129374
rect 280540 129372 280546 129436
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 214005 129298 214071 129301
rect 231761 129298 231827 129301
rect 214005 129296 217212 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 214005 129240 214010 129296
rect 214066 129240 217212 129296
rect 214005 129238 217212 129240
rect 228804 129296 231827 129298
rect 228804 129240 231766 129296
rect 231822 129240 231827 129296
rect 228804 129238 231827 129240
rect 66161 129235 66227 129238
rect 214005 129235 214071 129238
rect 231761 129235 231827 129238
rect 264973 129298 265039 129301
rect 264973 129296 268180 129298
rect 264973 129240 264978 129296
rect 265034 129240 268180 129296
rect 264973 129238 268180 129240
rect 264973 129235 265039 129238
rect 231669 128890 231735 128893
rect 228804 128888 231735 128890
rect 228804 128832 231674 128888
rect 231730 128832 231735 128888
rect 228804 128830 231735 128832
rect 231669 128827 231735 128830
rect 258574 128828 258580 128892
rect 258644 128890 258650 128892
rect 258644 128830 268180 128890
rect 258644 128828 258650 128830
rect 213913 128754 213979 128757
rect 213913 128752 217212 128754
rect 213913 128696 213918 128752
rect 213974 128696 217212 128752
rect 213913 128694 217212 128696
rect 213913 128691 213979 128694
rect 282821 128618 282887 128621
rect 279956 128616 282887 128618
rect 279956 128560 282826 128616
rect 282882 128560 282887 128616
rect 279956 128558 282887 128560
rect 282821 128555 282887 128558
rect 267774 128420 267780 128484
rect 267844 128482 267850 128484
rect 267844 128422 268180 128482
rect 267844 128420 267850 128422
rect 231761 128346 231827 128349
rect 228804 128344 231827 128346
rect 228804 128288 231766 128344
rect 231822 128288 231827 128344
rect 228804 128286 231827 128288
rect 231761 128283 231827 128286
rect 66069 128074 66135 128077
rect 68142 128074 68816 128080
rect 66069 128072 68816 128074
rect 66069 128016 66074 128072
rect 66130 128020 68816 128072
rect 214005 128074 214071 128077
rect 214005 128072 217212 128074
rect 66130 128016 68202 128020
rect 66069 128014 68202 128016
rect 214005 128016 214010 128072
rect 214066 128016 217212 128072
rect 214005 128014 217212 128016
rect 66069 128011 66135 128014
rect 214005 128011 214071 128014
rect 230841 127938 230907 127941
rect 228804 127936 230907 127938
rect 228804 127880 230846 127936
rect 230902 127880 230907 127936
rect 228804 127878 230907 127880
rect 230841 127875 230907 127878
rect 267590 127876 267596 127940
rect 267660 127938 267666 127940
rect 267660 127878 268180 127938
rect 267660 127876 267666 127878
rect 281717 127802 281783 127805
rect 279956 127800 281783 127802
rect 279956 127744 281722 127800
rect 281778 127744 281783 127800
rect 279956 127742 281783 127744
rect 281717 127739 281783 127742
rect 265801 127530 265867 127533
rect 265801 127528 268180 127530
rect 265801 127472 265806 127528
rect 265862 127472 268180 127528
rect 265801 127470 268180 127472
rect 265801 127467 265867 127470
rect 213913 127394 213979 127397
rect 230974 127394 230980 127396
rect 213913 127392 217212 127394
rect 213913 127336 213918 127392
rect 213974 127336 217212 127392
rect 213913 127334 217212 127336
rect 228804 127334 230980 127394
rect 213913 127331 213979 127334
rect 230974 127332 230980 127334
rect 231044 127332 231050 127396
rect 264973 127122 265039 127125
rect 282821 127122 282887 127125
rect 264973 127120 268180 127122
rect 264973 127064 264978 127120
rect 265034 127064 268180 127120
rect 264973 127062 268180 127064
rect 279956 127120 282887 127122
rect 279956 127064 282826 127120
rect 282882 127064 282887 127120
rect 279956 127062 282887 127064
rect 264973 127059 265039 127062
rect 282821 127059 282887 127062
rect 231761 126986 231827 126989
rect 228804 126984 231827 126986
rect 228804 126928 231766 126984
rect 231822 126928 231827 126984
rect 228804 126926 231827 126928
rect 231761 126923 231827 126926
rect 214005 126714 214071 126717
rect 265157 126714 265223 126717
rect 214005 126712 217212 126714
rect 214005 126656 214010 126712
rect 214066 126656 217212 126712
rect 214005 126654 217212 126656
rect 265157 126712 268180 126714
rect 265157 126656 265162 126712
rect 265218 126656 268180 126712
rect 265157 126654 268180 126656
rect 214005 126651 214071 126654
rect 265157 126651 265223 126654
rect 583569 126578 583635 126581
rect 583526 126576 583635 126578
rect 583526 126520 583574 126576
rect 583630 126520 583635 126576
rect 583526 126515 583635 126520
rect 231669 126442 231735 126445
rect 228804 126440 231735 126442
rect 228804 126384 231674 126440
rect 231730 126384 231735 126440
rect 228804 126382 231735 126384
rect 231669 126379 231735 126382
rect 67449 126306 67515 126309
rect 68142 126306 68816 126312
rect 67449 126304 68816 126306
rect 67449 126248 67454 126304
rect 67510 126252 68816 126304
rect 265065 126306 265131 126309
rect 281901 126306 281967 126309
rect 265065 126304 268180 126306
rect 67510 126248 68202 126252
rect 67449 126246 68202 126248
rect 265065 126248 265070 126304
rect 265126 126248 268180 126304
rect 265065 126246 268180 126248
rect 279956 126304 281967 126306
rect 279956 126248 281906 126304
rect 281962 126248 281967 126304
rect 279956 126246 281967 126248
rect 67449 126243 67515 126246
rect 265065 126243 265131 126246
rect 281901 126243 281967 126246
rect 583526 126170 583586 126515
rect 583342 126124 583586 126170
rect 583342 126110 584960 126124
rect 213913 126034 213979 126037
rect 231117 126034 231183 126037
rect 213913 126032 217212 126034
rect 213913 125976 213918 126032
rect 213974 125976 217212 126032
rect 213913 125974 217212 125976
rect 228804 126032 231183 126034
rect 228804 125976 231122 126032
rect 231178 125976 231183 126032
rect 228804 125974 231183 125976
rect 583342 126034 583402 126110
rect 583520 126034 584960 126110
rect 583342 125974 584960 126034
rect 213913 125971 213979 125974
rect 231117 125971 231183 125974
rect 264973 125898 265039 125901
rect 264973 125896 268180 125898
rect 264973 125840 264978 125896
rect 265034 125840 268180 125896
rect 583520 125884 584960 125974
rect 264973 125838 268180 125840
rect 264973 125835 265039 125838
rect 231761 125490 231827 125493
rect 282821 125490 282887 125493
rect 228804 125488 231827 125490
rect 228804 125432 231766 125488
rect 231822 125432 231827 125488
rect 228804 125430 231827 125432
rect 279956 125488 282887 125490
rect 279956 125432 282826 125488
rect 282882 125432 282887 125488
rect 279956 125430 282887 125432
rect 231761 125427 231827 125430
rect 282821 125427 282887 125430
rect 214005 125354 214071 125357
rect 265157 125354 265223 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 265157 125352 268180 125354
rect 265157 125296 265162 125352
rect 265218 125296 268180 125352
rect 265157 125294 268180 125296
rect 214005 125291 214071 125294
rect 265157 125291 265223 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect 231761 125082 231827 125085
rect 228804 125080 231827 125082
rect 228804 125024 231766 125080
rect 231822 125024 231827 125080
rect 228804 125022 231827 125024
rect 231761 125019 231827 125022
rect 265065 124946 265131 124949
rect 265065 124944 268180 124946
rect 265065 124888 265070 124944
rect 265126 124888 268180 124944
rect 265065 124886 268180 124888
rect 265065 124883 265131 124886
rect 282729 124810 282795 124813
rect 279956 124808 282795 124810
rect 279956 124752 282734 124808
rect 282790 124752 282795 124808
rect 279956 124750 282795 124752
rect 282729 124747 282795 124750
rect 213913 124674 213979 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 213913 124611 213979 124614
rect 231485 124538 231551 124541
rect 228804 124536 231551 124538
rect 228804 124480 231490 124536
rect 231546 124480 231551 124536
rect 228804 124478 231551 124480
rect 231485 124475 231551 124478
rect 264973 124538 265039 124541
rect 264973 124536 268180 124538
rect 264973 124480 264978 124536
rect 265034 124480 268180 124536
rect 264973 124478 268180 124480
rect 264973 124475 265039 124478
rect 214005 124130 214071 124133
rect 230749 124130 230815 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 228804 124128 230815 124130
rect 228804 124072 230754 124128
rect 230810 124072 230815 124128
rect 228804 124070 230815 124072
rect 214005 124067 214071 124070
rect 230749 124067 230815 124070
rect 265157 124130 265223 124133
rect 265157 124128 268180 124130
rect 265157 124072 265162 124128
rect 265218 124072 268180 124128
rect 265157 124070 268180 124072
rect 265157 124067 265223 124070
rect 282821 123994 282887 123997
rect 279956 123992 282887 123994
rect 279956 123936 282826 123992
rect 282882 123936 282887 123992
rect 279956 123934 282887 123936
rect 282821 123931 282887 123934
rect -960 123572 480 123812
rect 265065 123722 265131 123725
rect 265065 123720 268180 123722
rect 265065 123664 265070 123720
rect 265126 123664 268180 123720
rect 265065 123662 268180 123664
rect 265065 123659 265131 123662
rect 67541 123586 67607 123589
rect 68142 123586 68816 123592
rect 230933 123586 230999 123589
rect 67541 123584 68816 123586
rect 67541 123528 67546 123584
rect 67602 123532 68816 123584
rect 228804 123584 230999 123586
rect 67602 123528 68202 123532
rect 67541 123526 68202 123528
rect 228804 123528 230938 123584
rect 230994 123528 230999 123584
rect 228804 123526 230999 123528
rect 67541 123523 67607 123526
rect 230933 123523 230999 123526
rect 213913 123450 213979 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 213913 123387 213979 123390
rect 264973 123314 265039 123317
rect 264973 123312 268180 123314
rect 264973 123256 264978 123312
rect 265034 123256 268180 123312
rect 264973 123254 268180 123256
rect 264973 123251 265039 123254
rect 231577 123178 231643 123181
rect 282637 123178 282703 123181
rect 228804 123176 231643 123178
rect 228804 123120 231582 123176
rect 231638 123120 231643 123176
rect 228804 123118 231643 123120
rect 279956 123176 282703 123178
rect 279956 123120 282642 123176
rect 282698 123120 282703 123176
rect 279956 123118 282703 123120
rect 231577 123115 231643 123118
rect 282637 123115 282703 123118
rect 265709 122906 265775 122909
rect 265709 122904 268180 122906
rect 265709 122848 265714 122904
rect 265770 122848 268180 122904
rect 265709 122846 268180 122848
rect 265709 122843 265775 122846
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 65977 122634 66043 122637
rect 68142 122634 68816 122640
rect 231761 122634 231827 122637
rect 65977 122632 68816 122634
rect 65977 122576 65982 122632
rect 66038 122580 68816 122632
rect 228804 122632 231827 122634
rect 66038 122576 68202 122580
rect 65977 122574 68202 122576
rect 228804 122576 231766 122632
rect 231822 122576 231827 122632
rect 228804 122574 231827 122576
rect 65977 122571 66043 122574
rect 231761 122571 231827 122574
rect 265065 122362 265131 122365
rect 265065 122360 268180 122362
rect 265065 122304 265070 122360
rect 265126 122304 268180 122360
rect 265065 122302 268180 122304
rect 265065 122299 265131 122302
rect 231669 122226 231735 122229
rect 228804 122224 231735 122226
rect 228804 122168 231674 122224
rect 231730 122168 231735 122224
rect 228804 122166 231735 122168
rect 231669 122163 231735 122166
rect 213913 122090 213979 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 213913 122027 213979 122030
rect 265157 121954 265223 121957
rect 265157 121952 268180 121954
rect 265157 121896 265162 121952
rect 265218 121896 268180 121952
rect 265157 121894 268180 121896
rect 265157 121891 265223 121894
rect 279926 121818 279986 122468
rect 287094 121818 287100 121820
rect 279926 121758 287100 121818
rect 287094 121756 287100 121758
rect 287164 121756 287170 121820
rect 230749 121682 230815 121685
rect 282821 121682 282887 121685
rect 228804 121680 230815 121682
rect 228804 121624 230754 121680
rect 230810 121624 230815 121680
rect 228804 121622 230815 121624
rect 279956 121680 282887 121682
rect 279956 121624 282826 121680
rect 282882 121624 282887 121680
rect 279956 121622 282887 121624
rect 230749 121619 230815 121622
rect 282821 121619 282887 121622
rect 264973 121546 265039 121549
rect 264973 121544 268180 121546
rect 264973 121488 264978 121544
rect 265034 121488 268180 121544
rect 264973 121486 268180 121488
rect 264973 121483 265039 121486
rect 214005 121410 214071 121413
rect 214005 121408 217212 121410
rect 214005 121352 214010 121408
rect 214066 121352 217212 121408
rect 214005 121350 217212 121352
rect 214005 121347 214071 121350
rect 231761 121274 231827 121277
rect 228804 121272 231827 121274
rect 228804 121216 231766 121272
rect 231822 121216 231827 121272
rect 228804 121214 231827 121216
rect 231761 121211 231827 121214
rect 265157 121138 265223 121141
rect 265157 121136 268180 121138
rect 265157 121080 265162 121136
rect 265218 121080 268180 121136
rect 265157 121078 268180 121080
rect 265157 121075 265223 121078
rect 65885 120866 65951 120869
rect 68142 120866 68816 120872
rect 281533 120866 281599 120869
rect 65885 120864 68816 120866
rect 65885 120808 65890 120864
rect 65946 120812 68816 120864
rect 279956 120864 281599 120866
rect 65946 120808 68202 120812
rect 65885 120806 68202 120808
rect 279956 120808 281538 120864
rect 281594 120808 281599 120864
rect 279956 120806 281599 120808
rect 65885 120803 65951 120806
rect 281533 120803 281599 120806
rect 213913 120730 213979 120733
rect 231577 120730 231643 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 228804 120728 231643 120730
rect 228804 120672 231582 120728
rect 231638 120672 231643 120728
rect 228804 120670 231643 120672
rect 213913 120667 213979 120670
rect 231577 120667 231643 120670
rect 264973 120730 265039 120733
rect 264973 120728 268180 120730
rect 264973 120672 264978 120728
rect 265034 120672 268180 120728
rect 264973 120670 268180 120672
rect 264973 120667 265039 120670
rect 231669 120322 231735 120325
rect 228804 120320 231735 120322
rect 228804 120264 231674 120320
rect 231730 120264 231735 120320
rect 228804 120262 231735 120264
rect 231669 120259 231735 120262
rect 265065 120322 265131 120325
rect 265065 120320 268180 120322
rect 265065 120264 265070 120320
rect 265126 120264 268180 120320
rect 265065 120262 268180 120264
rect 265065 120259 265131 120262
rect 282729 120186 282795 120189
rect 279956 120184 282795 120186
rect 279956 120128 282734 120184
rect 282790 120128 282795 120184
rect 279956 120126 282795 120128
rect 282729 120123 282795 120126
rect 214097 120050 214163 120053
rect 214097 120048 217212 120050
rect 214097 119992 214102 120048
rect 214158 119992 217212 120048
rect 214097 119990 217212 119992
rect 214097 119987 214163 119990
rect 230933 119778 230999 119781
rect 228804 119776 230999 119778
rect 228804 119720 230938 119776
rect 230994 119720 230999 119776
rect 228804 119718 230999 119720
rect 230933 119715 230999 119718
rect 264973 119778 265039 119781
rect 264973 119776 268180 119778
rect 264973 119720 264978 119776
rect 265034 119720 268180 119776
rect 264973 119718 268180 119720
rect 264973 119715 265039 119718
rect 214005 119506 214071 119509
rect 214005 119504 217212 119506
rect 214005 119448 214010 119504
rect 214066 119448 217212 119504
rect 214005 119446 217212 119448
rect 214005 119443 214071 119446
rect 231393 119370 231459 119373
rect 282085 119370 282151 119373
rect 228804 119368 231459 119370
rect 228804 119312 231398 119368
rect 231454 119312 231459 119368
rect 279956 119368 282151 119370
rect 228804 119310 231459 119312
rect 231393 119307 231459 119310
rect 251766 119036 251772 119100
rect 251836 119098 251842 119100
rect 268150 119098 268210 119340
rect 279956 119312 282090 119368
rect 282146 119312 282151 119368
rect 279956 119310 282151 119312
rect 282085 119307 282151 119310
rect 251836 119038 268210 119098
rect 251836 119036 251842 119038
rect 230749 118962 230815 118965
rect 228804 118960 230815 118962
rect 228804 118904 230754 118960
rect 230810 118904 230815 118960
rect 228804 118902 230815 118904
rect 230749 118899 230815 118902
rect 264237 118962 264303 118965
rect 264237 118960 268180 118962
rect 264237 118904 264242 118960
rect 264298 118904 268180 118960
rect 264237 118902 268180 118904
rect 264237 118899 264303 118902
rect 213913 118826 213979 118829
rect 213913 118824 217212 118826
rect 213913 118768 213918 118824
rect 213974 118768 217212 118824
rect 213913 118766 217212 118768
rect 213913 118763 213979 118766
rect 264973 118554 265039 118557
rect 282821 118554 282887 118557
rect 264973 118552 268180 118554
rect 264973 118496 264978 118552
rect 265034 118496 268180 118552
rect 264973 118494 268180 118496
rect 279956 118552 282887 118554
rect 279956 118496 282826 118552
rect 282882 118496 282887 118552
rect 279956 118494 282887 118496
rect 264973 118491 265039 118494
rect 282821 118491 282887 118494
rect 231669 118418 231735 118421
rect 228804 118416 231735 118418
rect 228804 118360 231674 118416
rect 231730 118360 231735 118416
rect 228804 118358 231735 118360
rect 231669 118355 231735 118358
rect 214005 118146 214071 118149
rect 266997 118146 267063 118149
rect 214005 118144 217212 118146
rect 214005 118088 214010 118144
rect 214066 118088 217212 118144
rect 214005 118086 217212 118088
rect 266997 118144 268180 118146
rect 266997 118088 267002 118144
rect 267058 118088 268180 118144
rect 266997 118086 268180 118088
rect 214005 118083 214071 118086
rect 266997 118083 267063 118086
rect 231761 118010 231827 118013
rect 228804 118008 231827 118010
rect 228804 117952 231766 118008
rect 231822 117952 231827 118008
rect 228804 117950 231827 117952
rect 231761 117947 231827 117950
rect 282729 117874 282795 117877
rect 279956 117872 282795 117874
rect 279956 117816 282734 117872
rect 282790 117816 282795 117872
rect 279956 117814 282795 117816
rect 282729 117811 282795 117814
rect 265065 117738 265131 117741
rect 265065 117736 268180 117738
rect 265065 117680 265070 117736
rect 265126 117680 268180 117736
rect 265065 117678 268180 117680
rect 265065 117675 265131 117678
rect 213913 117466 213979 117469
rect 231485 117466 231551 117469
rect 213913 117464 217212 117466
rect 213913 117408 213918 117464
rect 213974 117408 217212 117464
rect 213913 117406 217212 117408
rect 228804 117464 231551 117466
rect 228804 117408 231490 117464
rect 231546 117408 231551 117464
rect 228804 117406 231551 117408
rect 213913 117403 213979 117406
rect 231485 117403 231551 117406
rect 265157 117194 265223 117197
rect 265157 117192 268180 117194
rect 265157 117136 265162 117192
rect 265218 117136 268180 117192
rect 265157 117134 268180 117136
rect 265157 117131 265223 117134
rect 231761 117058 231827 117061
rect 282821 117058 282887 117061
rect 228804 117056 231827 117058
rect 228804 117000 231766 117056
rect 231822 117000 231827 117056
rect 228804 116998 231827 117000
rect 279956 117056 282887 117058
rect 279956 117000 282826 117056
rect 282882 117000 282887 117056
rect 279956 116998 282887 117000
rect 231761 116995 231827 116998
rect 282821 116995 282887 116998
rect 213913 116786 213979 116789
rect 264973 116786 265039 116789
rect 213913 116784 217212 116786
rect 213913 116728 213918 116784
rect 213974 116728 217212 116784
rect 213913 116726 217212 116728
rect 264973 116784 268180 116786
rect 264973 116728 264978 116784
rect 265034 116728 268180 116784
rect 264973 116726 268180 116728
rect 213913 116723 213979 116726
rect 264973 116723 265039 116726
rect 230974 116588 230980 116652
rect 231044 116650 231050 116652
rect 265801 116650 265867 116653
rect 231044 116648 265867 116650
rect 231044 116592 265806 116648
rect 265862 116592 265867 116648
rect 231044 116590 265867 116592
rect 231044 116588 231050 116590
rect 265801 116587 265867 116590
rect 231209 116514 231275 116517
rect 228804 116512 231275 116514
rect 228804 116456 231214 116512
rect 231270 116456 231275 116512
rect 228804 116454 231275 116456
rect 231209 116451 231275 116454
rect 265065 116378 265131 116381
rect 282729 116378 282795 116381
rect 265065 116376 268180 116378
rect 265065 116320 265070 116376
rect 265126 116320 268180 116376
rect 265065 116318 268180 116320
rect 279956 116376 282795 116378
rect 279956 116320 282734 116376
rect 282790 116320 282795 116376
rect 279956 116318 282795 116320
rect 265065 116315 265131 116318
rect 282729 116315 282795 116318
rect 216213 116106 216279 116109
rect 230657 116106 230723 116109
rect 216213 116104 217212 116106
rect 216213 116048 216218 116104
rect 216274 116048 217212 116104
rect 216213 116046 217212 116048
rect 228804 116104 230723 116106
rect 228804 116048 230662 116104
rect 230718 116048 230723 116104
rect 228804 116046 230723 116048
rect 216213 116043 216279 116046
rect 230657 116043 230723 116046
rect 264973 115970 265039 115973
rect 264973 115968 268180 115970
rect 264973 115912 264978 115968
rect 265034 115912 268180 115968
rect 264973 115910 268180 115912
rect 264973 115907 265039 115910
rect 231761 115562 231827 115565
rect 228804 115560 231827 115562
rect 228804 115504 231766 115560
rect 231822 115504 231827 115560
rect 228804 115502 231827 115504
rect 231761 115499 231827 115502
rect 264973 115562 265039 115565
rect 282085 115562 282151 115565
rect 264973 115560 268180 115562
rect 264973 115504 264978 115560
rect 265034 115504 268180 115560
rect 264973 115502 268180 115504
rect 279956 115560 282151 115562
rect 279956 115504 282090 115560
rect 282146 115504 282151 115560
rect 279956 115502 282151 115504
rect 264973 115499 265039 115502
rect 282085 115499 282151 115502
rect 214005 115426 214071 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 214005 115363 214071 115366
rect 231158 115154 231164 115156
rect 228804 115094 231164 115154
rect 231158 115092 231164 115094
rect 231228 115092 231234 115156
rect 262806 115092 262812 115156
rect 262876 115154 262882 115156
rect 262876 115094 268180 115154
rect 262876 115092 262882 115094
rect 213913 114882 213979 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 213913 114819 213979 114822
rect 281717 114746 281783 114749
rect 279956 114744 281783 114746
rect 279956 114688 281722 114744
rect 281778 114688 281783 114744
rect 279956 114686 281783 114688
rect 281717 114683 281783 114686
rect 231669 114610 231735 114613
rect 228804 114608 231735 114610
rect 228804 114552 231674 114608
rect 231730 114552 231735 114608
rect 228804 114550 231735 114552
rect 231669 114547 231735 114550
rect 265801 114610 265867 114613
rect 265801 114608 268180 114610
rect 265801 114552 265806 114608
rect 265862 114552 268180 114608
rect 265801 114550 268180 114552
rect 265801 114547 265867 114550
rect 234061 114474 234127 114477
rect 237414 114474 237420 114476
rect 234061 114472 237420 114474
rect 234061 114416 234066 114472
rect 234122 114416 237420 114472
rect 234061 114414 237420 114416
rect 234061 114411 234127 114414
rect 237414 114412 237420 114414
rect 237484 114412 237490 114476
rect 214005 114202 214071 114205
rect 231761 114202 231827 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 228804 114200 231827 114202
rect 228804 114144 231766 114200
rect 231822 114144 231827 114200
rect 228804 114142 231827 114144
rect 214005 114139 214071 114142
rect 231761 114139 231827 114142
rect 253054 113868 253060 113932
rect 253124 113930 253130 113932
rect 268150 113930 268210 114172
rect 282821 114066 282887 114069
rect 279956 114064 282887 114066
rect 279956 114008 282826 114064
rect 282882 114008 282887 114064
rect 279956 114006 282887 114008
rect 282821 114003 282887 114006
rect 253124 113870 268210 113930
rect 253124 113868 253130 113870
rect 231485 113658 231551 113661
rect 228804 113656 231551 113658
rect 228804 113600 231490 113656
rect 231546 113600 231551 113656
rect 228804 113598 231551 113600
rect 231485 113595 231551 113598
rect 213913 113522 213979 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 213913 113459 213979 113462
rect 250294 113460 250300 113524
rect 250364 113522 250370 113524
rect 268150 113522 268210 113764
rect 250364 113462 268210 113522
rect 250364 113460 250370 113462
rect 267641 113386 267707 113389
rect 267641 113384 268180 113386
rect 267641 113328 267646 113384
rect 267702 113328 268180 113384
rect 267641 113326 268180 113328
rect 267641 113323 267707 113326
rect 229921 113250 229987 113253
rect 282729 113250 282795 113253
rect 228804 113248 229987 113250
rect 228804 113192 229926 113248
rect 229982 113192 229987 113248
rect 228804 113190 229987 113192
rect 279956 113248 282795 113250
rect 279956 113192 282734 113248
rect 282790 113192 282795 113248
rect 279956 113190 282795 113192
rect 229921 113187 229987 113190
rect 282729 113187 282795 113190
rect 265065 112978 265131 112981
rect 265065 112976 268180 112978
rect 265065 112920 265070 112976
rect 265126 112920 268180 112976
rect 265065 112918 268180 112920
rect 265065 112915 265131 112918
rect 214005 112842 214071 112845
rect 583017 112842 583083 112845
rect 583520 112842 584960 112932
rect 214005 112840 217212 112842
rect 214005 112784 214010 112840
rect 214066 112784 217212 112840
rect 214005 112782 217212 112784
rect 583017 112840 584960 112842
rect 583017 112784 583022 112840
rect 583078 112784 584960 112840
rect 583017 112782 584960 112784
rect 214005 112779 214071 112782
rect 583017 112779 583083 112782
rect 231761 112706 231827 112709
rect 228804 112704 231827 112706
rect 228804 112648 231766 112704
rect 231822 112648 231827 112704
rect 583520 112692 584960 112782
rect 228804 112646 231827 112648
rect 231761 112643 231827 112646
rect 264973 112570 265039 112573
rect 264973 112568 268180 112570
rect 264973 112512 264978 112568
rect 265034 112512 268180 112568
rect 264973 112510 268180 112512
rect 264973 112507 265039 112510
rect 282085 112434 282151 112437
rect 279956 112432 282151 112434
rect 279956 112376 282090 112432
rect 282146 112376 282151 112432
rect 279956 112374 282151 112376
rect 282085 112371 282151 112374
rect 231669 112298 231735 112301
rect 228804 112296 231735 112298
rect 228804 112240 231674 112296
rect 231730 112240 231735 112296
rect 228804 112238 231735 112240
rect 231669 112235 231735 112238
rect 213913 112162 213979 112165
rect 213913 112160 217212 112162
rect 213913 112104 213918 112160
rect 213974 112104 217212 112160
rect 213913 112102 217212 112104
rect 213913 112099 213979 112102
rect 265157 112026 265223 112029
rect 265157 112024 268180 112026
rect 265157 111968 265162 112024
rect 265218 111968 268180 112024
rect 265157 111966 268180 111968
rect 265157 111963 265223 111966
rect 164724 111754 165354 111760
rect 167821 111754 167887 111757
rect 231301 111754 231367 111757
rect 282821 111754 282887 111757
rect 164724 111752 167887 111754
rect 164724 111700 167826 111752
rect 165294 111696 167826 111700
rect 167882 111696 167887 111752
rect 165294 111694 167887 111696
rect 228804 111752 231367 111754
rect 228804 111696 231306 111752
rect 231362 111696 231367 111752
rect 228804 111694 231367 111696
rect 279956 111752 282887 111754
rect 279956 111696 282826 111752
rect 282882 111696 282887 111752
rect 279956 111694 282887 111696
rect 167821 111691 167887 111694
rect 231301 111691 231367 111694
rect 282821 111691 282887 111694
rect 265065 111618 265131 111621
rect 265065 111616 268180 111618
rect 265065 111560 265070 111616
rect 265126 111560 268180 111616
rect 265065 111558 268180 111560
rect 265065 111555 265131 111558
rect 214005 111482 214071 111485
rect 214005 111480 217212 111482
rect 214005 111424 214010 111480
rect 214066 111424 217212 111480
rect 214005 111422 217212 111424
rect 214005 111419 214071 111422
rect 231761 111346 231827 111349
rect 228804 111344 231827 111346
rect 228804 111288 231766 111344
rect 231822 111288 231827 111344
rect 228804 111286 231827 111288
rect 231761 111283 231827 111286
rect 265157 111210 265223 111213
rect 265157 111208 268180 111210
rect 265157 111152 265162 111208
rect 265218 111152 268180 111208
rect 265157 111150 268180 111152
rect 265157 111147 265223 111150
rect 282729 110938 282795 110941
rect 279956 110936 282795 110938
rect 279956 110880 282734 110936
rect 282790 110880 282795 110936
rect 279956 110878 282795 110880
rect 282729 110875 282795 110878
rect 213913 110802 213979 110805
rect 230565 110802 230631 110805
rect 213913 110800 217212 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217212 110800
rect 213913 110742 217212 110744
rect 228804 110800 230631 110802
rect 228804 110744 230570 110800
rect 230626 110744 230631 110800
rect 228804 110742 230631 110744
rect 213913 110739 213979 110742
rect 230565 110739 230631 110742
rect 264973 110802 265039 110805
rect 264973 110800 268180 110802
rect 264973 110744 264978 110800
rect 265034 110744 268180 110800
rect 264973 110742 268180 110744
rect 264973 110739 265039 110742
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 231761 110394 231827 110397
rect 228804 110392 231827 110394
rect 228804 110336 231766 110392
rect 231822 110336 231827 110392
rect 228804 110334 231827 110336
rect 231761 110331 231827 110334
rect 265065 110394 265131 110397
rect 265065 110392 268180 110394
rect 265065 110336 265070 110392
rect 265126 110336 268180 110392
rect 265065 110334 268180 110336
rect 265065 110331 265131 110334
rect 214005 110258 214071 110261
rect 214005 110256 217212 110258
rect 214005 110200 214010 110256
rect 214066 110200 217212 110256
rect 214005 110198 217212 110200
rect 214005 110195 214071 110198
rect 164724 110122 165354 110128
rect 167821 110122 167887 110125
rect 282085 110122 282151 110125
rect 164724 110120 167887 110122
rect 164724 110068 167826 110120
rect 165294 110064 167826 110068
rect 167882 110064 167887 110120
rect 165294 110062 167887 110064
rect 279956 110120 282151 110122
rect 279956 110064 282090 110120
rect 282146 110064 282151 110120
rect 279956 110062 282151 110064
rect 167821 110059 167887 110062
rect 282085 110059 282151 110062
rect 264973 109986 265039 109989
rect 264973 109984 268180 109986
rect 264973 109928 264978 109984
rect 265034 109928 268180 109984
rect 264973 109926 268180 109928
rect 264973 109923 265039 109926
rect 231669 109850 231735 109853
rect 228804 109848 231735 109850
rect 228804 109792 231674 109848
rect 231730 109792 231735 109848
rect 228804 109790 231735 109792
rect 231669 109787 231735 109790
rect 213913 109578 213979 109581
rect 265157 109578 265223 109581
rect 213913 109576 217212 109578
rect 213913 109520 213918 109576
rect 213974 109520 217212 109576
rect 213913 109518 217212 109520
rect 265157 109576 268180 109578
rect 265157 109520 265162 109576
rect 265218 109520 268180 109576
rect 265157 109518 268180 109520
rect 213913 109515 213979 109518
rect 265157 109515 265223 109518
rect 230565 109442 230631 109445
rect 282269 109442 282335 109445
rect 228804 109440 230631 109442
rect 228804 109384 230570 109440
rect 230626 109384 230631 109440
rect 228804 109382 230631 109384
rect 279956 109440 282335 109442
rect 279956 109384 282274 109440
rect 282330 109384 282335 109440
rect 279956 109382 282335 109384
rect 230565 109379 230631 109382
rect 282269 109379 282335 109382
rect 265157 109034 265223 109037
rect 265157 109032 268180 109034
rect 265157 108976 265162 109032
rect 265218 108976 268180 109032
rect 265157 108974 268180 108976
rect 265157 108971 265223 108974
rect 214005 108898 214071 108901
rect 231761 108898 231827 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 228804 108896 231827 108898
rect 228804 108840 231766 108896
rect 231822 108840 231827 108896
rect 228804 108838 231827 108840
rect 214005 108835 214071 108838
rect 231761 108835 231827 108838
rect 164724 108762 165354 108768
rect 167821 108762 167887 108765
rect 164724 108760 167887 108762
rect 164724 108708 167826 108760
rect 165294 108704 167826 108708
rect 167882 108704 167887 108760
rect 165294 108702 167887 108704
rect 167821 108699 167887 108702
rect 265065 108626 265131 108629
rect 282085 108626 282151 108629
rect 265065 108624 268180 108626
rect 265065 108568 265070 108624
rect 265126 108568 268180 108624
rect 265065 108566 268180 108568
rect 279956 108624 282151 108626
rect 279956 108568 282090 108624
rect 282146 108568 282151 108624
rect 279956 108566 282151 108568
rect 265065 108563 265131 108566
rect 282085 108563 282151 108566
rect 231485 108490 231551 108493
rect 228804 108488 231551 108490
rect 228804 108432 231490 108488
rect 231546 108432 231551 108488
rect 228804 108430 231551 108432
rect 231485 108427 231551 108430
rect 213913 108218 213979 108221
rect 264513 108218 264579 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 264513 108216 268180 108218
rect 264513 108160 264518 108216
rect 264574 108160 268180 108216
rect 264513 108158 268180 108160
rect 213913 108155 213979 108158
rect 264513 108155 264579 108158
rect 230841 107946 230907 107949
rect 228804 107944 230907 107946
rect 228804 107888 230846 107944
rect 230902 107888 230907 107944
rect 228804 107886 230907 107888
rect 230841 107883 230907 107886
rect 264973 107810 265039 107813
rect 281717 107810 281783 107813
rect 264973 107808 268180 107810
rect 264973 107752 264978 107808
rect 265034 107752 268180 107808
rect 264973 107750 268180 107752
rect 279956 107808 281783 107810
rect 279956 107752 281722 107808
rect 281778 107752 281783 107808
rect 279956 107750 281783 107752
rect 264973 107747 265039 107750
rect 281717 107747 281783 107750
rect 214005 107538 214071 107541
rect 231761 107538 231827 107541
rect 214005 107536 217212 107538
rect 214005 107480 214010 107536
rect 214066 107480 217212 107536
rect 214005 107478 217212 107480
rect 228804 107536 231827 107538
rect 228804 107480 231766 107536
rect 231822 107480 231827 107536
rect 228804 107478 231827 107480
rect 214005 107475 214071 107478
rect 231761 107475 231827 107478
rect 265065 107402 265131 107405
rect 265065 107400 268180 107402
rect 265065 107344 265070 107400
rect 265126 107344 268180 107400
rect 265065 107342 268180 107344
rect 265065 107339 265131 107342
rect 231301 107130 231367 107133
rect 228804 107128 231367 107130
rect 228804 107072 231306 107128
rect 231362 107072 231367 107128
rect 228804 107070 231367 107072
rect 231301 107067 231367 107070
rect 264973 106994 265039 106997
rect 264973 106992 268180 106994
rect 264973 106936 264978 106992
rect 265034 106936 268180 106992
rect 264973 106934 268180 106936
rect 264973 106931 265039 106934
rect 213913 106858 213979 106861
rect 213913 106856 217212 106858
rect 213913 106800 213918 106856
rect 213974 106800 217212 106856
rect 213913 106798 217212 106800
rect 213913 106795 213979 106798
rect 231485 106586 231551 106589
rect 228804 106584 231551 106586
rect 228804 106528 231490 106584
rect 231546 106528 231551 106584
rect 228804 106526 231551 106528
rect 231485 106523 231551 106526
rect 264421 106450 264487 106453
rect 279926 106450 279986 107100
rect 288382 106450 288388 106452
rect 264421 106448 268180 106450
rect 264421 106392 264426 106448
rect 264482 106392 268180 106448
rect 264421 106390 268180 106392
rect 279926 106390 288388 106450
rect 264421 106387 264487 106390
rect 288382 106388 288388 106390
rect 288452 106388 288458 106452
rect 287278 106314 287284 106316
rect 279956 106254 287284 106314
rect 287278 106252 287284 106254
rect 287348 106252 287354 106316
rect 214005 106178 214071 106181
rect 231761 106178 231827 106181
rect 214005 106176 217212 106178
rect 214005 106120 214010 106176
rect 214066 106120 217212 106176
rect 214005 106118 217212 106120
rect 228804 106176 231827 106178
rect 228804 106120 231766 106176
rect 231822 106120 231827 106176
rect 228804 106118 231827 106120
rect 214005 106115 214071 106118
rect 231761 106115 231827 106118
rect 265433 106042 265499 106045
rect 265433 106040 268180 106042
rect 265433 105984 265438 106040
rect 265494 105984 268180 106040
rect 265433 105982 268180 105984
rect 265433 105979 265499 105982
rect 215017 105634 215083 105637
rect 231669 105634 231735 105637
rect 215017 105632 217212 105634
rect 215017 105576 215022 105632
rect 215078 105576 217212 105632
rect 215017 105574 217212 105576
rect 228804 105632 231735 105634
rect 228804 105576 231674 105632
rect 231730 105576 231735 105632
rect 228804 105574 231735 105576
rect 215017 105571 215083 105574
rect 231669 105571 231735 105574
rect 264973 105634 265039 105637
rect 264973 105632 268180 105634
rect 264973 105576 264978 105632
rect 265034 105576 268180 105632
rect 264973 105574 268180 105576
rect 264973 105571 265039 105574
rect 281533 105498 281599 105501
rect 279956 105496 281599 105498
rect 279956 105440 281538 105496
rect 281594 105440 281599 105496
rect 279956 105438 281599 105440
rect 281533 105435 281599 105438
rect 230565 105226 230631 105229
rect 228804 105224 230631 105226
rect 228804 105168 230570 105224
rect 230626 105168 230631 105224
rect 228804 105166 230631 105168
rect 230565 105163 230631 105166
rect 265065 105226 265131 105229
rect 265065 105224 268180 105226
rect 265065 105168 265070 105224
rect 265126 105168 268180 105224
rect 265065 105166 268180 105168
rect 265065 105163 265131 105166
rect 213913 104954 213979 104957
rect 213913 104952 217212 104954
rect 213913 104896 213918 104952
rect 213974 104896 217212 104952
rect 213913 104894 217212 104896
rect 213913 104891 213979 104894
rect 265157 104818 265223 104821
rect 285806 104818 285812 104820
rect 265157 104816 268180 104818
rect 265157 104760 265162 104816
rect 265218 104760 268180 104816
rect 265157 104758 268180 104760
rect 279956 104758 285812 104818
rect 265157 104755 265223 104758
rect 285806 104756 285812 104758
rect 285876 104756 285882 104820
rect 231761 104682 231827 104685
rect 228804 104680 231827 104682
rect 228804 104624 231766 104680
rect 231822 104624 231827 104680
rect 228804 104622 231827 104624
rect 231761 104619 231827 104622
rect 265065 104410 265131 104413
rect 265065 104408 268180 104410
rect 265065 104352 265070 104408
rect 265126 104352 268180 104408
rect 265065 104350 268180 104352
rect 265065 104347 265131 104350
rect 214833 104274 214899 104277
rect 230841 104274 230907 104277
rect 214833 104272 217212 104274
rect 214833 104216 214838 104272
rect 214894 104216 217212 104272
rect 214833 104214 217212 104216
rect 228804 104272 230907 104274
rect 228804 104216 230846 104272
rect 230902 104216 230907 104272
rect 228804 104214 230907 104216
rect 214833 104211 214899 104214
rect 230841 104211 230907 104214
rect 282821 104002 282887 104005
rect 279956 104000 282887 104002
rect 279956 103944 282826 104000
rect 282882 103944 282887 104000
rect 279956 103942 282887 103944
rect 282821 103939 282887 103942
rect 264973 103866 265039 103869
rect 264973 103864 268180 103866
rect 264973 103808 264978 103864
rect 265034 103808 268180 103864
rect 264973 103806 268180 103808
rect 264973 103803 265039 103806
rect 231485 103730 231551 103733
rect 228804 103728 231551 103730
rect 228804 103672 231490 103728
rect 231546 103672 231551 103728
rect 228804 103670 231551 103672
rect 231485 103667 231551 103670
rect 213913 103594 213979 103597
rect 213913 103592 217212 103594
rect 213913 103536 213918 103592
rect 213974 103536 217212 103592
rect 213913 103534 217212 103536
rect 213913 103531 213979 103534
rect 265249 103458 265315 103461
rect 265249 103456 268180 103458
rect 265249 103400 265254 103456
rect 265310 103400 268180 103456
rect 265249 103398 268180 103400
rect 265249 103395 265315 103398
rect 231761 103322 231827 103325
rect 228804 103320 231827 103322
rect 228804 103264 231766 103320
rect 231822 103264 231827 103320
rect 228804 103262 231827 103264
rect 231761 103259 231827 103262
rect 265065 103050 265131 103053
rect 265065 103048 268180 103050
rect 265065 102992 265070 103048
rect 265126 102992 268180 103048
rect 265065 102990 268180 102992
rect 265065 102987 265131 102990
rect 213453 102914 213519 102917
rect 213453 102912 217212 102914
rect 213453 102856 213458 102912
rect 213514 102856 217212 102912
rect 213453 102854 217212 102856
rect 213453 102851 213519 102854
rect 166206 102716 166212 102780
rect 166276 102778 166282 102780
rect 214557 102778 214623 102781
rect 231669 102778 231735 102781
rect 166276 102776 214623 102778
rect 166276 102720 214562 102776
rect 214618 102720 214623 102776
rect 166276 102718 214623 102720
rect 228804 102776 231735 102778
rect 228804 102720 231674 102776
rect 231730 102720 231735 102776
rect 228804 102718 231735 102720
rect 166276 102716 166282 102718
rect 214557 102715 214623 102718
rect 231669 102715 231735 102718
rect 265157 102642 265223 102645
rect 279926 102642 279986 103156
rect 265157 102640 268180 102642
rect 265157 102584 265162 102640
rect 265218 102584 268180 102640
rect 265157 102582 268180 102584
rect 279926 102582 287070 102642
rect 265157 102579 265223 102582
rect 282821 102506 282887 102509
rect 279956 102504 282887 102506
rect 279956 102448 282826 102504
rect 282882 102448 282887 102504
rect 279956 102446 282887 102448
rect 282821 102443 282887 102446
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 231577 102370 231643 102373
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 228804 102368 231643 102370
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 228804 102312 231582 102368
rect 231638 102312 231643 102368
rect 228804 102310 231643 102312
rect 65977 102307 66043 102310
rect 231577 102307 231643 102310
rect 213913 102234 213979 102237
rect 264973 102234 265039 102237
rect 287010 102234 287070 102582
rect 295374 102234 295380 102236
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 264973 102232 268180 102234
rect 264973 102176 264978 102232
rect 265034 102176 268180 102232
rect 264973 102174 268180 102176
rect 287010 102174 295380 102234
rect 213913 102171 213979 102174
rect 264973 102171 265039 102174
rect 295374 102172 295380 102174
rect 295444 102172 295450 102236
rect 231117 101826 231183 101829
rect 228804 101824 231183 101826
rect 228804 101768 231122 101824
rect 231178 101768 231183 101824
rect 228804 101766 231183 101768
rect 231117 101763 231183 101766
rect 265341 101826 265407 101829
rect 265341 101824 268180 101826
rect 265341 101768 265346 101824
rect 265402 101768 268180 101824
rect 265341 101766 268180 101768
rect 265341 101763 265407 101766
rect 281809 101690 281875 101693
rect 279956 101688 281875 101690
rect 279956 101632 281814 101688
rect 281870 101632 281875 101688
rect 279956 101630 281875 101632
rect 281809 101627 281875 101630
rect 214741 101554 214807 101557
rect 214741 101552 217212 101554
rect 214741 101496 214746 101552
rect 214802 101496 217212 101552
rect 214741 101494 217212 101496
rect 214741 101491 214807 101494
rect 231761 101418 231827 101421
rect 228804 101416 231827 101418
rect 228804 101360 231766 101416
rect 231822 101360 231827 101416
rect 228804 101358 231827 101360
rect 231761 101355 231827 101358
rect 264973 101282 265039 101285
rect 264973 101280 268180 101282
rect 264973 101224 264978 101280
rect 265034 101224 268180 101280
rect 264973 101222 268180 101224
rect 264973 101219 265039 101222
rect 213913 101010 213979 101013
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 213913 100947 213979 100950
rect 231301 100874 231367 100877
rect 228804 100872 231367 100874
rect 228804 100816 231306 100872
rect 231362 100816 231367 100872
rect 228804 100814 231367 100816
rect 231301 100811 231367 100814
rect 265065 100874 265131 100877
rect 281533 100874 281599 100877
rect 265065 100872 268180 100874
rect 265065 100816 265070 100872
rect 265126 100816 268180 100872
rect 265065 100814 268180 100816
rect 279956 100872 281599 100874
rect 279956 100816 281538 100872
rect 281594 100816 281599 100872
rect 279956 100814 281599 100816
rect 265065 100811 265131 100814
rect 281533 100811 281599 100814
rect 67633 100738 67699 100741
rect 68142 100738 68816 100744
rect 67633 100736 68816 100738
rect 67633 100680 67638 100736
rect 67694 100684 68816 100736
rect 67694 100680 68202 100684
rect 67633 100678 68202 100680
rect 67633 100675 67699 100678
rect 230749 100466 230815 100469
rect 228804 100464 230815 100466
rect 228804 100408 230754 100464
rect 230810 100408 230815 100464
rect 228804 100406 230815 100408
rect 230749 100403 230815 100406
rect 214005 100330 214071 100333
rect 214005 100328 217212 100330
rect 214005 100272 214010 100328
rect 214066 100272 217212 100328
rect 214005 100270 217212 100272
rect 214005 100267 214071 100270
rect 267958 100132 267964 100196
rect 268028 100194 268034 100196
rect 268150 100194 268210 100436
rect 281717 100194 281783 100197
rect 268028 100134 268210 100194
rect 279956 100192 281783 100194
rect 279956 100136 281722 100192
rect 281778 100136 281783 100192
rect 279956 100134 281783 100136
rect 268028 100132 268034 100134
rect 281717 100131 281783 100134
rect 265065 100058 265131 100061
rect 265065 100056 268180 100058
rect 265065 100000 265070 100056
rect 265126 100000 268180 100056
rect 265065 99998 268180 100000
rect 265065 99995 265131 99998
rect 231117 99922 231183 99925
rect 228804 99920 231183 99922
rect 228804 99864 231122 99920
rect 231178 99864 231183 99920
rect 228804 99862 231183 99864
rect 231117 99859 231183 99862
rect 213913 99650 213979 99653
rect 264973 99650 265039 99653
rect 213913 99648 217212 99650
rect 213913 99592 213918 99648
rect 213974 99592 217212 99648
rect 213913 99590 217212 99592
rect 264973 99648 268180 99650
rect 264973 99592 264978 99648
rect 265034 99592 268180 99648
rect 264973 99590 268180 99592
rect 213913 99587 213979 99590
rect 264973 99587 265039 99590
rect 231577 99514 231643 99517
rect 228804 99512 231643 99514
rect 228804 99456 231582 99512
rect 231638 99456 231643 99512
rect 228804 99454 231643 99456
rect 231577 99451 231643 99454
rect 583293 99514 583359 99517
rect 583520 99514 584960 99604
rect 583293 99512 584960 99514
rect 583293 99456 583298 99512
rect 583354 99456 584960 99512
rect 583293 99454 584960 99456
rect 583293 99451 583359 99454
rect 282821 99378 282887 99381
rect 279956 99376 282887 99378
rect 279956 99320 282826 99376
rect 282882 99320 282887 99376
rect 583520 99364 584960 99454
rect 279956 99318 282887 99320
rect 282821 99315 282887 99318
rect 265065 99242 265131 99245
rect 265065 99240 268180 99242
rect 265065 99184 265070 99240
rect 265126 99184 268180 99240
rect 265065 99182 268180 99184
rect 265065 99179 265131 99182
rect 214005 98970 214071 98973
rect 231209 98970 231275 98973
rect 214005 98968 217212 98970
rect 214005 98912 214010 98968
rect 214066 98912 217212 98968
rect 214005 98910 217212 98912
rect 228804 98968 231275 98970
rect 228804 98912 231214 98968
rect 231270 98912 231275 98968
rect 228804 98910 231275 98912
rect 214005 98907 214071 98910
rect 231209 98907 231275 98910
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 264973 98635 265039 98638
rect 230657 98562 230723 98565
rect 228804 98560 230723 98562
rect 228804 98504 230662 98560
rect 230718 98504 230723 98560
rect 228804 98502 230723 98504
rect 230657 98499 230723 98502
rect 213913 98290 213979 98293
rect 213913 98288 217212 98290
rect 213913 98232 213918 98288
rect 213974 98232 217212 98288
rect 213913 98230 217212 98232
rect 213913 98227 213979 98230
rect 229134 98228 229140 98292
rect 229204 98290 229210 98292
rect 229204 98230 268180 98290
rect 229204 98228 229210 98230
rect 279374 98157 279434 98532
rect 279325 98152 279434 98157
rect 279325 98096 279330 98152
rect 279386 98096 279434 98152
rect 279325 98094 279434 98096
rect 279325 98091 279391 98094
rect 231117 98018 231183 98021
rect 228804 98016 231183 98018
rect 228804 97960 231122 98016
rect 231178 97960 231183 98016
rect 228804 97958 231183 97960
rect 231117 97955 231183 97958
rect 264973 97882 265039 97885
rect 282821 97882 282887 97885
rect 264973 97880 268180 97882
rect 264973 97824 264978 97880
rect 265034 97824 268180 97880
rect 264973 97822 268180 97824
rect 279956 97880 282887 97882
rect 279956 97824 282826 97880
rect 282882 97824 282887 97880
rect 279956 97822 282887 97824
rect 264973 97819 265039 97822
rect 282821 97819 282887 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 213913 97610 213979 97613
rect 231669 97610 231735 97613
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 228804 97608 231735 97610
rect 228804 97552 231674 97608
rect 231730 97552 231735 97608
rect 228804 97550 231735 97552
rect 213913 97547 213979 97550
rect 231669 97547 231735 97550
rect 265157 97474 265223 97477
rect 265157 97472 268180 97474
rect 265157 97416 265162 97472
rect 265218 97416 268180 97472
rect 265157 97414 268180 97416
rect 265157 97411 265223 97414
rect 229185 97204 229251 97205
rect 229134 97202 229140 97204
rect 229094 97142 229140 97202
rect 229204 97200 229251 97204
rect 229246 97144 229251 97200
rect 229134 97140 229140 97142
rect 229204 97140 229251 97144
rect 229185 97139 229251 97140
rect 229093 97066 229159 97069
rect 228804 97064 229159 97066
rect 228804 97008 229098 97064
rect 229154 97008 229159 97064
rect 228804 97006 229159 97008
rect 229093 97003 229159 97006
rect 265065 97066 265131 97069
rect 282177 97066 282243 97069
rect 265065 97064 268180 97066
rect 265065 97008 265070 97064
rect 265126 97008 268180 97064
rect 265065 97006 268180 97008
rect 279956 97064 282243 97066
rect 279956 97008 282182 97064
rect 282238 97008 282243 97064
rect 279956 97006 282243 97008
rect 265065 97003 265131 97006
rect 282177 97003 282243 97006
rect 214005 96930 214071 96933
rect 214005 96928 217212 96930
rect 214005 96872 214010 96928
rect 214066 96872 217212 96928
rect 214005 96870 217212 96872
rect 214005 96867 214071 96870
rect 229185 96658 229251 96661
rect 228804 96656 229251 96658
rect 228804 96600 229190 96656
rect 229246 96600 229251 96656
rect 228804 96598 229251 96600
rect 229185 96595 229251 96598
rect 264973 96658 265039 96661
rect 264973 96656 268180 96658
rect 264973 96600 264978 96656
rect 265034 96600 268180 96656
rect 264973 96598 268180 96600
rect 264973 96595 265039 96598
rect 214097 96386 214163 96389
rect 214097 96384 217212 96386
rect 214097 96328 214102 96384
rect 214158 96328 217212 96384
rect 214097 96326 217212 96328
rect 214097 96323 214163 96326
rect 231117 96250 231183 96253
rect 228804 96248 231183 96250
rect 228804 96192 231122 96248
rect 231178 96192 231183 96248
rect 228804 96190 231183 96192
rect 231117 96187 231183 96190
rect 264973 96250 265039 96253
rect 264973 96248 268180 96250
rect 264973 96192 264978 96248
rect 265034 96192 268180 96248
rect 264973 96190 268180 96192
rect 264973 96187 265039 96190
rect 279233 96114 279299 96117
rect 279374 96114 279434 96356
rect 279233 96112 279434 96114
rect 279233 96056 279238 96112
rect 279294 96056 279434 96112
rect 279233 96054 279434 96056
rect 279233 96051 279299 96054
rect 226374 95916 226380 95980
rect 226444 95978 226450 95980
rect 228950 95978 228956 95980
rect 226444 95918 228956 95978
rect 226444 95916 226450 95918
rect 228950 95916 228956 95918
rect 229020 95916 229026 95980
rect 197118 95100 197124 95164
rect 197188 95162 197194 95164
rect 281533 95162 281599 95165
rect 197188 95160 281599 95162
rect 197188 95104 281538 95160
rect 281594 95104 281599 95160
rect 197188 95102 281599 95104
rect 197188 95100 197194 95102
rect 281533 95099 281599 95102
rect 59261 95026 59327 95029
rect 215017 95026 215083 95029
rect 59261 95024 215083 95026
rect 59261 94968 59266 95024
rect 59322 94968 215022 95024
rect 215078 94968 215083 95024
rect 59261 94966 215083 94968
rect 59261 94963 59327 94966
rect 215017 94963 215083 94966
rect 151629 94892 151695 94893
rect 151624 94890 151630 94892
rect 151538 94830 151630 94890
rect 151624 94828 151630 94830
rect 151694 94828 151700 94892
rect 151629 94827 151695 94828
rect 109033 94756 109099 94757
rect 110689 94756 110755 94757
rect 115841 94756 115907 94757
rect 119429 94756 119495 94757
rect 109033 94754 109062 94756
rect 108970 94752 109062 94754
rect 108970 94696 109038 94752
rect 108970 94694 109062 94696
rect 109033 94692 109062 94694
rect 109126 94692 109132 94756
rect 110688 94754 110694 94756
rect 110602 94694 110694 94754
rect 110688 94692 110694 94694
rect 110758 94692 110764 94756
rect 115841 94754 115862 94756
rect 115770 94752 115862 94754
rect 115770 94696 115846 94752
rect 115770 94694 115862 94696
rect 115841 94692 115862 94694
rect 115926 94692 115932 94756
rect 119392 94692 119398 94756
rect 119462 94754 119495 94756
rect 119462 94752 119554 94754
rect 119490 94696 119554 94752
rect 119462 94694 119554 94696
rect 119462 94692 119495 94694
rect 109033 94691 109099 94692
rect 110689 94691 110755 94692
rect 115841 94691 115907 94692
rect 119429 94691 119495 94692
rect 267590 94420 267596 94484
rect 267660 94482 267666 94484
rect 270585 94482 270651 94485
rect 267660 94480 270651 94482
rect 267660 94424 270590 94480
rect 270646 94424 270651 94480
rect 267660 94422 270651 94424
rect 267660 94420 267666 94422
rect 270585 94419 270651 94422
rect 104566 93876 104572 93940
rect 104636 93938 104642 93940
rect 167729 93938 167795 93941
rect 104636 93936 167795 93938
rect 104636 93880 167734 93936
rect 167790 93880 167795 93936
rect 104636 93878 167795 93880
rect 104636 93876 104642 93878
rect 167729 93875 167795 93878
rect 224217 93938 224283 93941
rect 229686 93938 229692 93940
rect 224217 93936 229692 93938
rect 224217 93880 224222 93936
rect 224278 93880 229692 93936
rect 224217 93878 229692 93880
rect 224217 93875 224283 93878
rect 229686 93876 229692 93878
rect 229756 93876 229762 93940
rect 66069 93802 66135 93805
rect 180149 93802 180215 93805
rect 66069 93800 180215 93802
rect 66069 93744 66074 93800
rect 66130 93744 180154 93800
rect 180210 93744 180215 93800
rect 66069 93742 180215 93744
rect 66069 93739 66135 93742
rect 180149 93739 180215 93742
rect 116710 93604 116716 93668
rect 116780 93666 116786 93668
rect 169017 93666 169083 93669
rect 116780 93664 169083 93666
rect 116780 93608 169022 93664
rect 169078 93608 169083 93664
rect 116780 93606 169083 93608
rect 116780 93604 116786 93606
rect 169017 93603 169083 93606
rect 100569 93532 100635 93533
rect 105537 93532 105603 93533
rect 118233 93532 118299 93533
rect 125409 93532 125475 93533
rect 151537 93532 151603 93533
rect 152089 93532 152155 93533
rect 100518 93530 100524 93532
rect 100478 93470 100524 93530
rect 100588 93528 100635 93532
rect 105486 93530 105492 93532
rect 100630 93472 100635 93528
rect 100518 93468 100524 93470
rect 100588 93468 100635 93472
rect 105446 93470 105492 93530
rect 105556 93528 105603 93532
rect 118182 93530 118188 93532
rect 105598 93472 105603 93528
rect 105486 93468 105492 93470
rect 105556 93468 105603 93472
rect 118142 93470 118188 93530
rect 118252 93528 118299 93532
rect 125358 93530 125364 93532
rect 118294 93472 118299 93528
rect 118182 93468 118188 93470
rect 118252 93468 118299 93472
rect 125318 93470 125364 93530
rect 125428 93528 125475 93532
rect 151486 93530 151492 93532
rect 125470 93472 125475 93528
rect 125358 93468 125364 93470
rect 125428 93468 125475 93472
rect 151446 93470 151492 93530
rect 151556 93528 151603 93532
rect 152038 93530 152044 93532
rect 151598 93472 151603 93528
rect 151486 93468 151492 93470
rect 151556 93468 151603 93472
rect 151998 93470 152044 93530
rect 152108 93528 152155 93532
rect 152150 93472 152155 93528
rect 152038 93468 152044 93470
rect 152108 93468 152155 93472
rect 100569 93467 100635 93468
rect 105537 93467 105603 93468
rect 118233 93467 118299 93468
rect 125409 93467 125475 93468
rect 151537 93467 151603 93468
rect 152089 93467 152155 93468
rect 110137 93260 110203 93261
rect 113817 93260 113883 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 113766 93258 113772 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 113726 93198 113772 93258
rect 113836 93256 113883 93260
rect 113878 93200 113883 93256
rect 113766 93196 113772 93198
rect 113836 93196 113883 93200
rect 110137 93195 110203 93196
rect 113817 93195 113883 93196
rect 74809 92444 74875 92445
rect 85849 92444 85915 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 85798 92442 85804 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 85758 92382 85804 92442
rect 85868 92440 85915 92444
rect 85910 92384 85915 92440
rect 85798 92380 85804 92382
rect 85868 92380 85915 92384
rect 91318 92380 91324 92444
rect 91388 92442 91394 92444
rect 91461 92442 91527 92445
rect 91388 92440 91527 92442
rect 91388 92384 91466 92440
rect 91522 92384 91527 92440
rect 91388 92382 91527 92384
rect 91388 92380 91394 92382
rect 74809 92379 74875 92380
rect 85849 92379 85915 92380
rect 91461 92379 91527 92382
rect 98494 92380 98500 92444
rect 98564 92442 98570 92444
rect 99005 92442 99071 92445
rect 98564 92440 99071 92442
rect 98564 92384 99010 92440
rect 99066 92384 99071 92440
rect 98564 92382 99071 92384
rect 98564 92380 98570 92382
rect 99005 92379 99071 92382
rect 104198 92380 104204 92444
rect 104268 92442 104274 92444
rect 104433 92442 104499 92445
rect 105721 92444 105787 92445
rect 105670 92442 105676 92444
rect 104268 92440 104499 92442
rect 104268 92384 104438 92440
rect 104494 92384 104499 92440
rect 104268 92382 104499 92384
rect 105630 92382 105676 92442
rect 105740 92440 105787 92444
rect 105782 92384 105787 92440
rect 104268 92380 104274 92382
rect 104433 92379 104499 92382
rect 105670 92380 105676 92382
rect 105740 92380 105787 92384
rect 106406 92380 106412 92444
rect 106476 92442 106482 92444
rect 106733 92442 106799 92445
rect 109585 92444 109651 92445
rect 113265 92444 113331 92445
rect 109534 92442 109540 92444
rect 106476 92440 106799 92442
rect 106476 92384 106738 92440
rect 106794 92384 106799 92440
rect 106476 92382 106799 92384
rect 109494 92382 109540 92442
rect 109604 92440 109651 92444
rect 113214 92442 113220 92444
rect 109646 92384 109651 92440
rect 106476 92380 106482 92382
rect 105721 92379 105787 92380
rect 106733 92379 106799 92382
rect 109534 92380 109540 92382
rect 109604 92380 109651 92384
rect 113174 92382 113220 92442
rect 113284 92440 113331 92444
rect 113326 92384 113331 92440
rect 113214 92380 113220 92382
rect 113284 92380 113331 92384
rect 115422 92380 115428 92444
rect 115492 92442 115498 92444
rect 115749 92442 115815 92445
rect 115492 92440 115815 92442
rect 115492 92384 115754 92440
rect 115810 92384 115815 92440
rect 115492 92382 115815 92384
rect 115492 92380 115498 92382
rect 109585 92379 109651 92380
rect 113265 92379 113331 92380
rect 115749 92379 115815 92382
rect 120574 92380 120580 92444
rect 120644 92442 120650 92444
rect 121177 92442 121243 92445
rect 123017 92444 123083 92445
rect 125777 92444 125843 92445
rect 122966 92442 122972 92444
rect 120644 92440 121243 92442
rect 120644 92384 121182 92440
rect 121238 92384 121243 92440
rect 120644 92382 121243 92384
rect 122926 92382 122972 92442
rect 123036 92440 123083 92444
rect 125726 92442 125732 92444
rect 123078 92384 123083 92440
rect 120644 92380 120650 92382
rect 121177 92379 121243 92382
rect 122966 92380 122972 92382
rect 123036 92380 123083 92384
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 125838 92384 125843 92440
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 136030 92380 136036 92444
rect 136100 92442 136106 92444
rect 136173 92442 136239 92445
rect 136100 92440 136239 92442
rect 136100 92384 136178 92440
rect 136234 92384 136239 92440
rect 136100 92382 136239 92384
rect 136100 92380 136106 92382
rect 123017 92379 123083 92380
rect 125777 92379 125843 92380
rect 136173 92379 136239 92382
rect 117998 92244 118004 92308
rect 118068 92306 118074 92308
rect 166206 92306 166212 92308
rect 118068 92246 166212 92306
rect 118068 92244 118074 92246
rect 166206 92244 166212 92246
rect 166276 92244 166282 92308
rect 103830 92108 103836 92172
rect 103900 92170 103906 92172
rect 174629 92170 174695 92173
rect 103900 92168 174695 92170
rect 103900 92112 174634 92168
rect 174690 92112 174695 92168
rect 103900 92110 174695 92112
rect 103900 92108 103906 92110
rect 174629 92107 174695 92110
rect 90214 91836 90220 91900
rect 90284 91898 90290 91900
rect 91001 91898 91067 91901
rect 90284 91896 91067 91898
rect 90284 91840 91006 91896
rect 91062 91840 91067 91896
rect 90284 91838 91067 91840
rect 90284 91836 90290 91838
rect 91001 91835 91067 91838
rect 84326 91700 84332 91764
rect 84396 91762 84402 91764
rect 85021 91762 85087 91765
rect 84396 91760 85087 91762
rect 84396 91704 85026 91760
rect 85082 91704 85087 91760
rect 84396 91702 85087 91704
rect 84396 91700 84402 91702
rect 85021 91699 85087 91702
rect 97206 91700 97212 91764
rect 97276 91762 97282 91764
rect 97349 91762 97415 91765
rect 101857 91764 101923 91765
rect 117129 91764 117195 91765
rect 101806 91762 101812 91764
rect 97276 91760 97415 91762
rect 97276 91704 97354 91760
rect 97410 91704 97415 91760
rect 97276 91702 97415 91704
rect 101766 91702 101812 91762
rect 101876 91760 101923 91764
rect 117078 91762 117084 91764
rect 101918 91704 101923 91760
rect 97276 91700 97282 91702
rect 97349 91699 97415 91702
rect 101806 91700 101812 91702
rect 101876 91700 101923 91704
rect 117038 91702 117084 91762
rect 117148 91760 117195 91764
rect 117190 91704 117195 91760
rect 117078 91700 117084 91702
rect 117148 91700 117195 91704
rect 101857 91699 101923 91700
rect 117129 91699 117195 91700
rect 222929 91762 222995 91765
rect 230974 91762 230980 91764
rect 222929 91760 230980 91762
rect 222929 91704 222934 91760
rect 222990 91704 230980 91760
rect 222929 91702 230980 91704
rect 222929 91699 222995 91702
rect 230974 91700 230980 91702
rect 231044 91700 231050 91764
rect 86769 91628 86835 91629
rect 86718 91626 86724 91628
rect 86678 91566 86724 91626
rect 86788 91624 86835 91628
rect 86830 91568 86835 91624
rect 86718 91564 86724 91566
rect 86788 91564 86835 91568
rect 126462 91564 126468 91628
rect 126532 91626 126538 91628
rect 126605 91626 126671 91629
rect 126532 91624 126671 91626
rect 126532 91568 126610 91624
rect 126666 91568 126671 91624
rect 126532 91566 126671 91568
rect 126532 91564 126538 91566
rect 86769 91563 86835 91564
rect 126605 91563 126671 91566
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 101949 91354 102015 91357
rect 100956 91352 102015 91354
rect 100956 91296 101954 91352
rect 102010 91296 102015 91352
rect 100956 91294 102015 91296
rect 100956 91292 100962 91294
rect 101949 91291 102015 91294
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89161 91218 89227 91221
rect 88996 91216 89227 91218
rect 88996 91160 89166 91216
rect 89222 91160 89227 91216
rect 88996 91158 89227 91160
rect 88996 91156 89002 91158
rect 88057 91155 88123 91156
rect 89161 91155 89227 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93117 91218 93183 91221
rect 92676 91216 93183 91218
rect 92676 91160 93122 91216
rect 93178 91160 93183 91216
rect 92676 91158 93183 91160
rect 92676 91156 92682 91158
rect 93117 91155 93183 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 94405 91218 94471 91221
rect 93964 91216 94471 91218
rect 93964 91160 94410 91216
rect 94466 91160 94471 91216
rect 93964 91158 94471 91160
rect 93964 91156 93970 91158
rect 94405 91155 94471 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 96337 91220 96403 91221
rect 96286 91218 96292 91220
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 96246 91158 96292 91218
rect 96356 91216 96403 91220
rect 96398 91160 96403 91216
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91158
rect 96356 91156 96403 91160
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97809 91218 97875 91221
rect 96724 91216 97875 91218
rect 96724 91160 97814 91216
rect 97870 91160 97875 91216
rect 96724 91158 97875 91160
rect 96724 91156 96730 91158
rect 96337 91155 96403 91156
rect 97809 91155 97875 91158
rect 98126 91156 98132 91220
rect 98196 91218 98202 91220
rect 98729 91218 98795 91221
rect 99097 91220 99163 91221
rect 99046 91218 99052 91220
rect 98196 91216 98795 91218
rect 98196 91160 98734 91216
rect 98790 91160 98795 91216
rect 98196 91158 98795 91160
rect 99006 91158 99052 91218
rect 99116 91216 99163 91220
rect 99158 91160 99163 91216
rect 98196 91156 98202 91158
rect 98729 91155 98795 91158
rect 99046 91156 99052 91158
rect 99116 91156 99163 91160
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100201 91218 100267 91221
rect 102041 91220 102107 91221
rect 101990 91218 101996 91220
rect 100036 91216 100267 91218
rect 100036 91160 100206 91216
rect 100262 91160 100267 91216
rect 100036 91158 100267 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 102102 91160 102107 91216
rect 100036 91156 100042 91158
rect 99097 91155 99163 91156
rect 100201 91155 100267 91158
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 102869 91218 102935 91221
rect 102796 91216 102935 91218
rect 102796 91160 102874 91216
rect 102930 91160 102935 91216
rect 102796 91158 102935 91160
rect 102796 91156 102802 91158
rect 102041 91155 102107 91156
rect 102869 91155 102935 91158
rect 106774 91156 106780 91220
rect 106844 91218 106850 91220
rect 107561 91218 107627 91221
rect 106844 91216 107627 91218
rect 106844 91160 107566 91216
rect 107622 91160 107627 91216
rect 106844 91158 107627 91160
rect 106844 91156 106850 91158
rect 107561 91155 107627 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 107929 91218 107995 91221
rect 107764 91216 107995 91218
rect 107764 91160 107934 91216
rect 107990 91160 107995 91216
rect 107764 91158 107995 91160
rect 107764 91156 107770 91158
rect 107929 91155 107995 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111333 91218 111399 91221
rect 111260 91216 111399 91218
rect 111260 91160 111338 91216
rect 111394 91160 111399 91216
rect 111260 91158 111399 91160
rect 111260 91156 111266 91158
rect 111333 91155 111399 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 112069 91218 112135 91221
rect 111996 91216 112135 91218
rect 111996 91160 112074 91216
rect 112130 91160 112135 91216
rect 111996 91158 112135 91160
rect 111996 91156 112002 91158
rect 112069 91155 112135 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112713 91218 112779 91221
rect 112364 91216 112779 91218
rect 112364 91160 112718 91216
rect 112774 91160 112779 91216
rect 112364 91158 112779 91160
rect 112364 91156 112370 91158
rect 112713 91155 112779 91158
rect 114318 91156 114324 91220
rect 114388 91218 114394 91220
rect 114461 91218 114527 91221
rect 114388 91216 114527 91218
rect 114388 91160 114466 91216
rect 114522 91160 114527 91216
rect 114388 91158 114527 91160
rect 114388 91156 114394 91158
rect 114461 91155 114527 91158
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115013 91218 115079 91221
rect 119705 91220 119771 91221
rect 119654 91218 119660 91220
rect 114940 91216 115079 91218
rect 114940 91160 115018 91216
rect 115074 91160 115079 91216
rect 114940 91158 115079 91160
rect 119614 91158 119660 91218
rect 119724 91216 119771 91220
rect 119766 91160 119771 91216
rect 114940 91156 114946 91158
rect 115013 91155 115079 91158
rect 119654 91156 119660 91158
rect 119724 91156 119771 91160
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121269 91218 121335 91221
rect 120276 91216 121335 91218
rect 120276 91160 121274 91216
rect 121330 91160 121335 91216
rect 120276 91158 121335 91160
rect 120276 91156 120282 91158
rect 119705 91155 119771 91156
rect 121269 91155 121335 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 121913 91218 121979 91221
rect 121748 91216 121979 91218
rect 121748 91160 121918 91216
rect 121974 91160 121979 91216
rect 121748 91158 121979 91160
rect 121748 91156 121754 91158
rect 121913 91155 121979 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 123293 91218 123359 91221
rect 124121 91220 124187 91221
rect 124070 91218 124076 91220
rect 123220 91216 123359 91218
rect 123220 91160 123298 91216
rect 123354 91160 123359 91216
rect 123220 91158 123359 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 124182 91160 124187 91216
rect 123220 91156 123226 91158
rect 123293 91155 123359 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 124121 91155 124187 91156
rect 126881 91155 126947 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 127636 91156 127642 91158
rect 128261 91155 128327 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 132401 91220 132467 91221
rect 132350 91218 132356 91220
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133781 91218 133847 91221
rect 133156 91216 133847 91218
rect 133156 91160 133786 91216
rect 133842 91160 133847 91216
rect 133156 91158 133847 91160
rect 133156 91156 133162 91158
rect 132401 91155 132467 91156
rect 133781 91155 133847 91158
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 135161 91218 135227 91221
rect 151721 91220 151787 91221
rect 151670 91218 151676 91220
rect 134444 91216 135227 91218
rect 134444 91160 135166 91216
rect 135222 91160 135227 91216
rect 134444 91158 135227 91160
rect 151630 91158 151676 91218
rect 151740 91216 151787 91220
rect 151782 91160 151787 91216
rect 134444 91156 134450 91158
rect 135161 91155 135227 91158
rect 151670 91156 151676 91158
rect 151740 91156 151787 91160
rect 151721 91155 151787 91156
rect 67449 91082 67515 91085
rect 214833 91082 214899 91085
rect 67449 91080 214899 91082
rect 67449 91024 67454 91080
rect 67510 91024 214838 91080
rect 214894 91024 214899 91080
rect 67449 91022 214899 91024
rect 67449 91019 67515 91022
rect 214833 91019 214899 91022
rect 124438 90884 124444 90948
rect 124508 90946 124514 90948
rect 177389 90946 177455 90949
rect 124508 90944 177455 90946
rect 124508 90888 177394 90944
rect 177450 90888 177455 90944
rect 124508 90886 177455 90888
rect 124508 90884 124514 90886
rect 177389 90883 177455 90886
rect 91001 89722 91067 89725
rect 184381 89722 184447 89725
rect 91001 89720 184447 89722
rect 91001 89664 91006 89720
rect 91062 89664 184386 89720
rect 184442 89664 184447 89720
rect 91001 89662 184447 89664
rect 91001 89659 91067 89662
rect 184381 89659 184447 89662
rect 85021 89586 85087 89589
rect 176009 89586 176075 89589
rect 85021 89584 176075 89586
rect 85021 89528 85026 89584
rect 85082 89528 176014 89584
rect 176070 89528 176075 89584
rect 85021 89526 176075 89528
rect 85021 89523 85087 89526
rect 176009 89523 176075 89526
rect 214557 89042 214623 89045
rect 244774 89042 244780 89044
rect 214557 89040 244780 89042
rect 214557 88984 214562 89040
rect 214618 88984 244780 89040
rect 214557 88982 244780 88984
rect 214557 88979 214623 88982
rect 244774 88980 244780 88982
rect 244844 88980 244850 89044
rect 123293 88226 123359 88229
rect 189717 88226 189783 88229
rect 123293 88224 189783 88226
rect 123293 88168 123298 88224
rect 123354 88168 189722 88224
rect 189778 88168 189783 88224
rect 123293 88166 189783 88168
rect 123293 88163 123359 88166
rect 189717 88163 189783 88166
rect 62021 86866 62087 86869
rect 214741 86866 214807 86869
rect 62021 86864 214807 86866
rect 62021 86808 62026 86864
rect 62082 86808 214746 86864
rect 214802 86808 214807 86864
rect 62021 86806 214807 86808
rect 62021 86803 62087 86806
rect 214741 86803 214807 86806
rect 582833 86186 582899 86189
rect 583520 86186 584960 86276
rect 582833 86184 584960 86186
rect 582833 86128 582838 86184
rect 582894 86128 584960 86184
rect 582833 86126 584960 86128
rect 582833 86123 582899 86126
rect 583520 86036 584960 86126
rect 119981 84826 120047 84829
rect 257521 84826 257587 84829
rect 119981 84824 257587 84826
rect -960 84690 480 84780
rect 119981 84768 119986 84824
rect 120042 84768 257526 84824
rect 257582 84768 257587 84824
rect 119981 84766 257587 84768
rect 119981 84763 120047 84766
rect 257521 84763 257587 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 19241 66874 19307 66877
rect 250294 66874 250300 66876
rect 19241 66872 250300 66874
rect 19241 66816 19246 66872
rect 19302 66816 250300 66872
rect 19241 66814 250300 66816
rect 19241 66811 19307 66814
rect 250294 66812 250300 66814
rect 250364 66812 250370 66876
rect 23381 65514 23447 65517
rect 253054 65514 253060 65516
rect 23381 65512 253060 65514
rect 23381 65456 23386 65512
rect 23442 65456 253060 65512
rect 23381 65454 253060 65456
rect 23381 65451 23447 65454
rect 253054 65452 253060 65454
rect 253124 65452 253130 65516
rect 57881 61434 57947 61437
rect 232446 61434 232452 61436
rect 57881 61432 232452 61434
rect 57881 61376 57886 61432
rect 57942 61376 232452 61432
rect 57881 61374 232452 61376
rect 57881 61371 57947 61374
rect 232446 61372 232452 61374
rect 232516 61372 232522 61436
rect 22001 59938 22067 59941
rect 267958 59938 267964 59940
rect 22001 59936 267964 59938
rect 22001 59880 22006 59936
rect 22062 59880 267964 59936
rect 22001 59878 267964 59880
rect 22001 59875 22067 59878
rect 267958 59876 267964 59878
rect 268028 59876 268034 59940
rect 582741 59666 582807 59669
rect 583520 59666 584960 59756
rect 582741 59664 584960 59666
rect 582741 59608 582746 59664
rect 582802 59608 584960 59664
rect 582741 59606 584960 59608
rect 582741 59603 582807 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 33041 57218 33107 57221
rect 258574 57218 258580 57220
rect 33041 57216 258580 57218
rect 33041 57160 33046 57216
rect 33102 57160 258580 57216
rect 33041 57158 258580 57160
rect 33041 57155 33107 57158
rect 258574 57156 258580 57158
rect 258644 57156 258650 57220
rect 16481 50282 16547 50285
rect 226374 50282 226380 50284
rect 16481 50280 226380 50282
rect 16481 50224 16486 50280
rect 16542 50224 226380 50280
rect 16481 50222 226380 50224
rect 16481 50219 16547 50222
rect 226374 50220 226380 50222
rect 226444 50220 226450 50284
rect 582649 46338 582715 46341
rect 583520 46338 584960 46428
rect 582649 46336 584960 46338
rect 582649 46280 582654 46336
rect 582710 46280 584960 46336
rect 582649 46278 584960 46280
rect 582649 46275 582715 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 67541 43482 67607 43485
rect 251766 43482 251772 43484
rect 67541 43480 251772 43482
rect 67541 43424 67546 43480
rect 67602 43424 251772 43480
rect 67541 43422 251772 43424
rect 67541 43419 67607 43422
rect 251766 43420 251772 43422
rect 251836 43420 251842 43484
rect 582557 33146 582623 33149
rect 583520 33146 584960 33236
rect 582557 33144 584960 33146
rect 582557 33088 582562 33144
rect 582618 33088 584960 33144
rect 582557 33086 584960 33088
rect 582557 33083 582623 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 31661 30970 31727 30973
rect 262806 30970 262812 30972
rect 31661 30968 262812 30970
rect 31661 30912 31666 30968
rect 31722 30912 262812 30968
rect 31661 30910 262812 30912
rect 31661 30907 31727 30910
rect 262806 30908 262812 30910
rect 262876 30908 262882 30972
rect 28901 24170 28967 24173
rect 267774 24170 267780 24172
rect 28901 24168 267780 24170
rect 28901 24112 28906 24168
rect 28962 24112 267780 24168
rect 28901 24110 267780 24112
rect 28901 24107 28967 24110
rect 267774 24108 267780 24110
rect 267844 24108 267850 24172
rect 20621 21314 20687 21317
rect 228214 21314 228220 21316
rect 20621 21312 228220 21314
rect 20621 21256 20626 21312
rect 20682 21256 228220 21312
rect 20621 21254 228220 21256
rect 20621 21251 20687 21254
rect 228214 21252 228220 21254
rect 228284 21252 228290 21316
rect 13 19954 79 19957
rect 13 19952 122 19954
rect 13 19896 18 19952
rect 74 19896 122 19952
rect 13 19891 122 19896
rect 62 19546 122 19891
rect 582373 19818 582439 19821
rect 583520 19818 584960 19908
rect 582373 19816 584960 19818
rect 582373 19760 582378 19816
rect 582434 19760 584960 19816
rect 582373 19758 584960 19760
rect 582373 19755 582439 19758
rect 583520 19668 584960 19758
rect 62 19500 674 19546
rect -960 19486 674 19500
rect -960 19410 480 19486
rect 614 19410 674 19486
rect -960 19350 674 19410
rect -960 19260 480 19350
rect 582465 6626 582531 6629
rect 583520 6626 584960 6716
rect 582465 6624 584960 6626
rect -960 6490 480 6580
rect 582465 6568 582470 6624
rect 582526 6568 584960 6624
rect 582465 6566 584960 6568
rect 582465 6563 582531 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 121085 3362 121151 3365
rect 246246 3362 246252 3364
rect 121085 3360 246252 3362
rect 121085 3304 121090 3360
rect 121146 3304 246252 3360
rect 121085 3302 246252 3304
rect 121085 3299 121151 3302
rect 246246 3300 246252 3302
rect 246316 3300 246322 3364
<< via3 >>
rect 213132 699756 213196 699820
rect 285628 295292 285692 295356
rect 248460 291212 248524 291276
rect 278820 288628 278884 288692
rect 288388 288492 288452 288556
rect 280292 287132 280356 287196
rect 228220 286044 228284 286108
rect 244412 286044 244476 286108
rect 220860 285636 220924 285700
rect 287100 284412 287164 284476
rect 233188 284276 233252 284340
rect 201356 284004 201420 284068
rect 218100 284004 218164 284068
rect 231716 284004 231780 284068
rect 244228 284004 244292 284068
rect 204852 283928 204916 283932
rect 204852 283872 204902 283928
rect 204902 283872 204916 283928
rect 204852 283868 204916 283872
rect 210740 283928 210804 283932
rect 210740 283872 210754 283928
rect 210754 283872 210804 283928
rect 210740 283868 210804 283872
rect 212396 283868 212460 283932
rect 217548 283928 217612 283932
rect 217548 283872 217598 283928
rect 217598 283872 217612 283928
rect 217548 283868 217612 283872
rect 223436 283868 223500 283932
rect 224172 283928 224236 283932
rect 224172 283872 224222 283928
rect 224222 283872 224236 283928
rect 224172 283868 224236 283872
rect 226196 283868 226260 283932
rect 226380 283868 226444 283932
rect 229692 283868 229756 283932
rect 231532 283868 231596 283932
rect 249748 283188 249812 283252
rect 281580 279652 281644 279716
rect 198780 259388 198844 259452
rect 197124 252180 197188 252244
rect 248644 248644 248708 248708
rect 243492 246196 243556 246260
rect 244228 244216 244292 244220
rect 244228 244160 244242 244216
rect 244242 244160 244292 244216
rect 244228 244156 244292 244160
rect 244228 244020 244292 244084
rect 245884 243476 245948 243540
rect 198780 241436 198844 241500
rect 245884 240212 245948 240276
rect 204852 240076 204916 240140
rect 218100 240076 218164 240140
rect 229692 240136 229756 240140
rect 229692 240080 229742 240136
rect 229742 240080 229756 240136
rect 229692 240076 229756 240080
rect 213132 238580 213196 238644
rect 243492 238580 243556 238644
rect 237420 237356 237484 237420
rect 231532 235996 231596 236060
rect 244228 234696 244292 234700
rect 244228 234640 244242 234696
rect 244242 234640 244292 234696
rect 244228 234636 244292 234640
rect 284340 225524 284404 225588
rect 212396 224164 212460 224228
rect 231900 208932 231964 208996
rect 295380 206212 295444 206276
rect 231716 196012 231780 196076
rect 236500 196012 236564 196076
rect 287284 192476 287348 192540
rect 281764 190980 281828 191044
rect 274588 189620 274652 189684
rect 229692 187036 229756 187100
rect 245700 186900 245764 186964
rect 232084 185676 232148 185740
rect 280292 185540 280356 185604
rect 234660 184180 234724 184244
rect 210740 182956 210804 183020
rect 230428 182820 230492 182884
rect 288572 182820 288636 182884
rect 237604 181460 237668 181524
rect 284524 181324 284588 181388
rect 217548 180100 217612 180164
rect 240364 179964 240428 180028
rect 226380 178740 226444 178804
rect 201356 178060 201420 178124
rect 97028 177924 97092 177988
rect 226196 177924 226260 177988
rect 101996 177576 102060 177580
rect 101996 177520 102046 177576
rect 102046 177520 102060 177576
rect 101996 177516 102060 177520
rect 130700 177516 130764 177580
rect 228220 177380 228284 177444
rect 285812 177380 285876 177444
rect 120764 177244 120828 177308
rect 123156 177244 123220 177308
rect 129412 177304 129476 177308
rect 129412 177248 129462 177304
rect 129462 177248 129476 177304
rect 129412 177244 129476 177248
rect 233372 177244 233436 177308
rect 291148 177244 291212 177308
rect 100708 177108 100772 177172
rect 104572 176836 104636 176900
rect 105676 176760 105740 176764
rect 105676 176704 105726 176760
rect 105726 176704 105740 176760
rect 105676 176700 105740 176704
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176760 109604 176764
rect 109540 176704 109590 176760
rect 109590 176704 109604 176760
rect 109540 176700 109604 176704
rect 110644 176760 110708 176764
rect 110644 176704 110694 176760
rect 110694 176704 110708 176760
rect 110644 176700 110708 176704
rect 112116 176700 112180 176764
rect 113220 176700 113284 176764
rect 116900 176760 116964 176764
rect 116900 176704 116950 176760
rect 116950 176704 116964 176760
rect 116900 176700 116964 176704
rect 119476 176760 119540 176764
rect 119476 176704 119526 176760
rect 119526 176704 119540 176760
rect 119476 176700 119540 176704
rect 125732 176700 125796 176764
rect 127020 176700 127084 176764
rect 132356 176760 132420 176764
rect 132356 176704 132406 176760
rect 132406 176704 132420 176760
rect 132356 176700 132420 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176760 158916 176764
rect 158852 176704 158902 176760
rect 158902 176704 158916 176760
rect 158852 176700 158916 176704
rect 229140 176700 229204 176764
rect 283788 176564 283852 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 241652 176428 241716 176492
rect 238524 176020 238588 176084
rect 220860 175944 220924 175948
rect 220860 175888 220910 175944
rect 220910 175888 220924 175944
rect 220860 175884 220924 175888
rect 223436 175884 223500 175948
rect 224172 175808 224236 175812
rect 224172 175752 224222 175808
rect 224222 175752 224236 175808
rect 224172 175748 224236 175752
rect 114324 175612 114388 175676
rect 124444 175672 124508 175676
rect 124444 175616 124494 175672
rect 124494 175616 124508 175672
rect 118372 175536 118436 175540
rect 118372 175480 118422 175536
rect 118422 175480 118436 175536
rect 118372 175476 118436 175480
rect 121868 175536 121932 175540
rect 121868 175480 121918 175536
rect 121918 175480 121932 175536
rect 121868 175476 121932 175480
rect 124444 175612 124508 175616
rect 133092 175672 133156 175676
rect 133092 175616 133142 175672
rect 133142 175616 133156 175672
rect 133092 175612 133156 175616
rect 274588 175748 274652 175812
rect 279188 175748 279252 175812
rect 98316 175340 98380 175404
rect 115726 174992 115790 174996
rect 115726 174936 115754 174992
rect 115754 174936 115790 174992
rect 115726 174932 115790 174936
rect 230612 174932 230676 174996
rect 281764 173980 281828 174044
rect 279372 172076 279436 172140
rect 279372 166772 279436 166836
rect 230612 163372 230676 163436
rect 283788 163100 283852 163164
rect 229692 161604 229756 161668
rect 238524 159564 238588 159628
rect 281580 157796 281644 157860
rect 230428 156164 230492 156228
rect 240364 153852 240428 153916
rect 244228 153716 244292 153780
rect 231900 150996 231964 151060
rect 245700 147732 245764 147796
rect 233188 147188 233252 147252
rect 291148 146372 291212 146436
rect 249748 145556 249812 145620
rect 233372 145284 233436 145348
rect 230428 144740 230492 144804
rect 234660 144740 234724 144804
rect 284340 144740 284404 144804
rect 248644 143380 248708 143444
rect 285628 143108 285692 143172
rect 248460 142020 248524 142084
rect 230428 141612 230492 141676
rect 230980 141340 231044 141404
rect 229692 139980 229756 140044
rect 236500 139708 236564 139772
rect 246252 139572 246316 139636
rect 232084 139164 232148 139228
rect 237604 138756 237668 138820
rect 284524 138484 284588 138548
rect 229140 137260 229204 137324
rect 231164 137260 231228 137324
rect 241652 136308 241716 136372
rect 288572 134132 288636 134196
rect 280108 133996 280172 134060
rect 244780 131956 244844 132020
rect 232452 131548 232516 131612
rect 280476 129372 280540 129436
rect 258580 128828 258644 128892
rect 267780 128420 267844 128484
rect 267596 127876 267660 127940
rect 230980 127332 231044 127396
rect 287100 121756 287164 121820
rect 251772 119036 251836 119100
rect 230980 116588 231044 116652
rect 231164 115092 231228 115156
rect 262812 115092 262876 115156
rect 237420 114412 237484 114476
rect 253060 113868 253124 113932
rect 250300 113460 250364 113524
rect 288388 106388 288452 106452
rect 287284 106252 287348 106316
rect 285812 104756 285876 104820
rect 166212 102716 166276 102780
rect 295380 102172 295444 102236
rect 267964 100132 268028 100196
rect 229140 98228 229204 98292
rect 229140 97200 229204 97204
rect 229140 97144 229190 97200
rect 229190 97144 229204 97200
rect 229140 97140 229204 97144
rect 226380 95916 226444 95980
rect 228956 95916 229020 95980
rect 197124 95100 197188 95164
rect 151630 94888 151694 94892
rect 151630 94832 151634 94888
rect 151634 94832 151690 94888
rect 151690 94832 151694 94888
rect 151630 94828 151694 94832
rect 109062 94752 109126 94756
rect 109062 94696 109094 94752
rect 109094 94696 109126 94752
rect 109062 94692 109126 94696
rect 110694 94752 110758 94756
rect 110694 94696 110750 94752
rect 110750 94696 110758 94752
rect 110694 94692 110758 94696
rect 115862 94752 115926 94756
rect 115862 94696 115902 94752
rect 115902 94696 115926 94752
rect 115862 94692 115926 94696
rect 119398 94752 119462 94756
rect 119398 94696 119434 94752
rect 119434 94696 119462 94752
rect 119398 94692 119462 94696
rect 267596 94420 267660 94484
rect 104572 93876 104636 93940
rect 229692 93876 229756 93940
rect 116716 93604 116780 93668
rect 100524 93528 100588 93532
rect 100524 93472 100574 93528
rect 100574 93472 100588 93528
rect 100524 93468 100588 93472
rect 105492 93528 105556 93532
rect 105492 93472 105542 93528
rect 105542 93472 105556 93528
rect 105492 93468 105556 93472
rect 118188 93528 118252 93532
rect 118188 93472 118238 93528
rect 118238 93472 118252 93528
rect 118188 93468 118252 93472
rect 125364 93528 125428 93532
rect 125364 93472 125414 93528
rect 125414 93472 125428 93528
rect 125364 93468 125428 93472
rect 151492 93528 151556 93532
rect 151492 93472 151542 93528
rect 151542 93472 151556 93528
rect 151492 93468 151556 93472
rect 152044 93528 152108 93532
rect 152044 93472 152094 93528
rect 152094 93472 152108 93528
rect 152044 93468 152108 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 113772 93256 113836 93260
rect 113772 93200 113822 93256
rect 113822 93200 113836 93256
rect 113772 93196 113836 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 85804 92440 85868 92444
rect 85804 92384 85854 92440
rect 85854 92384 85868 92440
rect 85804 92380 85868 92384
rect 91324 92380 91388 92444
rect 98500 92380 98564 92444
rect 104204 92380 104268 92444
rect 105676 92440 105740 92444
rect 105676 92384 105726 92440
rect 105726 92384 105740 92440
rect 105676 92380 105740 92384
rect 106412 92380 106476 92444
rect 109540 92440 109604 92444
rect 109540 92384 109590 92440
rect 109590 92384 109604 92440
rect 109540 92380 109604 92384
rect 113220 92440 113284 92444
rect 113220 92384 113270 92440
rect 113270 92384 113284 92440
rect 113220 92380 113284 92384
rect 115428 92380 115492 92444
rect 120580 92380 120644 92444
rect 122972 92440 123036 92444
rect 122972 92384 123022 92440
rect 123022 92384 123036 92440
rect 122972 92380 123036 92384
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 136036 92380 136100 92444
rect 118004 92244 118068 92308
rect 166212 92244 166276 92308
rect 103836 92108 103900 92172
rect 90220 91836 90284 91900
rect 84332 91700 84396 91764
rect 97212 91700 97276 91764
rect 101812 91760 101876 91764
rect 101812 91704 101862 91760
rect 101862 91704 101876 91760
rect 101812 91700 101876 91704
rect 117084 91760 117148 91764
rect 117084 91704 117134 91760
rect 117134 91704 117148 91760
rect 117084 91700 117148 91704
rect 230980 91700 231044 91764
rect 86724 91624 86788 91628
rect 86724 91568 86774 91624
rect 86774 91568 86788 91624
rect 86724 91564 86788 91568
rect 126468 91564 126532 91628
rect 100892 91292 100956 91356
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 88932 91156 88996 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 95004 91156 95068 91220
rect 96292 91216 96356 91220
rect 96292 91160 96342 91216
rect 96342 91160 96356 91216
rect 96292 91156 96356 91160
rect 96660 91156 96724 91220
rect 98132 91156 98196 91220
rect 99052 91216 99116 91220
rect 99052 91160 99102 91216
rect 99102 91160 99116 91216
rect 99052 91156 99116 91160
rect 99972 91156 100036 91220
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 106780 91156 106844 91220
rect 107700 91156 107764 91220
rect 108068 91156 108132 91220
rect 111196 91156 111260 91220
rect 111932 91156 111996 91220
rect 112300 91156 112364 91220
rect 114324 91156 114388 91220
rect 114876 91156 114940 91220
rect 119660 91216 119724 91220
rect 119660 91160 119710 91216
rect 119710 91160 119724 91216
rect 119660 91156 119724 91160
rect 120212 91156 120276 91220
rect 121684 91156 121748 91220
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 126652 91156 126716 91220
rect 127572 91156 127636 91220
rect 129412 91156 129476 91220
rect 130700 91156 130764 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 133092 91156 133156 91220
rect 134380 91156 134444 91220
rect 151676 91216 151740 91220
rect 151676 91160 151726 91216
rect 151726 91160 151740 91216
rect 151676 91156 151740 91160
rect 124444 90884 124508 90948
rect 244780 88980 244844 89044
rect 250300 66812 250364 66876
rect 253060 65452 253124 65516
rect 232452 61372 232516 61436
rect 267964 59876 268028 59940
rect 258580 57156 258644 57220
rect 226380 50220 226444 50284
rect 251772 43420 251836 43484
rect 262812 30908 262876 30972
rect 267780 24108 267844 24172
rect 228220 21252 228284 21316
rect 246252 3300 246316 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 99234 176600 99854 208338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 101995 177580 102061 177581
rect 101995 177516 101996 177580
rect 102060 177516 102061 177580
rect 101995 177515 102061 177516
rect 100707 177172 100773 177173
rect 100707 177108 100708 177172
rect 100772 177108 100773 177172
rect 100707 177107 100773 177108
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177107
rect 101998 175130 102058 177515
rect 102954 176600 103574 212058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 104571 176900 104637 176901
rect 104571 176836 104572 176900
rect 104636 176836 104637 176900
rect 104571 176835 104637 176836
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 176835
rect 105675 176764 105741 176765
rect 105675 176700 105676 176764
rect 105740 176700 105741 176764
rect 105675 176699 105741 176700
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 105678 175130 105738 176699
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 176764 110709 176765
rect 110643 176700 110644 176764
rect 110708 176700 110709 176764
rect 110643 176699 110709 176700
rect 112115 176764 112181 176765
rect 112115 176700 112116 176764
rect 112180 176700 112181 176764
rect 112115 176699 112181 176700
rect 113219 176764 113285 176765
rect 113219 176700 113220 176764
rect 113284 176700 113285 176764
rect 113219 176699 113285 176700
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 176699
rect 112118 175130 112178 176699
rect 113222 175130 113282 176699
rect 113514 176600 114134 186618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 116899 176764 116965 176765
rect 116899 176700 116900 176764
rect 116964 176700 116965 176764
rect 116899 176699 116965 176700
rect 114323 175676 114389 175677
rect 114323 175612 114324 175676
rect 114388 175612 114389 175676
rect 114323 175611 114389 175612
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175611
rect 116902 175130 116962 176699
rect 117234 176600 117854 190338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120763 177308 120829 177309
rect 120763 177244 120764 177308
rect 120828 177244 120829 177308
rect 120763 177243 120829 177244
rect 119475 176764 119541 176765
rect 119475 176700 119476 176764
rect 119540 176700 119541 176764
rect 119475 176699 119541 176700
rect 118371 175540 118437 175541
rect 118371 175476 118372 175540
rect 118436 175476 118437 175540
rect 118371 175475 118437 175476
rect 118374 175130 118434 175475
rect 119478 175130 119538 176699
rect 120766 175130 120826 177243
rect 120954 176600 121574 194058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 123155 177308 123221 177309
rect 123155 177244 123156 177308
rect 123220 177244 123221 177308
rect 123155 177243 123221 177244
rect 121867 175540 121933 175541
rect 121867 175476 121868 175540
rect 121932 175476 121933 175540
rect 121867 175475 121933 175476
rect 121870 175130 121930 175475
rect 123158 175130 123218 177243
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 124443 175676 124509 175677
rect 124443 175612 124444 175676
rect 124508 175612 124509 175676
rect 124443 175611 124509 175612
rect 124446 175130 124506 175611
rect 125734 175130 125794 176699
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 177580 130765 177581
rect 130699 177516 130700 177580
rect 130764 177516 130765 177580
rect 130699 177515 130765 177516
rect 129411 177308 129477 177309
rect 129411 177244 129412 177308
rect 129476 177244 129477 177308
rect 129411 177243 129477 177244
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 114326 175070 114428 175130
rect 116902 175070 117012 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115725 174996 115791 174997
rect 115725 174932 115726 174996
rect 115790 174932 115791 174996
rect 115725 174931 115791 174932
rect 115728 174494 115788 174931
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177243
rect 130702 175130 130762 177515
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 176764 132421 176765
rect 132355 176700 132356 176764
rect 132420 176700 132421 176764
rect 132355 176699 132421 176700
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 132358 175130 132418 176699
rect 133091 175676 133157 175677
rect 133091 175612 133092 175676
rect 133156 175612 133157 175676
rect 133091 175611 133157 175612
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 175611
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 166211 102780 166277 102781
rect 166211 102716 166212 102780
rect 166276 102716 166277 102780
rect 166211 102715 166277 102716
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91765 84394 94830
rect 84331 91764 84397 91765
rect 84331 91700 84332 91764
rect 84396 91700 84397 91764
rect 84331 91699 84397 91700
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 92445 85866 94830
rect 85803 92444 85869 92445
rect 85803 92380 85804 92444
rect 85868 92380 85869 92444
rect 85803 92379 85869 92380
rect 86726 91629 86786 94830
rect 86723 91628 86789 91629
rect 86723 91564 86724 91628
rect 86788 91564 86789 91628
rect 86723 91563 86789 91564
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 91221 88994 94830
rect 90222 91901 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 92445 91386 94830
rect 91323 92444 91389 92445
rect 91323 92380 91324 92444
rect 91388 92380 91389 92444
rect 91323 92379 91389 92380
rect 90219 91900 90285 91901
rect 90219 91836 90220 91900
rect 90284 91836 90285 91900
rect 90219 91835 90285 91836
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91221 96722 94830
rect 97214 91765 97274 94830
rect 97211 91764 97277 91765
rect 97211 91700 97212 91764
rect 97276 91700 97277 91764
rect 97211 91699 97277 91700
rect 98134 91221 98194 94830
rect 98502 92445 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 92444 98565 92445
rect 98499 92380 98500 92444
rect 98564 92380 98565 92444
rect 98499 92379 98565 92380
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100526 93533 100586 94830
rect 100523 93532 100589 93533
rect 100523 93468 100524 93532
rect 100588 93468 100589 93532
rect 100523 93467 100589 93468
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91765 101874 94830
rect 101811 91764 101877 91765
rect 101811 91700 101812 91764
rect 101876 91700 101877 91764
rect 101811 91699 101877 91700
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 91221 102794 93810
rect 103286 93530 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103286 93470 103714 93530
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 103654 92170 103714 93470
rect 104206 92445 104266 94830
rect 104574 93941 104634 94830
rect 104571 93940 104637 93941
rect 104571 93876 104572 93940
rect 104636 93876 104637 93940
rect 104571 93875 104637 93876
rect 105494 93533 105554 94830
rect 105491 93532 105557 93533
rect 105491 93468 105492 93532
rect 105556 93468 105557 93532
rect 105491 93467 105557 93468
rect 105678 92445 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 92445 106474 94830
rect 104203 92444 104269 92445
rect 104203 92380 104204 92444
rect 104268 92380 104269 92444
rect 104203 92379 104269 92380
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106411 92444 106477 92445
rect 106411 92380 106412 92444
rect 106476 92380 106477 92444
rect 106411 92379 106477 92380
rect 103835 92172 103901 92173
rect 103835 92170 103836 92172
rect 103654 92110 103836 92170
rect 103835 92108 103836 92110
rect 103900 92108 103901 92172
rect 103835 92107 103901 92108
rect 106782 91221 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 107702 91221 107762 94830
rect 108070 91221 108130 94830
rect 109064 94757 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 109472 94830 109602 94890
rect 109061 94756 109127 94757
rect 109061 94692 109062 94756
rect 109126 94692 109127 94756
rect 109061 94691 109127 94692
rect 109542 92445 109602 94830
rect 110094 94830 110212 94890
rect 110094 93261 110154 94830
rect 110696 94757 110756 95200
rect 111240 94890 111300 95200
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110693 94756 110759 94757
rect 110693 94692 110694 94756
rect 110758 94692 110759 94756
rect 110693 94691 110759 94692
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 109539 92444 109605 92445
rect 109539 92380 109540 92444
rect 109604 92380 109605 92444
rect 109539 92379 109605 92380
rect 106779 91220 106845 91221
rect 106779 91156 106780 91220
rect 106844 91156 106845 91220
rect 106779 91155 106845 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 111198 91221 111258 94830
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 113834 94890
rect 112302 91221 112362 94830
rect 113222 92445 113282 94830
rect 113774 93261 113834 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 114776 94830 114938 94890
rect 113771 93260 113837 93261
rect 113771 93196 113772 93260
rect 113836 93196 113837 93260
rect 113771 93195 113837 93196
rect 113219 92444 113285 92445
rect 113219 92380 113220 92444
rect 113284 92380 113285 92444
rect 113219 92379 113285 92380
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115430 92445 115490 94830
rect 115864 94757 115924 95200
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115861 94756 115927 94757
rect 115861 94692 115862 94756
rect 115926 94692 115927 94756
rect 115861 94691 115927 94692
rect 116718 93669 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 93668 116781 93669
rect 116715 93604 116716 93668
rect 116780 93604 116781 93668
rect 116715 93603 116781 93604
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 117086 91765 117146 94830
rect 117083 91764 117149 91765
rect 117083 91700 117084 91764
rect 117148 91700 117149 91764
rect 117083 91699 117149 91700
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92309 118066 94830
rect 118190 93533 118250 94830
rect 119400 94757 119460 95200
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119397 94756 119463 94757
rect 119397 94692 119398 94756
rect 119462 94692 119463 94756
rect 119397 94691 119463 94692
rect 118187 93532 118253 93533
rect 118187 93468 118188 93532
rect 118252 93468 118253 93532
rect 118187 93467 118253 93468
rect 118003 92308 118069 92309
rect 118003 92244 118004 92308
rect 118068 92244 118069 92308
rect 118003 92243 118069 92244
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120214 91221 120274 94830
rect 120582 92445 120642 94830
rect 120579 92444 120645 92445
rect 120579 92380 120580 92444
rect 120644 92380 120645 92444
rect 120579 92379 120645 92380
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91221 121746 94830
rect 122054 91221 122114 94830
rect 122974 92445 123034 94830
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122971 92444 123037 92445
rect 122971 92380 122972 92444
rect 123036 92380 123037 92444
rect 122971 92379 123037 92380
rect 123158 91221 123218 94830
rect 124078 91221 124138 94830
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124446 90949 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 93533 125426 94830
rect 125363 93532 125429 93533
rect 125363 93468 125364 93532
rect 125428 93468 125429 93532
rect 125363 93467 125429 93468
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126470 91629 126530 94830
rect 126467 91628 126533 91629
rect 126467 91564 126468 91628
rect 126532 91564 126533 91628
rect 126467 91563 126533 91564
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 127574 91221 127634 94830
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 124443 90948 124509 90949
rect 124443 90884 124444 90948
rect 124508 90884 124509 90948
rect 124443 90883 124509 90884
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 91221 133154 94830
rect 134382 91221 134442 94830
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151496 94754 151556 95200
rect 151632 94893 151692 95200
rect 151629 94892 151695 94893
rect 151629 94828 151630 94892
rect 151694 94828 151695 94892
rect 151629 94827 151695 94828
rect 151768 94754 151828 95200
rect 151494 94694 151556 94754
rect 151678 94694 151828 94754
rect 151904 94754 151964 95200
rect 151904 94694 152106 94754
rect 151494 93533 151554 94694
rect 151491 93532 151557 93533
rect 151491 93468 151492 93532
rect 151556 93468 151557 93532
rect 151491 93467 151557 93468
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151678 91221 151738 94694
rect 152046 93533 152106 94694
rect 152043 93532 152109 93533
rect 152043 93468 152044 93532
rect 152108 93468 152109 93532
rect 152043 93467 152109 93468
rect 151675 91220 151741 91221
rect 151675 91156 151676 91220
rect 151740 91156 151741 91220
rect 151675 91155 151741 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 92309 166274 102715
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166211 92308 166277 92309
rect 166211 92244 166212 92308
rect 166276 92244 166277 92308
rect 166211 92243 166277 92244
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 286182 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 286182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 213131 699820 213197 699821
rect 213131 699756 213132 699820
rect 213196 699756 213197 699820
rect 213131 699755 213197 699756
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 201355 284068 201421 284069
rect 201355 284004 201356 284068
rect 201420 284004 201421 284068
rect 201355 284003 201421 284004
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 198779 259452 198845 259453
rect 198779 259388 198780 259452
rect 198844 259388 198845 259452
rect 198779 259387 198845 259388
rect 197123 252244 197189 252245
rect 197123 252180 197124 252244
rect 197188 252180 197189 252244
rect 197123 252179 197189 252180
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 197126 95165 197186 252179
rect 198782 241501 198842 259387
rect 198779 241500 198845 241501
rect 198779 241436 198780 241500
rect 198844 241436 198845 241500
rect 198779 241435 198845 241436
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 201358 178125 201418 284003
rect 204851 283932 204917 283933
rect 204851 283868 204852 283932
rect 204916 283868 204917 283932
rect 204851 283867 204917 283868
rect 210739 283932 210805 283933
rect 210739 283868 210740 283932
rect 210804 283868 210805 283932
rect 210739 283867 210805 283868
rect 212395 283932 212461 283933
rect 212395 283868 212396 283932
rect 212460 283868 212461 283932
rect 212395 283867 212461 283868
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 204854 240141 204914 283867
rect 204851 240140 204917 240141
rect 204851 240076 204852 240140
rect 204916 240076 204917 240140
rect 204851 240075 204917 240076
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 201355 178124 201421 178125
rect 201355 178060 201356 178124
rect 201420 178060 201421 178124
rect 201355 178059 201421 178060
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 197123 95164 197189 95165
rect 197123 95100 197124 95164
rect 197188 95100 197189 95164
rect 197123 95099 197189 95100
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238182
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 210742 183021 210802 283867
rect 210954 212614 211574 238182
rect 212398 224229 212458 283867
rect 213134 238645 213194 699755
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 286182 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 286182 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 286182 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 228219 286108 228285 286109
rect 228219 286044 228220 286108
rect 228284 286044 228285 286108
rect 228219 286043 228285 286044
rect 244411 286108 244477 286109
rect 244411 286044 244412 286108
rect 244476 286044 244477 286108
rect 244411 286043 244477 286044
rect 220859 285700 220925 285701
rect 220859 285636 220860 285700
rect 220924 285636 220925 285700
rect 220859 285635 220925 285636
rect 218099 284068 218165 284069
rect 218099 284004 218100 284068
rect 218164 284004 218165 284068
rect 218099 284003 218165 284004
rect 217547 283932 217613 283933
rect 217547 283868 217548 283932
rect 217612 283868 217613 283932
rect 217547 283867 217613 283868
rect 213131 238644 213197 238645
rect 213131 238580 213132 238644
rect 213196 238580 213197 238644
rect 213131 238579 213197 238580
rect 212395 224228 212461 224229
rect 212395 224164 212396 224228
rect 212460 224164 212461 224228
rect 212395 224163 212461 224164
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210739 183020 210805 183021
rect 210739 182956 210740 183020
rect 210804 182956 210805 183020
rect 210739 182955 210805 182956
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 212058
rect 217550 180165 217610 283867
rect 218102 240141 218162 284003
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 218099 240140 218165 240141
rect 218099 240076 218100 240140
rect 218164 240076 218165 240140
rect 218099 240075 218165 240076
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217547 180164 217613 180165
rect 217547 180100 217548 180164
rect 217612 180100 217613 180164
rect 217547 180099 217613 180100
rect 217794 178000 218414 182898
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 220862 175949 220922 285635
rect 223435 283932 223501 283933
rect 223435 283868 223436 283932
rect 223500 283868 223501 283932
rect 223435 283867 223501 283868
rect 224171 283932 224237 283933
rect 224171 283868 224172 283932
rect 224236 283868 224237 283932
rect 224171 283867 224237 283868
rect 226195 283932 226261 283933
rect 226195 283868 226196 283932
rect 226260 283868 226261 283932
rect 226195 283867 226261 283868
rect 226379 283932 226445 283933
rect 226379 283868 226380 283932
rect 226444 283868 226445 283932
rect 226379 283867 226445 283868
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 223438 175949 223498 283867
rect 220859 175948 220925 175949
rect 220859 175884 220860 175948
rect 220924 175884 220925 175948
rect 220859 175883 220925 175884
rect 223435 175948 223501 175949
rect 223435 175884 223436 175948
rect 223500 175884 223501 175948
rect 223435 175883 223501 175884
rect 224174 175813 224234 283867
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 226198 177989 226258 283867
rect 226382 178805 226442 283867
rect 226379 178804 226445 178805
rect 226379 178740 226380 178804
rect 226444 178740 226445 178804
rect 226379 178739 226445 178740
rect 226195 177988 226261 177989
rect 226195 177924 226196 177988
rect 226260 177924 226261 177988
rect 226195 177923 226261 177924
rect 228222 177445 228282 286043
rect 233187 284340 233253 284341
rect 233187 284276 233188 284340
rect 233252 284276 233253 284340
rect 233187 284275 233253 284276
rect 231715 284068 231781 284069
rect 231715 284004 231716 284068
rect 231780 284004 231781 284068
rect 231715 284003 231781 284004
rect 229691 283932 229757 283933
rect 229691 283868 229692 283932
rect 229756 283868 229757 283932
rect 229691 283867 229757 283868
rect 231531 283932 231597 283933
rect 231531 283868 231532 283932
rect 231596 283868 231597 283932
rect 231531 283867 231597 283868
rect 229694 240141 229754 283867
rect 229691 240140 229757 240141
rect 229691 240076 229692 240140
rect 229756 240076 229757 240140
rect 229691 240075 229757 240076
rect 228954 230614 229574 238182
rect 231534 236061 231594 283867
rect 231531 236060 231597 236061
rect 231531 235996 231532 236060
rect 231596 235996 231597 236060
rect 231531 235995 231597 235996
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 231718 196077 231778 284003
rect 231899 208996 231965 208997
rect 231899 208932 231900 208996
rect 231964 208932 231965 208996
rect 231899 208931 231965 208932
rect 231715 196076 231781 196077
rect 231715 196012 231716 196076
rect 231780 196012 231781 196076
rect 231715 196011 231781 196012
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 229691 187100 229757 187101
rect 229691 187036 229692 187100
rect 229756 187036 229757 187100
rect 229691 187035 229757 187036
rect 228219 177444 228285 177445
rect 228219 177380 228220 177444
rect 228284 177380 228285 177444
rect 228219 177379 228285 177380
rect 229139 176764 229205 176765
rect 229139 176700 229140 176764
rect 229204 176700 229205 176764
rect 229139 176699 229205 176700
rect 224171 175812 224237 175813
rect 224171 175748 224172 175812
rect 224236 175748 224237 175812
rect 224171 175747 224237 175748
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 229142 137325 229202 176699
rect 229694 161669 229754 187035
rect 230427 182884 230493 182885
rect 230427 182820 230428 182884
rect 230492 182820 230493 182884
rect 230427 182819 230493 182820
rect 229691 161668 229757 161669
rect 229691 161604 229692 161668
rect 229756 161604 229757 161668
rect 229691 161603 229757 161604
rect 230430 156229 230490 182819
rect 230611 174996 230677 174997
rect 230611 174932 230612 174996
rect 230676 174932 230677 174996
rect 230611 174931 230677 174932
rect 230614 163437 230674 174931
rect 230611 163436 230677 163437
rect 230611 163372 230612 163436
rect 230676 163372 230677 163436
rect 230611 163371 230677 163372
rect 230427 156228 230493 156229
rect 230427 156164 230428 156228
rect 230492 156164 230493 156228
rect 230427 156163 230493 156164
rect 231902 151061 231962 208931
rect 232083 185740 232149 185741
rect 232083 185676 232084 185740
rect 232148 185676 232149 185740
rect 232083 185675 232149 185676
rect 231899 151060 231965 151061
rect 231899 150996 231900 151060
rect 231964 150996 231965 151060
rect 231899 150995 231965 150996
rect 230427 144804 230493 144805
rect 230427 144740 230428 144804
rect 230492 144740 230493 144804
rect 230427 144739 230493 144740
rect 230430 141677 230490 144739
rect 230427 141676 230493 141677
rect 230427 141612 230428 141676
rect 230492 141612 230493 141676
rect 230427 141611 230493 141612
rect 230979 141404 231045 141405
rect 230979 141340 230980 141404
rect 231044 141340 231045 141404
rect 230979 141339 231045 141340
rect 229691 140044 229757 140045
rect 229691 139980 229692 140044
rect 229756 139980 229757 140044
rect 229691 139979 229757 139980
rect 229139 137324 229205 137325
rect 229139 137260 229140 137324
rect 229204 137260 229205 137324
rect 229139 137259 229205 137260
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 229139 98292 229205 98293
rect 229139 98290 229140 98292
rect 228958 98230 229140 98290
rect 228958 97202 229018 98230
rect 229139 98228 229140 98230
rect 229204 98228 229205 98292
rect 229139 98227 229205 98228
rect 228222 97142 229018 97202
rect 229139 97204 229205 97205
rect 226379 95980 226445 95981
rect 226379 95916 226380 95980
rect 226444 95916 226445 95980
rect 226379 95915 226445 95916
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 226382 50285 226442 95915
rect 226379 50284 226445 50285
rect 226379 50220 226380 50284
rect 226444 50220 226445 50284
rect 226379 50219 226445 50220
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 228222 21317 228282 97142
rect 229139 97140 229140 97204
rect 229204 97140 229205 97204
rect 229139 97139 229205 97140
rect 229142 96930 229202 97139
rect 228958 96870 229202 96930
rect 228958 95981 229018 96870
rect 228955 95980 229021 95981
rect 228955 95916 228956 95980
rect 229020 95916 229021 95980
rect 228955 95915 229021 95916
rect 228954 86614 229574 94000
rect 229694 93941 229754 139979
rect 230982 127397 231042 141339
rect 232086 139229 232146 185675
rect 233190 147253 233250 284275
rect 244227 284068 244293 284069
rect 244227 284004 244228 284068
rect 244292 284004 244293 284068
rect 244227 284003 244293 284004
rect 244230 280530 244290 284003
rect 244046 280470 244290 280530
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 243491 246260 243557 246261
rect 243491 246196 243492 246260
rect 243556 246196 243557 246260
rect 243491 246195 243557 246196
rect 243494 238645 243554 246195
rect 244046 243810 244106 280470
rect 244414 277410 244474 286043
rect 244230 277350 244474 277410
rect 246954 284614 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 248459 291276 248525 291277
rect 248459 291212 248460 291276
rect 248524 291212 248525 291276
rect 248459 291211 248525 291212
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 244230 244221 244290 277350
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 244227 244220 244293 244221
rect 244227 244156 244228 244220
rect 244292 244156 244293 244220
rect 244227 244155 244293 244156
rect 244227 244084 244293 244085
rect 244227 244020 244228 244084
rect 244292 244020 244293 244084
rect 244227 244019 244293 244020
rect 244230 243810 244290 244019
rect 244046 243750 244290 243810
rect 245883 243540 245949 243541
rect 245883 243476 245884 243540
rect 245948 243476 245949 243540
rect 245883 243475 245949 243476
rect 245886 240277 245946 243475
rect 245883 240276 245949 240277
rect 245883 240212 245884 240276
rect 245948 240212 245949 240276
rect 245883 240211 245949 240212
rect 243491 238644 243557 238645
rect 243491 238580 243492 238644
rect 243556 238580 243557 238644
rect 243491 238579 243557 238580
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 237419 237420 237485 237421
rect 237419 237356 237420 237420
rect 237484 237356 237485 237420
rect 237419 237355 237485 237356
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 234659 184244 234725 184245
rect 234659 184180 234660 184244
rect 234724 184180 234725 184244
rect 234659 184179 234725 184180
rect 233371 177308 233437 177309
rect 233371 177244 233372 177308
rect 233436 177244 233437 177308
rect 233371 177243 233437 177244
rect 233187 147252 233253 147253
rect 233187 147188 233188 147252
rect 233252 147188 233253 147252
rect 233187 147187 233253 147188
rect 233374 145349 233434 177243
rect 233371 145348 233437 145349
rect 233371 145284 233372 145348
rect 233436 145284 233437 145348
rect 233371 145283 233437 145284
rect 234662 144805 234722 184179
rect 235794 165454 236414 200898
rect 236499 196076 236565 196077
rect 236499 196012 236500 196076
rect 236564 196012 236565 196076
rect 236499 196011 236565 196012
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 144804 234725 144805
rect 234659 144740 234660 144804
rect 234724 144740 234725 144804
rect 234659 144739 234725 144740
rect 232083 139228 232149 139229
rect 232083 139164 232084 139228
rect 232148 139164 232149 139228
rect 232083 139163 232149 139164
rect 231163 137324 231229 137325
rect 231163 137260 231164 137324
rect 231228 137260 231229 137324
rect 231163 137259 231229 137260
rect 230979 127396 231045 127397
rect 230979 127332 230980 127396
rect 231044 127332 231045 127396
rect 230979 127331 231045 127332
rect 230979 116652 231045 116653
rect 230979 116588 230980 116652
rect 231044 116588 231045 116652
rect 230979 116587 231045 116588
rect 229691 93940 229757 93941
rect 229691 93876 229692 93940
rect 229756 93876 229757 93940
rect 229691 93875 229757 93876
rect 230982 91765 231042 116587
rect 231166 115157 231226 137259
rect 232451 131612 232517 131613
rect 232451 131548 232452 131612
rect 232516 131548 232517 131612
rect 232451 131547 232517 131548
rect 231163 115156 231229 115157
rect 231163 115092 231164 115156
rect 231228 115092 231229 115156
rect 231163 115091 231229 115092
rect 230979 91764 231045 91765
rect 230979 91700 230980 91764
rect 231044 91700 231045 91764
rect 230979 91699 231045 91700
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 232454 61437 232514 131547
rect 235794 129454 236414 164898
rect 236502 139773 236562 196011
rect 236499 139772 236565 139773
rect 236499 139708 236500 139772
rect 236564 139708 236565 139772
rect 236499 139707 236565 139708
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 237422 114477 237482 237355
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 237603 181524 237669 181525
rect 237603 181460 237604 181524
rect 237668 181460 237669 181524
rect 237603 181459 237669 181460
rect 237606 138821 237666 181459
rect 238523 176084 238589 176085
rect 238523 176020 238524 176084
rect 238588 176020 238589 176084
rect 238523 176019 238589 176020
rect 238526 159629 238586 176019
rect 239514 169174 240134 204618
rect 243234 208894 243854 238182
rect 244227 234700 244293 234701
rect 244227 234636 244228 234700
rect 244292 234636 244293 234700
rect 244227 234635 244293 234636
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 240363 180028 240429 180029
rect 240363 179964 240364 180028
rect 240428 179964 240429 180028
rect 240363 179963 240429 179964
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238523 159628 238589 159629
rect 238523 159564 238524 159628
rect 238588 159564 238589 159628
rect 238523 159563 238589 159564
rect 237603 138820 237669 138821
rect 237603 138756 237604 138820
rect 237668 138756 237669 138820
rect 237603 138755 237669 138756
rect 239514 133174 240134 168618
rect 240366 153917 240426 179963
rect 241651 176492 241717 176493
rect 241651 176428 241652 176492
rect 241716 176428 241717 176492
rect 241651 176427 241717 176428
rect 240363 153916 240429 153917
rect 240363 153852 240364 153916
rect 240428 153852 240429 153916
rect 240363 153851 240429 153852
rect 241654 136373 241714 176427
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 244230 153781 244290 234635
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 245699 186964 245765 186965
rect 245699 186900 245700 186964
rect 245764 186900 245765 186964
rect 245699 186899 245765 186900
rect 244227 153780 244293 153781
rect 244227 153716 244228 153780
rect 244292 153716 244293 153780
rect 244227 153715 244293 153716
rect 245702 147797 245762 186899
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 245699 147796 245765 147797
rect 245699 147732 245700 147796
rect 245764 147732 245765 147796
rect 245699 147731 245765 147732
rect 246954 140614 247574 176058
rect 248462 142085 248522 291211
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 249747 283252 249813 283253
rect 249747 283188 249748 283252
rect 249812 283188 249813 283252
rect 249747 283187 249813 283188
rect 248643 248708 248709 248709
rect 248643 248644 248644 248708
rect 248708 248644 248709 248708
rect 248643 248643 248709 248644
rect 248646 143445 248706 248643
rect 249750 145621 249810 283187
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 249747 145620 249813 145621
rect 249747 145556 249748 145620
rect 249812 145556 249813 145620
rect 249747 145555 249813 145556
rect 248643 143444 248709 143445
rect 248643 143380 248644 143444
rect 248708 143380 248709 143444
rect 248643 143379 248709 143380
rect 248459 142084 248525 142085
rect 248459 142020 248460 142084
rect 248524 142020 248525 142084
rect 248459 142019 248525 142020
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246251 139636 246317 139637
rect 246251 139572 246252 139636
rect 246316 139572 246317 139636
rect 246251 139571 246317 139572
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 241651 136372 241717 136373
rect 241651 136308 241652 136372
rect 241716 136308 241717 136372
rect 241651 136307 241717 136308
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 237419 114476 237485 114477
rect 237419 114412 237420 114476
rect 237484 114412 237485 114476
rect 237419 114411 237485 114412
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 232451 61436 232517 61437
rect 232451 61372 232452 61436
rect 232516 61372 232517 61436
rect 232451 61371 232517 61372
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228219 21316 228285 21317
rect 228219 21252 228220 21316
rect 228284 21252 228285 21316
rect 228219 21251 228285 21252
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 100894 243854 136338
rect 244779 132020 244845 132021
rect 244779 131956 244780 132020
rect 244844 131956 244845 132020
rect 244779 131955 244845 131956
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 244782 89045 244842 131955
rect 244779 89044 244845 89045
rect 244779 88980 244780 89044
rect 244844 88980 244845 89044
rect 244779 88979 244845 88980
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 246254 3365 246314 139571
rect 246954 104614 247574 140058
rect 251771 119100 251837 119101
rect 251771 119036 251772 119100
rect 251836 119036 251837 119100
rect 251771 119035 251837 119036
rect 250299 113524 250365 113525
rect 250299 113460 250300 113524
rect 250364 113460 250365 113524
rect 250299 113459 250365 113460
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 250302 66877 250362 113459
rect 250299 66876 250365 66877
rect 250299 66812 250300 66876
rect 250364 66812 250365 66876
rect 250299 66811 250365 66812
rect 251774 43485 251834 119035
rect 253059 113932 253125 113933
rect 253059 113868 253060 113932
rect 253124 113868 253125 113932
rect 253059 113867 253125 113868
rect 253062 65517 253122 113867
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253059 65516 253125 65517
rect 253059 65452 253060 65516
rect 253124 65452 253125 65516
rect 253059 65451 253125 65452
rect 251771 43484 251837 43485
rect 251771 43420 251772 43484
rect 251836 43420 251837 43484
rect 251771 43419 251837 43420
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246251 3364 246317 3365
rect 246251 3300 246252 3364
rect 246316 3300 246317 3364
rect 246251 3299 246317 3300
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 258579 128892 258645 128893
rect 258579 128828 258580 128892
rect 258644 128828 258645 128892
rect 258579 128827 258645 128828
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 258582 57221 258642 128827
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 278819 288692 278885 288693
rect 278819 288628 278820 288692
rect 278884 288628 278885 288692
rect 278819 288627 278885 288628
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 274587 189684 274653 189685
rect 274587 189620 274588 189684
rect 274652 189620 274653 189684
rect 274587 189619 274653 189620
rect 274590 175813 274650 189619
rect 275514 178000 276134 204618
rect 278822 176490 278882 288627
rect 279234 280894 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 280291 287196 280357 287197
rect 280291 287132 280292 287196
rect 280356 287132 280357 287196
rect 280291 287131 280357 287132
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 178000 279854 208338
rect 280294 190470 280354 287131
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 285627 295356 285693 295357
rect 285627 295292 285628 295356
rect 285692 295292 285693 295356
rect 285627 295291 285693 295292
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 281579 279716 281645 279717
rect 281579 279652 281580 279716
rect 281644 279652 281645 279716
rect 281579 279651 281645 279652
rect 280110 190410 280354 190470
rect 278822 176430 279434 176490
rect 274587 175812 274653 175813
rect 274587 175748 274588 175812
rect 274652 175748 274653 175812
rect 274587 175747 274653 175748
rect 279187 175812 279253 175813
rect 279187 175748 279188 175812
rect 279252 175748 279253 175812
rect 279187 175747 279253 175748
rect 279190 171150 279250 175747
rect 279374 172141 279434 176430
rect 279371 172140 279437 172141
rect 279371 172076 279372 172140
rect 279436 172076 279437 172140
rect 279371 172075 279437 172076
rect 279190 171090 279434 171150
rect 279374 166837 279434 171090
rect 279371 166836 279437 166837
rect 279371 166772 279372 166836
rect 279436 166772 279437 166836
rect 279371 166771 279437 166772
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 280110 134061 280170 190410
rect 280291 185604 280357 185605
rect 280291 185540 280292 185604
rect 280356 185540 280357 185604
rect 280291 185539 280357 185540
rect 280294 151830 280354 185539
rect 281582 157861 281642 279651
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 284339 225588 284405 225589
rect 284339 225524 284340 225588
rect 284404 225524 284405 225588
rect 284339 225523 284405 225524
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 281763 191044 281829 191045
rect 281763 190980 281764 191044
rect 281828 190980 281829 191044
rect 281763 190979 281829 190980
rect 281766 174045 281826 190979
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 283787 176628 283853 176629
rect 283787 176564 283788 176628
rect 283852 176564 283853 176628
rect 283787 176563 283853 176564
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281763 174044 281829 174045
rect 281763 173980 281764 174044
rect 281828 173980 281829 174044
rect 281763 173979 281829 173980
rect 281579 157860 281645 157861
rect 281579 157796 281580 157860
rect 281644 157796 281645 157860
rect 281579 157795 281645 157796
rect 280294 151770 280538 151830
rect 280107 134060 280173 134061
rect 280107 133996 280108 134060
rect 280172 133996 280173 134060
rect 280107 133995 280173 133996
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 280478 129437 280538 151770
rect 282954 140614 283574 176058
rect 283790 163165 283850 176563
rect 283787 163164 283853 163165
rect 283787 163100 283788 163164
rect 283852 163100 283853 163164
rect 283787 163099 283853 163100
rect 284342 144805 284402 225523
rect 284523 181388 284589 181389
rect 284523 181324 284524 181388
rect 284588 181324 284589 181388
rect 284523 181323 284589 181324
rect 284339 144804 284405 144805
rect 284339 144740 284340 144804
rect 284404 144740 284405 144804
rect 284339 144739 284405 144740
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280475 129436 280541 129437
rect 280475 129372 280476 129436
rect 280540 129372 280541 129436
rect 280475 129371 280541 129372
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 267779 128484 267845 128485
rect 267779 128420 267780 128484
rect 267844 128420 267845 128484
rect 267779 128419 267845 128420
rect 267595 127940 267661 127941
rect 267595 127876 267596 127940
rect 267660 127876 267661 127940
rect 267595 127875 267661 127876
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 262811 115156 262877 115157
rect 262811 115092 262812 115156
rect 262876 115092 262877 115156
rect 262811 115091 262877 115092
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 258579 57220 258645 57221
rect 258579 57156 258580 57220
rect 258644 57156 258645 57220
rect 258579 57155 258645 57156
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 262814 30973 262874 115091
rect 264954 86614 265574 122058
rect 267598 94485 267658 127875
rect 267595 94484 267661 94485
rect 267595 94420 267596 94484
rect 267660 94420 267661 94484
rect 267595 94419 267661 94420
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 262811 30972 262877 30973
rect 262811 30908 262812 30972
rect 262876 30908 262877 30972
rect 262811 30907 262877 30908
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 267782 24173 267842 128419
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 282954 104614 283574 140058
rect 284526 138549 284586 181323
rect 285630 143173 285690 295291
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288387 288556 288453 288557
rect 288387 288492 288388 288556
rect 288452 288492 288453 288556
rect 288387 288491 288453 288492
rect 287099 284476 287165 284477
rect 287099 284412 287100 284476
rect 287164 284412 287165 284476
rect 287099 284411 287165 284412
rect 285811 177444 285877 177445
rect 285811 177380 285812 177444
rect 285876 177380 285877 177444
rect 285811 177379 285877 177380
rect 285627 143172 285693 143173
rect 285627 143108 285628 143172
rect 285692 143108 285693 143172
rect 285627 143107 285693 143108
rect 284523 138548 284589 138549
rect 284523 138484 284524 138548
rect 284588 138484 284589 138548
rect 284523 138483 284589 138484
rect 285814 104821 285874 177379
rect 287102 121821 287162 284411
rect 287283 192540 287349 192541
rect 287283 192476 287284 192540
rect 287348 192476 287349 192540
rect 287283 192475 287349 192476
rect 287099 121820 287165 121821
rect 287099 121756 287100 121820
rect 287164 121756 287165 121820
rect 287099 121755 287165 121756
rect 287286 106317 287346 192475
rect 288390 106453 288450 288491
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 288571 182884 288637 182885
rect 288571 182820 288572 182884
rect 288636 182820 288637 182884
rect 288571 182819 288637 182820
rect 288574 134197 288634 182819
rect 289794 147454 290414 182898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 295379 206276 295445 206277
rect 295379 206212 295380 206276
rect 295444 206212 295445 206276
rect 295379 206211 295445 206212
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 291147 177308 291213 177309
rect 291147 177244 291148 177308
rect 291212 177244 291213 177308
rect 291147 177243 291213 177244
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288571 134196 288637 134197
rect 288571 134132 288572 134196
rect 288636 134132 288637 134196
rect 288571 134131 288637 134132
rect 289794 111454 290414 146898
rect 291150 146437 291210 177243
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 291147 146436 291213 146437
rect 291147 146372 291148 146436
rect 291212 146372 291213 146436
rect 291147 146371 291213 146372
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 288387 106452 288453 106453
rect 288387 106388 288388 106452
rect 288452 106388 288453 106452
rect 288387 106387 288453 106388
rect 287283 106316 287349 106317
rect 287283 106252 287284 106316
rect 287348 106252 287349 106316
rect 287283 106251 287349 106252
rect 285811 104820 285877 104821
rect 285811 104756 285812 104820
rect 285876 104756 285877 104820
rect 285811 104755 285877 104756
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 267963 100196 268029 100197
rect 267963 100132 267964 100196
rect 268028 100132 268029 100196
rect 267963 100131 268029 100132
rect 267966 59941 268026 100131
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 267963 59940 268029 59941
rect 267963 59876 267964 59940
rect 268028 59876 268029 59940
rect 267963 59875 268029 59876
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 267779 24172 267845 24173
rect 267779 24108 267780 24172
rect 267844 24108 267845 24172
rect 267779 24107 267845 24108
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 295382 102237 295442 206211
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 295379 102236 295445 102237
rect 295379 102172 295380 102236
rect 295444 102172 295445 102236
rect 295379 102171 295445 102172
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 275513 128898 275749 129134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1643900835
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1643900835
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1643900835
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1643900835
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
