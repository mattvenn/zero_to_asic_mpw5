magic
tech sky130A
magscale 1 2
timestamp 1647523150
<< metal1 >>
rect 201494 703196 201500 703248
rect 201552 703236 201558 703248
rect 202782 703236 202788 703248
rect 201552 703208 202788 703236
rect 201552 703196 201558 703208
rect 202782 703196 202788 703208
rect 202840 703196 202846 703248
rect 95142 703128 95148 703180
rect 95200 703168 95206 703180
rect 332502 703168 332508 703180
rect 95200 703140 332508 703168
rect 95200 703128 95206 703140
rect 332502 703128 332508 703140
rect 332560 703128 332566 703180
rect 116578 703060 116584 703112
rect 116636 703100 116642 703112
rect 397454 703100 397460 703112
rect 116636 703072 397460 703100
rect 116636 703060 116642 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 76558 702992 76564 703044
rect 76616 703032 76622 703044
rect 364978 703032 364984 703044
rect 76616 703004 364984 703032
rect 76616 702992 76622 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 104802 702924 104808 702976
rect 104860 702964 104866 702976
rect 413646 702964 413652 702976
rect 104860 702936 413652 702964
rect 104860 702924 104866 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 113082 702856 113088 702908
rect 113140 702896 113146 702908
rect 462314 702896 462320 702908
rect 113140 702868 462320 702896
rect 113140 702856 113146 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 75178 702788 75184 702840
rect 75236 702828 75242 702840
rect 429838 702828 429844 702840
rect 75236 702800 429844 702828
rect 75236 702788 75242 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 110322 702720 110328 702772
rect 110380 702760 110386 702772
rect 478506 702760 478512 702772
rect 110380 702732 478512 702760
rect 110380 702720 110386 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 115842 702652 115848 702704
rect 115900 702692 115906 702704
rect 494790 702692 494796 702704
rect 115900 702664 494796 702692
rect 115900 702652 115906 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 111702 702584 111708 702636
rect 111760 702624 111766 702636
rect 559650 702624 559656 702636
rect 111760 702596 559656 702624
rect 111760 702584 111766 702596
rect 559650 702584 559656 702596
rect 559708 702584 559714 702636
rect 79318 702516 79324 702568
rect 79376 702556 79382 702568
rect 527174 702556 527180 702568
rect 79376 702528 527180 702556
rect 79376 702516 79382 702528
rect 527174 702516 527180 702528
rect 527232 702516 527238 702568
rect 68922 702448 68928 702500
rect 68980 702488 68986 702500
rect 543458 702488 543464 702500
rect 68980 702460 543464 702488
rect 68980 702448 68986 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 85574 700380 85580 700392
rect 8168 700352 85580 700380
rect 8168 700340 8174 700352
rect 85574 700340 85580 700352
rect 85632 700340 85638 700392
rect 97258 700340 97264 700392
rect 97316 700380 97322 700392
rect 154114 700380 154120 700392
rect 97316 700352 154120 700380
rect 97316 700340 97322 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 155218 700340 155224 700392
rect 155276 700380 155282 700392
rect 218974 700380 218980 700392
rect 155276 700352 218980 700380
rect 155276 700340 155282 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 235166 700312 235172 700324
rect 62080 700284 235172 700312
rect 62080 700272 62086 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 106274 698952 106280 698964
rect 24360 698924 106280 698952
rect 24360 698912 24366 698924
rect 106274 698912 106280 698924
rect 106332 698912 106338 698964
rect 57882 697552 57888 697604
rect 57940 697592 57946 697604
rect 170306 697592 170312 697604
rect 57940 697564 170312 697592
rect 57940 697552 57946 697564
rect 170306 697552 170312 697564
rect 170364 697552 170370 697604
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 69014 696940 69020 696992
rect 69072 696980 69078 696992
rect 580166 696980 580172 696992
rect 69072 696952 580172 696980
rect 69072 696940 69078 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 122742 683136 122748 683188
rect 122800 683176 122806 683188
rect 580166 683176 580172 683188
rect 122800 683148 580172 683176
rect 122800 683136 122806 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 57974 670732 57980 670744
rect 3568 670704 57980 670732
rect 3568 670692 3574 670704
rect 57974 670692 57980 670704
rect 58032 670692 58038 670744
rect 83458 670692 83464 670744
rect 83516 670732 83522 670744
rect 580166 670732 580172 670744
rect 83516 670704 580172 670732
rect 83516 670692 83522 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 658112 3516 658164
rect 3568 658152 3574 658164
rect 7558 658152 7564 658164
rect 3568 658124 7564 658152
rect 3568 658112 3574 658124
rect 7558 658112 7564 658124
rect 7616 658112 7622 658164
rect 128998 643084 129004 643136
rect 129056 643124 129062 643136
rect 580166 643124 580172 643136
rect 129056 643096 580172 643124
rect 129056 643084 129062 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 87598 618304 87604 618316
rect 3568 618276 87604 618304
rect 3568 618264 3574 618276
rect 87598 618264 87604 618276
rect 87656 618264 87662 618316
rect 411898 616836 411904 616888
rect 411956 616876 411962 616888
rect 580166 616876 580172 616888
rect 411956 616848 580172 616876
rect 411956 616836 411962 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 35158 605860 35164 605872
rect 3568 605832 35164 605860
rect 3568 605820 3574 605832
rect 35158 605820 35164 605832
rect 35216 605820 35222 605872
rect 68830 596776 68836 596828
rect 68888 596816 68894 596828
rect 136634 596816 136640 596828
rect 68888 596788 136640 596816
rect 68888 596776 68894 596788
rect 136634 596776 136640 596788
rect 136692 596776 136698 596828
rect 78030 595416 78036 595468
rect 78088 595456 78094 595468
rect 266354 595456 266360 595468
rect 78088 595428 266360 595456
rect 78088 595416 78094 595428
rect 266354 595416 266360 595428
rect 266412 595416 266418 595468
rect 40034 591268 40040 591320
rect 40092 591308 40098 591320
rect 55858 591308 55864 591320
rect 40092 591280 55864 591308
rect 40092 591268 40098 591280
rect 55858 591268 55864 591280
rect 55916 591268 55922 591320
rect 111610 590656 111616 590708
rect 111668 590696 111674 590708
rect 580166 590696 580172 590708
rect 111668 590668 580172 590696
rect 111668 590656 111674 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 68462 589908 68468 589960
rect 68520 589948 68526 589960
rect 97258 589948 97264 589960
rect 68520 589920 97264 589948
rect 68520 589908 68526 589920
rect 97258 589908 97264 589920
rect 97316 589908 97322 589960
rect 7558 588548 7564 588600
rect 7616 588588 7622 588600
rect 87322 588588 87328 588600
rect 7616 588560 87328 588588
rect 7616 588548 7622 588560
rect 87322 588548 87328 588560
rect 87380 588548 87386 588600
rect 87598 587868 87604 587920
rect 87656 587908 87662 587920
rect 95234 587908 95240 587920
rect 87656 587880 95240 587908
rect 87656 587868 87662 587880
rect 95234 587868 95240 587880
rect 95292 587868 95298 587920
rect 81710 587800 81716 587852
rect 81768 587840 81774 587852
rect 83458 587840 83464 587852
rect 81768 587812 83464 587840
rect 81768 587800 81774 587812
rect 83458 587800 83464 587812
rect 83516 587800 83522 587852
rect 3418 587120 3424 587172
rect 3476 587160 3482 587172
rect 53834 587160 53840 587172
rect 3476 587132 53840 587160
rect 3476 587120 3482 587132
rect 53834 587120 53840 587132
rect 53892 587120 53898 587172
rect 88334 587120 88340 587172
rect 88392 587160 88398 587172
rect 111794 587160 111800 587172
rect 88392 587132 111800 587160
rect 88392 587120 88398 587132
rect 111794 587120 111800 587132
rect 111852 587120 111858 587172
rect 133230 587120 133236 587172
rect 133288 587160 133294 587172
rect 155218 587160 155224 587172
rect 133288 587132 155224 587160
rect 133288 587120 133294 587132
rect 155218 587120 155224 587132
rect 155276 587120 155282 587172
rect 94130 586780 94136 586832
rect 94188 586820 94194 586832
rect 117498 586820 117504 586832
rect 94188 586792 117504 586820
rect 94188 586780 94194 586792
rect 117498 586780 117504 586792
rect 117556 586780 117562 586832
rect 91554 586712 91560 586764
rect 91612 586752 91618 586764
rect 123110 586752 123116 586764
rect 91612 586724 123116 586752
rect 91612 586712 91618 586724
rect 123110 586712 123116 586724
rect 123168 586712 123174 586764
rect 94866 586644 94872 586696
rect 94924 586684 94930 586696
rect 127066 586684 127072 586696
rect 94924 586656 127072 586684
rect 94924 586644 94930 586656
rect 127066 586644 127072 586656
rect 127124 586644 127130 586696
rect 46842 586576 46848 586628
rect 46900 586616 46906 586628
rect 85114 586616 85120 586628
rect 46900 586588 85120 586616
rect 46900 586576 46906 586588
rect 85114 586576 85120 586588
rect 85172 586576 85178 586628
rect 90266 586576 90272 586628
rect 90324 586616 90330 586628
rect 124306 586616 124312 586628
rect 90324 586588 124312 586616
rect 90324 586576 90330 586588
rect 124306 586576 124312 586588
rect 124364 586576 124370 586628
rect 41230 586508 41236 586560
rect 41288 586548 41294 586560
rect 80606 586548 80612 586560
rect 41288 586520 80612 586548
rect 41288 586508 41294 586520
rect 80606 586508 80612 586520
rect 80664 586508 80670 586560
rect 98730 586508 98736 586560
rect 98788 586548 98794 586560
rect 133230 586548 133236 586560
rect 98788 586520 133236 586548
rect 98788 586508 98794 586520
rect 133230 586508 133236 586520
rect 133288 586508 133294 586560
rect 69106 585760 69112 585812
rect 69164 585800 69170 585812
rect 282914 585800 282920 585812
rect 69164 585772 282920 585800
rect 69164 585760 69170 585772
rect 282914 585760 282920 585772
rect 282972 585760 282978 585812
rect 54478 585352 54484 585404
rect 54536 585392 54542 585404
rect 76558 585392 76564 585404
rect 54536 585364 76564 585392
rect 54536 585352 54542 585364
rect 76558 585352 76564 585364
rect 76616 585352 76622 585404
rect 95234 585352 95240 585404
rect 95292 585392 95298 585404
rect 95878 585392 95884 585404
rect 95292 585364 95884 585392
rect 95292 585352 95298 585364
rect 95878 585352 95884 585364
rect 95936 585392 95942 585404
rect 118694 585392 118700 585404
rect 95936 585364 118700 585392
rect 95936 585352 95942 585364
rect 118694 585352 118700 585364
rect 118752 585352 118758 585404
rect 52178 585284 52184 585336
rect 52236 585324 52242 585336
rect 78030 585324 78036 585336
rect 52236 585296 78036 585324
rect 52236 585284 52242 585296
rect 78030 585284 78036 585296
rect 78088 585284 78094 585336
rect 95142 585284 95148 585336
rect 95200 585324 95206 585336
rect 122834 585324 122840 585336
rect 95200 585296 122840 585324
rect 95200 585284 95206 585296
rect 122834 585284 122840 585296
rect 122892 585284 122898 585336
rect 34238 585216 34244 585268
rect 34296 585256 34302 585268
rect 72234 585256 72240 585268
rect 34296 585228 72240 585256
rect 34296 585216 34302 585228
rect 72234 585216 72240 585228
rect 72292 585216 72298 585268
rect 92290 585216 92296 585268
rect 92348 585256 92354 585268
rect 125594 585256 125600 585268
rect 92348 585228 125600 585256
rect 92348 585216 92354 585228
rect 125594 585216 125600 585228
rect 125652 585216 125658 585268
rect 46750 585148 46756 585200
rect 46808 585188 46814 585200
rect 85574 585188 85580 585200
rect 46808 585160 85580 585188
rect 46808 585148 46814 585160
rect 85574 585148 85580 585160
rect 85632 585148 85638 585200
rect 87322 585148 87328 585200
rect 87380 585188 87386 585200
rect 87506 585188 87512 585200
rect 87380 585160 87512 585188
rect 87380 585148 87386 585160
rect 87506 585148 87512 585160
rect 87564 585188 87570 585200
rect 121454 585188 121460 585200
rect 87564 585160 121460 585188
rect 87564 585148 87570 585160
rect 121454 585148 121460 585160
rect 121512 585148 121518 585200
rect 103146 584400 103152 584452
rect 103204 584440 103210 584452
rect 104802 584440 104808 584452
rect 103204 584412 104808 584440
rect 103204 584400 103210 584412
rect 104802 584400 104808 584412
rect 104860 584440 104866 584452
rect 116302 584440 116308 584452
rect 104860 584412 116308 584440
rect 104860 584400 104866 584412
rect 116302 584400 116308 584412
rect 116360 584400 116366 584452
rect 36998 584060 37004 584112
rect 37056 584100 37062 584112
rect 75454 584100 75460 584112
rect 37056 584072 75460 584100
rect 37056 584060 37062 584072
rect 75454 584060 75460 584072
rect 75512 584060 75518 584112
rect 77846 584060 77852 584112
rect 77904 584100 77910 584112
rect 79318 584100 79324 584112
rect 77904 584072 79324 584100
rect 77904 584060 77910 584072
rect 79318 584060 79324 584072
rect 79376 584060 79382 584112
rect 59262 583992 59268 584044
rect 59320 584032 59326 584044
rect 77864 584032 77892 584060
rect 59320 584004 77892 584032
rect 59320 583992 59326 584004
rect 101306 583992 101312 584044
rect 101364 584032 101370 584044
rect 113174 584032 113180 584044
rect 101364 584004 113180 584032
rect 101364 583992 101370 584004
rect 113174 583992 113180 584004
rect 113232 583992 113238 584044
rect 53558 583924 53564 583976
rect 53616 583964 53622 583976
rect 75086 583964 75092 583976
rect 53616 583936 75092 583964
rect 53616 583924 53622 583936
rect 75086 583924 75092 583936
rect 75144 583924 75150 583976
rect 101858 583924 101864 583976
rect 101916 583964 101922 583976
rect 114554 583964 114560 583976
rect 101916 583936 114560 583964
rect 101916 583924 101922 583936
rect 114554 583924 114560 583936
rect 114612 583924 114618 583976
rect 57698 583856 57704 583908
rect 57756 583896 57762 583908
rect 81434 583896 81440 583908
rect 57756 583868 81440 583896
rect 57756 583856 57762 583868
rect 81434 583856 81440 583868
rect 81492 583896 81498 583908
rect 81710 583896 81716 583908
rect 81492 583868 81716 583896
rect 81492 583856 81498 583868
rect 81710 583856 81716 583868
rect 81768 583856 81774 583908
rect 88978 583856 88984 583908
rect 89036 583896 89042 583908
rect 100754 583896 100760 583908
rect 89036 583868 100760 583896
rect 89036 583856 89042 583868
rect 100754 583856 100760 583868
rect 100812 583856 100818 583908
rect 105538 583856 105544 583908
rect 105596 583896 105602 583908
rect 118786 583896 118792 583908
rect 105596 583868 118792 583896
rect 105596 583856 105602 583868
rect 118786 583856 118792 583868
rect 118844 583856 118850 583908
rect 61746 583788 61752 583840
rect 61804 583828 61810 583840
rect 87690 583828 87696 583840
rect 61804 583800 87696 583828
rect 61804 583788 61810 583800
rect 87690 583788 87696 583800
rect 87748 583788 87754 583840
rect 96522 583788 96528 583840
rect 96580 583828 96586 583840
rect 110690 583828 110696 583840
rect 96580 583800 110696 583828
rect 96580 583788 96586 583800
rect 110690 583788 110696 583800
rect 110748 583788 110754 583840
rect 69198 583720 69204 583772
rect 69256 583760 69262 583772
rect 73338 583760 73344 583772
rect 69256 583732 73344 583760
rect 69256 583720 69262 583732
rect 73338 583720 73344 583732
rect 73396 583720 73402 583772
rect 97442 583720 97448 583772
rect 97500 583760 97506 583772
rect 124214 583760 124220 583772
rect 97500 583732 124220 583760
rect 97500 583720 97506 583732
rect 124214 583720 124220 583732
rect 124272 583720 124278 583772
rect 59998 582972 60004 583024
rect 60056 583012 60062 583024
rect 71866 583012 71872 583024
rect 60056 582984 71872 583012
rect 60056 582972 60062 582984
rect 71866 582972 71872 582984
rect 71924 582972 71930 583024
rect 100754 582972 100760 583024
rect 100812 583012 100818 583024
rect 124490 583012 124496 583024
rect 100812 582984 124496 583012
rect 100812 582972 100818 582984
rect 124490 582972 124496 582984
rect 124548 582972 124554 583024
rect 11698 582700 11704 582752
rect 11756 582740 11762 582752
rect 107654 582740 107660 582752
rect 11756 582712 107660 582740
rect 11756 582700 11762 582712
rect 107654 582700 107660 582712
rect 107712 582700 107718 582752
rect 55122 582632 55128 582684
rect 55180 582672 55186 582684
rect 78674 582672 78680 582684
rect 55180 582644 78680 582672
rect 55180 582632 55186 582644
rect 78674 582632 78680 582644
rect 78732 582632 78738 582684
rect 56318 582564 56324 582616
rect 56376 582604 56382 582616
rect 81894 582604 81900 582616
rect 56376 582576 81900 582604
rect 56376 582564 56382 582576
rect 81894 582564 81900 582576
rect 81952 582564 81958 582616
rect 89622 582564 89628 582616
rect 89680 582604 89686 582616
rect 118970 582604 118976 582616
rect 89680 582576 118976 582604
rect 89680 582564 89686 582576
rect 118970 582564 118976 582576
rect 119028 582564 119034 582616
rect 52086 582496 52092 582548
rect 52144 582536 52150 582548
rect 79318 582536 79324 582548
rect 52144 582508 79324 582536
rect 52144 582496 52150 582508
rect 79318 582496 79324 582508
rect 79376 582496 79382 582548
rect 99282 582496 99288 582548
rect 99340 582536 99346 582548
rect 129734 582536 129740 582548
rect 99340 582508 129740 582536
rect 99340 582496 99346 582508
rect 129734 582496 129740 582508
rect 129792 582496 129798 582548
rect 103882 582428 103888 582480
rect 103940 582468 103946 582480
rect 116118 582468 116124 582480
rect 103940 582440 116124 582468
rect 103940 582428 103946 582440
rect 116118 582428 116124 582440
rect 116176 582428 116182 582480
rect 68738 582360 68744 582412
rect 68796 582400 68802 582412
rect 386322 582400 386328 582412
rect 68796 582372 386328 582400
rect 68796 582360 68802 582372
rect 386322 582360 386328 582372
rect 386380 582360 386386 582412
rect 82722 581788 82728 581800
rect 74506 581760 82728 581788
rect 70394 581680 70400 581732
rect 70452 581720 70458 581732
rect 70946 581720 70952 581732
rect 70452 581692 70952 581720
rect 70452 581680 70458 581692
rect 70946 581680 70952 581692
rect 71004 581680 71010 581732
rect 43806 581272 43812 581324
rect 43864 581312 43870 581324
rect 67634 581312 67640 581324
rect 43864 581284 67640 581312
rect 43864 581272 43870 581284
rect 67634 581272 67640 581284
rect 67692 581272 67698 581324
rect 59078 581204 59084 581256
rect 59136 581244 59142 581256
rect 70394 581244 70400 581256
rect 59136 581216 70400 581244
rect 59136 581204 59142 581216
rect 70394 581204 70400 581216
rect 70452 581204 70458 581256
rect 57790 581136 57796 581188
rect 57848 581176 57854 581188
rect 74506 581176 74534 581760
rect 82722 581748 82728 581760
rect 82780 581748 82786 581800
rect 104986 581748 104992 581800
rect 105044 581788 105050 581800
rect 111978 581788 111984 581800
rect 105044 581760 111984 581788
rect 105044 581748 105050 581760
rect 111978 581748 111984 581760
rect 112036 581748 112042 581800
rect 76742 581680 76748 581732
rect 76800 581680 76806 581732
rect 100570 581680 100576 581732
rect 100628 581720 100634 581732
rect 100628 581692 103514 581720
rect 100628 581680 100634 581692
rect 57848 581148 74534 581176
rect 57848 581136 57854 581148
rect 50798 581068 50804 581120
rect 50856 581108 50862 581120
rect 76760 581108 76788 581680
rect 50856 581080 76788 581108
rect 50856 581068 50862 581080
rect 35618 581000 35624 581052
rect 35676 581040 35682 581052
rect 70486 581040 70492 581052
rect 35676 581012 70492 581040
rect 35676 581000 35682 581012
rect 70486 581000 70492 581012
rect 70544 581000 70550 581052
rect 103486 581040 103514 581692
rect 104434 581680 104440 581732
rect 104492 581720 104498 581732
rect 104492 581692 113174 581720
rect 104492 581680 104498 581692
rect 113146 581108 113174 581692
rect 123018 581108 123024 581120
rect 113146 581080 123024 581108
rect 123018 581068 123024 581080
rect 123076 581068 123082 581120
rect 121546 581040 121552 581052
rect 103486 581012 121552 581040
rect 121546 581000 121552 581012
rect 121604 581000 121610 581052
rect 39942 580252 39948 580304
rect 40000 580292 40006 580304
rect 67910 580292 67916 580304
rect 40000 580264 67916 580292
rect 40000 580252 40006 580264
rect 67910 580252 67916 580264
rect 67968 580252 67974 580304
rect 3234 579708 3240 579760
rect 3292 579748 3298 579760
rect 7558 579748 7564 579760
rect 3292 579720 7564 579748
rect 3292 579708 3298 579720
rect 7558 579708 7564 579720
rect 7616 579708 7622 579760
rect 108942 579640 108948 579692
rect 109000 579680 109006 579692
rect 120166 579680 120172 579692
rect 109000 579652 120172 579680
rect 109000 579640 109006 579652
rect 120166 579640 120172 579652
rect 120224 579640 120230 579692
rect 106734 578892 106740 578944
rect 106792 578932 106798 578944
rect 121638 578932 121644 578944
rect 106792 578904 121644 578932
rect 106792 578892 106798 578904
rect 121638 578892 121644 578904
rect 121696 578892 121702 578944
rect 59170 578280 59176 578332
rect 59228 578320 59234 578332
rect 67634 578320 67640 578332
rect 59228 578292 67640 578320
rect 59228 578280 59234 578292
rect 67634 578280 67640 578292
rect 67692 578280 67698 578332
rect 108850 578280 108856 578332
rect 108908 578320 108914 578332
rect 117314 578320 117320 578332
rect 108908 578292 117320 578320
rect 108908 578280 108914 578292
rect 117314 578280 117320 578292
rect 117372 578280 117378 578332
rect 108942 578212 108948 578264
rect 109000 578252 109006 578264
rect 134058 578252 134064 578264
rect 109000 578224 134064 578252
rect 109000 578212 109006 578224
rect 134058 578212 134064 578224
rect 134116 578212 134122 578264
rect 108206 578144 108212 578196
rect 108264 578184 108270 578196
rect 111702 578184 111708 578196
rect 108264 578156 111708 578184
rect 108264 578144 108270 578156
rect 111702 578144 111708 578156
rect 111760 578144 111766 578196
rect 386322 578144 386328 578196
rect 386380 578184 386386 578196
rect 579798 578184 579804 578196
rect 386380 578156 579804 578184
rect 386380 578144 386386 578156
rect 579798 578144 579804 578156
rect 579856 578144 579862 578196
rect 63218 576852 63224 576904
rect 63276 576892 63282 576904
rect 67634 576892 67640 576904
rect 63276 576864 67640 576892
rect 63276 576852 63282 576864
rect 67634 576852 67640 576864
rect 67692 576852 67698 576904
rect 108942 575560 108948 575612
rect 109000 575600 109006 575612
rect 126238 575600 126244 575612
rect 109000 575572 126244 575600
rect 109000 575560 109006 575572
rect 126238 575560 126244 575572
rect 126296 575560 126302 575612
rect 34422 575492 34428 575544
rect 34480 575532 34486 575544
rect 67634 575532 67640 575544
rect 34480 575504 67640 575532
rect 34480 575492 34486 575504
rect 67634 575492 67640 575504
rect 67692 575492 67698 575544
rect 108850 575492 108856 575544
rect 108908 575532 108914 575544
rect 129826 575532 129832 575544
rect 108908 575504 129832 575532
rect 108908 575492 108914 575504
rect 129826 575492 129832 575504
rect 129884 575492 129890 575544
rect 64598 574132 64604 574184
rect 64656 574172 64662 574184
rect 67726 574172 67732 574184
rect 64656 574144 67732 574172
rect 64656 574132 64662 574144
rect 67726 574132 67732 574144
rect 67784 574132 67790 574184
rect 53742 574064 53748 574116
rect 53800 574104 53806 574116
rect 67634 574104 67640 574116
rect 53800 574076 67640 574104
rect 53800 574064 53806 574076
rect 67634 574064 67640 574076
rect 67692 574064 67698 574116
rect 108942 573996 108948 574048
rect 109000 574036 109006 574048
rect 121914 574036 121920 574048
rect 109000 574008 121920 574036
rect 109000 573996 109006 574008
rect 121914 573996 121920 574008
rect 121972 573996 121978 574048
rect 121914 573316 121920 573368
rect 121972 573356 121978 573368
rect 122742 573356 122748 573368
rect 121972 573328 122748 573356
rect 121972 573316 121978 573328
rect 122742 573316 122748 573328
rect 122800 573356 122806 573368
rect 131758 573356 131764 573368
rect 122800 573328 131764 573356
rect 122800 573316 122806 573328
rect 131758 573316 131764 573328
rect 131816 573316 131822 573368
rect 108942 572840 108948 572892
rect 109000 572880 109006 572892
rect 113358 572880 113364 572892
rect 109000 572852 113364 572880
rect 109000 572840 109006 572852
rect 113358 572840 113364 572852
rect 113416 572840 113422 572892
rect 64690 572772 64696 572824
rect 64748 572812 64754 572824
rect 67726 572812 67732 572824
rect 64748 572784 67732 572812
rect 64748 572772 64754 572784
rect 67726 572772 67732 572784
rect 67784 572772 67790 572824
rect 107838 572772 107844 572824
rect 107896 572812 107902 572824
rect 110506 572812 110512 572824
rect 107896 572784 110512 572812
rect 107896 572772 107902 572784
rect 110506 572772 110512 572784
rect 110564 572772 110570 572824
rect 61838 572704 61844 572756
rect 61896 572744 61902 572756
rect 67634 572744 67640 572756
rect 61896 572716 67640 572744
rect 61896 572704 61902 572716
rect 67634 572704 67640 572716
rect 67692 572704 67698 572756
rect 105630 572296 105636 572348
rect 105688 572336 105694 572348
rect 109218 572336 109224 572348
rect 105688 572308 109224 572336
rect 105688 572296 105694 572308
rect 109218 572296 109224 572308
rect 109276 572296 109282 572348
rect 66162 571548 66168 571600
rect 66220 571588 66226 571600
rect 68278 571588 68284 571600
rect 66220 571560 68284 571588
rect 66220 571548 66226 571560
rect 68278 571548 68284 571560
rect 68336 571548 68342 571600
rect 108942 571344 108948 571396
rect 109000 571384 109006 571396
rect 128354 571384 128360 571396
rect 109000 571356 128360 571384
rect 109000 571344 109006 571356
rect 128354 571344 128360 571356
rect 128412 571344 128418 571396
rect 108850 569984 108856 570036
rect 108908 570024 108914 570036
rect 132494 570024 132500 570036
rect 108908 569996 132500 570024
rect 108908 569984 108914 569996
rect 132494 569984 132500 569996
rect 132552 569984 132558 570036
rect 39298 569916 39304 569968
rect 39356 569956 39362 569968
rect 67634 569956 67640 569968
rect 39356 569928 67640 569956
rect 39356 569916 39362 569928
rect 67634 569916 67640 569928
rect 67692 569916 67698 569968
rect 108942 569916 108948 569968
rect 109000 569956 109006 569968
rect 135346 569956 135352 569968
rect 109000 569928 135352 569956
rect 109000 569916 109006 569928
rect 135346 569916 135352 569928
rect 135404 569916 135410 569968
rect 64782 568624 64788 568676
rect 64840 568664 64846 568676
rect 67634 568664 67640 568676
rect 64840 568636 67640 568664
rect 64840 568624 64846 568636
rect 67634 568624 67640 568636
rect 67692 568624 67698 568676
rect 108942 568556 108948 568608
rect 109000 568596 109006 568608
rect 120074 568596 120080 568608
rect 109000 568568 120080 568596
rect 109000 568556 109006 568568
rect 120074 568556 120080 568568
rect 120132 568556 120138 568608
rect 108942 567536 108948 567588
rect 109000 567576 109006 567588
rect 114646 567576 114652 567588
rect 109000 567548 114652 567576
rect 109000 567536 109006 567548
rect 114646 567536 114652 567548
rect 114704 567536 114710 567588
rect 66070 567196 66076 567248
rect 66128 567236 66134 567248
rect 67634 567236 67640 567248
rect 66128 567208 67640 567236
rect 66128 567196 66134 567208
rect 67634 567196 67640 567208
rect 67692 567196 67698 567248
rect 108942 567196 108948 567248
rect 109000 567236 109006 567248
rect 115934 567236 115940 567248
rect 109000 567208 115940 567236
rect 109000 567196 109006 567208
rect 115934 567196 115940 567208
rect 115992 567196 115998 567248
rect 108850 565904 108856 565956
rect 108908 565944 108914 565956
rect 117406 565944 117412 565956
rect 108908 565916 117412 565944
rect 108908 565904 108914 565916
rect 117406 565904 117412 565916
rect 117464 565904 117470 565956
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 22738 565876 22744 565888
rect 3476 565848 22744 565876
rect 3476 565836 3482 565848
rect 22738 565836 22744 565848
rect 22796 565836 22802 565888
rect 108942 565836 108948 565888
rect 109000 565876 109006 565888
rect 125870 565876 125876 565888
rect 109000 565848 125876 565876
rect 109000 565836 109006 565848
rect 125870 565836 125876 565848
rect 125928 565836 125934 565888
rect 65978 564476 65984 564528
rect 66036 564516 66042 564528
rect 67726 564516 67732 564528
rect 66036 564488 67732 564516
rect 66036 564476 66042 564488
rect 67726 564476 67732 564488
rect 67784 564476 67790 564528
rect 49602 564408 49608 564460
rect 49660 564448 49666 564460
rect 67634 564448 67640 564460
rect 49660 564420 67640 564448
rect 49660 564408 49666 564420
rect 67634 564408 67640 564420
rect 67692 564408 67698 564460
rect 108942 564408 108948 564460
rect 109000 564448 109006 564460
rect 131022 564448 131028 564460
rect 109000 564420 131028 564448
rect 109000 564408 109006 564420
rect 131022 564408 131028 564420
rect 131080 564448 131086 564460
rect 413278 564448 413284 564460
rect 131080 564420 413284 564448
rect 131080 564408 131086 564420
rect 413278 564408 413284 564420
rect 413336 564408 413342 564460
rect 108942 563728 108948 563780
rect 109000 563768 109006 563780
rect 110322 563768 110328 563780
rect 109000 563740 110328 563768
rect 109000 563728 109006 563740
rect 110322 563728 110328 563740
rect 110380 563768 110386 563780
rect 136818 563768 136824 563780
rect 110380 563740 136824 563768
rect 110380 563728 110386 563740
rect 136818 563728 136824 563740
rect 136876 563728 136882 563780
rect 126238 563660 126244 563712
rect 126296 563700 126302 563712
rect 580166 563700 580172 563712
rect 126296 563672 580172 563700
rect 126296 563660 126302 563672
rect 580166 563660 580172 563672
rect 580224 563660 580230 563712
rect 61930 563116 61936 563168
rect 61988 563156 61994 563168
rect 67634 563156 67640 563168
rect 61988 563128 67640 563156
rect 61988 563116 61994 563128
rect 67634 563116 67640 563128
rect 67692 563116 67698 563168
rect 48130 563048 48136 563100
rect 48188 563088 48194 563100
rect 67726 563088 67732 563100
rect 48188 563060 67732 563088
rect 48188 563048 48194 563060
rect 67726 563048 67732 563060
rect 67784 563048 67790 563100
rect 60734 562980 60740 563032
rect 60792 563020 60798 563032
rect 62022 563020 62028 563032
rect 60792 562992 62028 563020
rect 60792 562980 60798 562992
rect 62022 562980 62028 562992
rect 62080 563020 62086 563032
rect 67634 563020 67640 563032
rect 62080 562992 67640 563020
rect 62080 562980 62086 562992
rect 67634 562980 67640 562992
rect 67692 562980 67698 563032
rect 52270 562300 52276 562352
rect 52328 562340 52334 562352
rect 60734 562340 60740 562352
rect 52328 562312 60740 562340
rect 52328 562300 52334 562312
rect 60734 562300 60740 562312
rect 60792 562300 60798 562352
rect 107654 560328 107660 560380
rect 107712 560368 107718 560380
rect 120258 560368 120264 560380
rect 107712 560340 120264 560368
rect 107712 560328 107718 560340
rect 120258 560328 120264 560340
rect 120316 560328 120322 560380
rect 50982 560260 50988 560312
rect 51040 560300 51046 560312
rect 67634 560300 67640 560312
rect 51040 560272 67640 560300
rect 51040 560260 51046 560272
rect 67634 560260 67640 560272
rect 67692 560260 67698 560312
rect 108942 560260 108948 560312
rect 109000 560300 109006 560312
rect 139486 560300 139492 560312
rect 109000 560272 139492 560300
rect 109000 560260 109006 560272
rect 139486 560260 139492 560272
rect 139544 560260 139550 560312
rect 128630 559512 128636 559564
rect 128688 559552 128694 559564
rect 201494 559552 201500 559564
rect 128688 559524 201500 559552
rect 128688 559512 128694 559524
rect 201494 559512 201500 559524
rect 201552 559512 201558 559564
rect 108850 558968 108856 559020
rect 108908 559008 108914 559020
rect 128630 559008 128636 559020
rect 108908 558980 128636 559008
rect 108908 558968 108914 558980
rect 128630 558968 128636 558980
rect 128688 558968 128694 559020
rect 45462 558900 45468 558952
rect 45520 558940 45526 558952
rect 67634 558940 67640 558952
rect 45520 558912 67640 558940
rect 45520 558900 45526 558912
rect 67634 558900 67640 558912
rect 67692 558900 67698 558952
rect 108942 558900 108948 558952
rect 109000 558940 109006 558952
rect 138106 558940 138112 558952
rect 109000 558912 138112 558940
rect 109000 558900 109006 558912
rect 138106 558900 138112 558912
rect 138164 558900 138170 558952
rect 108574 558016 108580 558068
rect 108632 558056 108638 558068
rect 111886 558056 111892 558068
rect 108632 558028 111892 558056
rect 108632 558016 108638 558028
rect 111886 558016 111892 558028
rect 111944 558016 111950 558068
rect 62758 557540 62764 557592
rect 62816 557580 62822 557592
rect 67634 557580 67640 557592
rect 62816 557552 67640 557580
rect 62816 557540 62822 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 108942 556520 108948 556572
rect 109000 556560 109006 556572
rect 113266 556560 113272 556572
rect 109000 556532 113272 556560
rect 109000 556520 109006 556532
rect 113266 556520 113272 556532
rect 113324 556520 113330 556572
rect 53650 556248 53656 556300
rect 53708 556288 53714 556300
rect 67726 556288 67732 556300
rect 53708 556260 67732 556288
rect 53708 556248 53714 556260
rect 67726 556248 67732 556260
rect 67784 556248 67790 556300
rect 43898 556180 43904 556232
rect 43956 556220 43962 556232
rect 67634 556220 67640 556232
rect 43956 556192 67640 556220
rect 43956 556180 43962 556192
rect 67634 556180 67640 556192
rect 67692 556180 67698 556232
rect 57882 556112 57888 556164
rect 57940 556152 57946 556164
rect 67726 556152 67732 556164
rect 57940 556124 67732 556152
rect 57940 556112 57946 556124
rect 67726 556112 67732 556124
rect 67784 556112 67790 556164
rect 48222 555432 48228 555484
rect 48280 555472 48286 555484
rect 57882 555472 57888 555484
rect 48280 555444 57888 555472
rect 48280 555432 48286 555444
rect 57882 555432 57888 555444
rect 57940 555432 57946 555484
rect 35710 554752 35716 554804
rect 35768 554792 35774 554804
rect 67634 554792 67640 554804
rect 35768 554764 67640 554792
rect 35768 554752 35774 554764
rect 67634 554752 67640 554764
rect 67692 554752 67698 554804
rect 109218 554752 109224 554804
rect 109276 554792 109282 554804
rect 115198 554792 115204 554804
rect 109276 554764 115204 554792
rect 109276 554752 109282 554764
rect 115198 554752 115204 554764
rect 115256 554752 115262 554804
rect 3142 554684 3148 554736
rect 3200 554724 3206 554736
rect 11698 554724 11704 554736
rect 3200 554696 11704 554724
rect 3200 554684 3206 554696
rect 11698 554684 11704 554696
rect 11756 554684 11762 554736
rect 108942 554004 108948 554056
rect 109000 554044 109006 554056
rect 111610 554044 111616 554056
rect 109000 554016 111616 554044
rect 109000 554004 109006 554016
rect 111610 554004 111616 554016
rect 111668 554044 111674 554056
rect 133966 554044 133972 554056
rect 111668 554016 133972 554044
rect 111668 554004 111674 554016
rect 133966 554004 133972 554016
rect 134024 554004 134030 554056
rect 57238 553392 57244 553444
rect 57296 553432 57302 553444
rect 67634 553432 67640 553444
rect 57296 553404 67640 553432
rect 57296 553392 57302 553404
rect 67634 553392 67640 553404
rect 67692 553392 67698 553444
rect 108942 553392 108948 553444
rect 109000 553432 109006 553444
rect 127250 553432 127256 553444
rect 109000 553404 127256 553432
rect 109000 553392 109006 553404
rect 127250 553392 127256 553404
rect 127308 553432 127314 553444
rect 128998 553432 129004 553444
rect 127308 553404 129004 553432
rect 127308 553392 127314 553404
rect 128998 553392 129004 553404
rect 129056 553392 129062 553444
rect 50890 552032 50896 552084
rect 50948 552072 50954 552084
rect 67634 552072 67640 552084
rect 50948 552044 67640 552072
rect 50948 552032 50954 552044
rect 67634 552032 67640 552044
rect 67692 552032 67698 552084
rect 108942 552032 108948 552084
rect 109000 552072 109006 552084
rect 136634 552072 136640 552084
rect 109000 552044 136640 552072
rect 109000 552032 109006 552044
rect 136634 552032 136640 552044
rect 136692 552032 136698 552084
rect 42702 550604 42708 550656
rect 42760 550644 42766 550656
rect 67634 550644 67640 550656
rect 42760 550616 67640 550644
rect 42760 550604 42766 550616
rect 67634 550604 67640 550616
rect 67692 550604 67698 550656
rect 108942 550604 108948 550656
rect 109000 550644 109006 550656
rect 131114 550644 131120 550656
rect 109000 550616 131120 550644
rect 109000 550604 109006 550616
rect 131114 550604 131120 550616
rect 131172 550604 131178 550656
rect 63402 549312 63408 549364
rect 63460 549352 63466 549364
rect 67634 549352 67640 549364
rect 63460 549324 67640 549352
rect 63460 549312 63466 549324
rect 67634 549312 67640 549324
rect 67692 549312 67698 549364
rect 108942 549312 108948 549364
rect 109000 549352 109006 549364
rect 139394 549352 139400 549364
rect 109000 549324 139400 549352
rect 109000 549312 109006 549324
rect 139394 549312 139400 549324
rect 139452 549312 139458 549364
rect 44082 549244 44088 549296
rect 44140 549284 44146 549296
rect 67726 549284 67732 549296
rect 44140 549256 67732 549284
rect 44140 549244 44146 549256
rect 67726 549244 67732 549256
rect 67784 549244 67790 549296
rect 108850 549244 108856 549296
rect 108908 549284 108914 549296
rect 140958 549284 140964 549296
rect 108908 549256 140964 549284
rect 108908 549244 108914 549256
rect 140958 549244 140964 549256
rect 141016 549244 141022 549296
rect 67266 549108 67272 549160
rect 67324 549148 67330 549160
rect 68370 549148 68376 549160
rect 67324 549120 68376 549148
rect 67324 549108 67330 549120
rect 68370 549108 68376 549120
rect 68428 549108 68434 549160
rect 107838 548360 107844 548412
rect 107896 548400 107902 548412
rect 110598 548400 110604 548412
rect 107896 548372 110604 548400
rect 107896 548360 107902 548372
rect 110598 548360 110604 548372
rect 110656 548360 110662 548412
rect 107654 548224 107660 548276
rect 107712 548264 107718 548276
rect 107838 548264 107844 548276
rect 107712 548236 107844 548264
rect 107712 548224 107718 548236
rect 107838 548224 107844 548236
rect 107896 548224 107902 548276
rect 41138 547884 41144 547936
rect 41196 547924 41202 547936
rect 67634 547924 67640 547936
rect 41196 547896 67640 547924
rect 41196 547884 41202 547896
rect 67634 547884 67640 547896
rect 67692 547884 67698 547936
rect 133782 547136 133788 547188
rect 133840 547176 133846 547188
rect 299474 547176 299480 547188
rect 133840 547148 299480 547176
rect 133840 547136 133846 547148
rect 299474 547136 299480 547148
rect 299532 547136 299538 547188
rect 63310 546524 63316 546576
rect 63368 546564 63374 546576
rect 67726 546564 67732 546576
rect 63368 546536 67732 546564
rect 63368 546524 63374 546536
rect 67726 546524 67732 546536
rect 67784 546524 67790 546576
rect 109678 546524 109684 546576
rect 109736 546564 109742 546576
rect 133138 546564 133144 546576
rect 109736 546536 133144 546564
rect 109736 546524 109742 546536
rect 133138 546524 133144 546536
rect 133196 546564 133202 546576
rect 133782 546564 133788 546576
rect 133196 546536 133788 546564
rect 133196 546524 133202 546536
rect 133782 546524 133788 546536
rect 133840 546524 133846 546576
rect 60642 546456 60648 546508
rect 60700 546496 60706 546508
rect 67634 546496 67640 546508
rect 60700 546468 67640 546496
rect 60700 546456 60706 546468
rect 67634 546456 67640 546468
rect 67692 546456 67698 546508
rect 108942 546456 108948 546508
rect 109000 546496 109006 546508
rect 142338 546496 142344 546508
rect 109000 546468 142344 546496
rect 109000 546456 109006 546468
rect 142338 546456 142344 546468
rect 142396 546456 142402 546508
rect 37182 545708 37188 545760
rect 37240 545748 37246 545760
rect 68738 545748 68744 545760
rect 37240 545720 68744 545748
rect 37240 545708 37246 545720
rect 68738 545708 68744 545720
rect 68796 545708 68802 545760
rect 108942 545708 108948 545760
rect 109000 545748 109006 545760
rect 115842 545748 115848 545760
rect 109000 545720 115848 545748
rect 109000 545708 109006 545720
rect 115842 545708 115848 545720
rect 115900 545748 115906 545760
rect 124398 545748 124404 545760
rect 115900 545720 124404 545748
rect 115900 545708 115906 545720
rect 124398 545708 124404 545720
rect 124456 545708 124462 545760
rect 108942 545096 108948 545148
rect 109000 545136 109006 545148
rect 135438 545136 135444 545148
rect 109000 545108 135444 545136
rect 109000 545096 109006 545108
rect 135438 545096 135444 545108
rect 135496 545096 135502 545148
rect 22738 544348 22744 544400
rect 22796 544388 22802 544400
rect 33134 544388 33140 544400
rect 22796 544360 33140 544388
rect 22796 544348 22802 544360
rect 33134 544348 33140 544360
rect 33192 544348 33198 544400
rect 108942 544348 108948 544400
rect 109000 544388 109006 544400
rect 113082 544388 113088 544400
rect 109000 544360 113088 544388
rect 109000 544348 109006 544360
rect 113082 544348 113088 544360
rect 113140 544388 113146 544400
rect 136726 544388 136732 544400
rect 113140 544360 136732 544388
rect 113140 544348 113146 544360
rect 136726 544348 136732 544360
rect 136784 544348 136790 544400
rect 38562 543804 38568 543856
rect 38620 543844 38626 543856
rect 67726 543844 67732 543856
rect 38620 543816 67732 543844
rect 38620 543804 38626 543816
rect 67726 543804 67732 543816
rect 67784 543804 67790 543856
rect 33134 543736 33140 543788
rect 33192 543776 33198 543788
rect 34330 543776 34336 543788
rect 33192 543748 34336 543776
rect 33192 543736 33198 543748
rect 34330 543736 34336 543748
rect 34388 543776 34394 543788
rect 67634 543776 67640 543788
rect 34388 543748 67640 543776
rect 34388 543736 34394 543748
rect 67634 543736 67640 543748
rect 67692 543736 67698 543788
rect 60550 542444 60556 542496
rect 60608 542484 60614 542496
rect 67634 542484 67640 542496
rect 60608 542456 67640 542484
rect 60608 542444 60614 542456
rect 67634 542444 67640 542456
rect 67692 542444 67698 542496
rect 49418 542376 49424 542428
rect 49476 542416 49482 542428
rect 68922 542416 68928 542428
rect 49476 542388 68928 542416
rect 49476 542376 49482 542388
rect 68922 542376 68928 542388
rect 68980 542376 68986 542428
rect 108942 542376 108948 542428
rect 109000 542416 109006 542428
rect 142154 542416 142160 542428
rect 109000 542388 142160 542416
rect 109000 542376 109006 542388
rect 142154 542376 142160 542388
rect 142212 542376 142218 542428
rect 109770 541628 109776 541680
rect 109828 541668 109834 541680
rect 580258 541668 580264 541680
rect 109828 541640 580264 541668
rect 109828 541628 109834 541640
rect 580258 541628 580264 541640
rect 580316 541628 580322 541680
rect 62022 540948 62028 541000
rect 62080 540988 62086 541000
rect 67634 540988 67640 541000
rect 62080 540960 67640 540988
rect 62080 540948 62086 540960
rect 67634 540948 67640 540960
rect 67692 540948 67698 541000
rect 108942 540948 108948 541000
rect 109000 540988 109006 541000
rect 140774 540988 140780 541000
rect 109000 540960 140780 540988
rect 109000 540948 109006 540960
rect 140774 540948 140780 540960
rect 140832 540948 140838 541000
rect 41322 539656 41328 539708
rect 41380 539696 41386 539708
rect 59998 539696 60004 539708
rect 41380 539668 60004 539696
rect 41380 539656 41386 539668
rect 59998 539656 60004 539668
rect 60056 539656 60062 539708
rect 37090 539588 37096 539640
rect 37148 539628 37154 539640
rect 67634 539628 67640 539640
rect 37148 539600 67640 539628
rect 37148 539588 37154 539600
rect 67634 539588 67640 539600
rect 67692 539588 67698 539640
rect 4798 539520 4804 539572
rect 4856 539560 4862 539572
rect 99006 539560 99012 539572
rect 4856 539532 99012 539560
rect 4856 539520 4862 539532
rect 99006 539520 99012 539532
rect 99064 539520 99070 539572
rect 57974 539452 57980 539504
rect 58032 539492 58038 539504
rect 91278 539492 91284 539504
rect 58032 539464 91284 539492
rect 58032 539452 58038 539464
rect 91278 539452 91284 539464
rect 91336 539452 91342 539504
rect 99190 539044 99196 539096
rect 99248 539084 99254 539096
rect 111978 539084 111984 539096
rect 99248 539056 111984 539084
rect 99248 539044 99254 539056
rect 111978 539044 111984 539056
rect 112036 539044 112042 539096
rect 99006 538976 99012 539028
rect 99064 539016 99070 539028
rect 122926 539016 122932 539028
rect 99064 538988 122932 539016
rect 99064 538976 99070 538988
rect 122926 538976 122932 538988
rect 122984 538976 122990 539028
rect 95142 538908 95148 538960
rect 95200 538948 95206 538960
rect 121638 538948 121644 538960
rect 95200 538920 121644 538948
rect 95200 538908 95206 538920
rect 121638 538908 121644 538920
rect 121696 538908 121702 538960
rect 61746 538840 61752 538892
rect 61804 538880 61810 538892
rect 82998 538880 83004 538892
rect 61804 538852 83004 538880
rect 61804 538840 61810 538852
rect 82998 538840 83004 538852
rect 83056 538840 83062 538892
rect 88058 538840 88064 538892
rect 88116 538880 88122 538892
rect 122098 538880 122104 538892
rect 88116 538852 122104 538880
rect 88116 538840 88122 538852
rect 122098 538840 122104 538852
rect 122156 538880 122162 538892
rect 411898 538880 411904 538892
rect 122156 538852 411904 538880
rect 122156 538840 122162 538852
rect 411898 538840 411904 538852
rect 411956 538840 411962 538892
rect 413278 538840 413284 538892
rect 413336 538880 413342 538892
rect 580902 538880 580908 538892
rect 413336 538852 580908 538880
rect 413336 538840 413342 538852
rect 580902 538840 580908 538852
rect 580960 538840 580966 538892
rect 57514 538568 57520 538620
rect 57572 538608 57578 538620
rect 57974 538608 57980 538620
rect 57572 538580 57980 538608
rect 57572 538568 57578 538580
rect 57974 538568 57980 538580
rect 58032 538568 58038 538620
rect 7558 538160 7564 538212
rect 7616 538200 7622 538212
rect 98362 538200 98368 538212
rect 7616 538172 98368 538200
rect 7616 538160 7622 538172
rect 98362 538160 98368 538172
rect 98420 538160 98426 538212
rect 103514 538160 103520 538212
rect 103572 538200 103578 538212
rect 109678 538200 109684 538212
rect 103572 538172 109684 538200
rect 103572 538160 103578 538172
rect 109678 538160 109684 538172
rect 109736 538160 109742 538212
rect 59998 538092 60004 538144
rect 60056 538132 60062 538144
rect 73890 538132 73896 538144
rect 60056 538104 73896 538132
rect 60056 538092 60062 538104
rect 73890 538092 73896 538104
rect 73948 538092 73954 538144
rect 94498 538092 94504 538144
rect 94556 538132 94562 538144
rect 104710 538132 104716 538144
rect 94556 538104 104716 538132
rect 94556 538092 94562 538104
rect 104710 538092 104716 538104
rect 104768 538092 104774 538144
rect 102226 537752 102232 537804
rect 102284 537792 102290 537804
rect 127158 537792 127164 537804
rect 102284 537764 127164 537792
rect 102284 537752 102290 537764
rect 127158 537752 127164 537764
rect 127216 537752 127222 537804
rect 95786 537684 95792 537736
rect 95844 537724 95850 537736
rect 121730 537724 121736 537736
rect 95844 537696 121736 537724
rect 95844 537684 95850 537696
rect 121730 537684 121736 537696
rect 121788 537684 121794 537736
rect 59078 537616 59084 537668
rect 59136 537656 59142 537668
rect 69750 537656 69756 537668
rect 59136 537628 69756 537656
rect 59136 537616 59142 537628
rect 69750 537616 69756 537628
rect 69808 537616 69814 537668
rect 85482 537616 85488 537668
rect 85540 537656 85546 537668
rect 98638 537656 98644 537668
rect 85540 537628 98644 537656
rect 85540 537616 85546 537628
rect 98638 537616 98644 537628
rect 98696 537616 98702 537668
rect 102870 537616 102876 537668
rect 102928 537656 102934 537668
rect 132586 537656 132592 537668
rect 102928 537628 132592 537656
rect 102928 537616 102934 537628
rect 132586 537616 132592 537628
rect 132644 537616 132650 537668
rect 52362 537548 52368 537600
rect 52420 537588 52426 537600
rect 82906 537588 82912 537600
rect 52420 537560 82912 537588
rect 52420 537548 52426 537560
rect 82906 537548 82912 537560
rect 82964 537548 82970 537600
rect 98362 537548 98368 537600
rect 98420 537588 98426 537600
rect 128538 537588 128544 537600
rect 98420 537560 128544 537588
rect 98420 537548 98426 537560
rect 128538 537548 128544 537560
rect 128596 537548 128602 537600
rect 57790 537480 57796 537532
rect 57848 537520 57854 537532
rect 74718 537520 74724 537532
rect 57848 537492 74724 537520
rect 57848 537480 57854 537492
rect 74718 537480 74724 537492
rect 74776 537480 74782 537532
rect 116578 537520 116584 537532
rect 84166 537492 116584 537520
rect 80330 537412 80336 537464
rect 80388 537452 80394 537464
rect 81434 537452 81440 537464
rect 80388 537424 81440 537452
rect 80388 537412 80394 537424
rect 81434 537412 81440 537424
rect 81492 537452 81498 537464
rect 84166 537452 84194 537492
rect 116578 537480 116584 537492
rect 116636 537480 116642 537532
rect 81492 537424 84194 537452
rect 81492 537412 81498 537424
rect 83458 536800 83464 536852
rect 83516 536840 83522 536852
rect 84838 536840 84844 536852
rect 83516 536812 84844 536840
rect 83516 536800 83522 536812
rect 84838 536800 84844 536812
rect 84896 536800 84902 536852
rect 35158 536732 35164 536784
rect 35216 536772 35222 536784
rect 106090 536772 106096 536784
rect 35216 536744 106096 536772
rect 35216 536732 35222 536744
rect 106090 536732 106096 536744
rect 106148 536732 106154 536784
rect 111794 536528 111800 536580
rect 111852 536568 111858 536580
rect 114738 536568 114744 536580
rect 111852 536540 114744 536568
rect 111852 536528 111858 536540
rect 114738 536528 114744 536540
rect 114796 536528 114802 536580
rect 38470 536052 38476 536104
rect 38528 536092 38534 536104
rect 71314 536092 71320 536104
rect 38528 536064 71320 536092
rect 38528 536052 38534 536064
rect 71314 536052 71320 536064
rect 71372 536052 71378 536104
rect 106090 536052 106096 536104
rect 106148 536092 106154 536104
rect 134150 536092 134156 536104
rect 106148 536064 134156 536092
rect 106148 536052 106154 536064
rect 134150 536052 134156 536064
rect 134208 536052 134214 536104
rect 71038 534964 71044 535016
rect 71096 535004 71102 535016
rect 79686 535004 79692 535016
rect 71096 534976 79692 535004
rect 71096 534964 71102 534976
rect 79686 534964 79692 534976
rect 79744 534964 79750 535016
rect 101950 534964 101956 535016
rect 102008 535004 102014 535016
rect 107930 535004 107936 535016
rect 102008 534976 107936 535004
rect 102008 534964 102014 534976
rect 107930 534964 107936 534976
rect 107988 534964 107994 535016
rect 56410 534896 56416 534948
rect 56468 534936 56474 534948
rect 75178 534936 75184 534948
rect 56468 534908 75184 534936
rect 56468 534896 56474 534908
rect 75178 534896 75184 534908
rect 75236 534896 75242 534948
rect 97810 534896 97816 534948
rect 97868 534936 97874 534948
rect 116118 534936 116124 534948
rect 97868 534908 116124 534936
rect 97868 534896 97874 534908
rect 116118 534896 116124 534908
rect 116176 534896 116182 534948
rect 42610 534828 42616 534880
rect 42668 534868 42674 534880
rect 73246 534868 73252 534880
rect 42668 534840 73252 534868
rect 42668 534828 42674 534840
rect 73246 534828 73252 534840
rect 73304 534828 73310 534880
rect 89990 534828 89996 534880
rect 90048 534868 90054 534880
rect 111978 534868 111984 534880
rect 90048 534840 111984 534868
rect 90048 534828 90054 534840
rect 111978 534828 111984 534840
rect 112036 534828 112042 534880
rect 50706 534760 50712 534812
rect 50764 534800 50770 534812
rect 83550 534800 83556 534812
rect 50764 534772 83556 534800
rect 50764 534760 50770 534772
rect 83550 534760 83556 534772
rect 83608 534760 83614 534812
rect 95050 534760 95056 534812
rect 95108 534800 95114 534812
rect 121546 534800 121552 534812
rect 95108 534772 121552 534800
rect 95108 534760 95114 534772
rect 121546 534760 121552 534772
rect 121604 534760 121610 534812
rect 45278 534692 45284 534744
rect 45336 534732 45342 534744
rect 78398 534732 78404 534744
rect 45336 534704 78404 534732
rect 45336 534692 45342 534704
rect 78398 534692 78404 534704
rect 78456 534692 78462 534744
rect 93854 534692 93860 534744
rect 93912 534732 93918 534744
rect 125778 534732 125784 534744
rect 93912 534704 125784 534732
rect 93912 534692 93918 534704
rect 125778 534692 125784 534704
rect 125836 534692 125842 534744
rect 97074 532176 97080 532228
rect 97132 532216 97138 532228
rect 109218 532216 109224 532228
rect 97132 532188 109224 532216
rect 97132 532176 97138 532188
rect 109218 532176 109224 532188
rect 109276 532176 109282 532228
rect 93762 532108 93768 532160
rect 93820 532148 93826 532160
rect 117498 532148 117504 532160
rect 93820 532120 117504 532148
rect 93820 532108 93826 532120
rect 117498 532108 117504 532120
rect 117556 532108 117562 532160
rect 87414 532040 87420 532092
rect 87472 532080 87478 532092
rect 111794 532080 111800 532092
rect 87472 532052 111800 532080
rect 87472 532040 87478 532052
rect 111794 532040 111800 532052
rect 111852 532040 111858 532092
rect 92566 531972 92572 532024
rect 92624 532012 92630 532024
rect 121638 532012 121644 532024
rect 92624 531984 121644 532012
rect 92624 531972 92630 531984
rect 121638 531972 121644 531984
rect 121696 531972 121702 532024
rect 49326 529252 49332 529304
rect 49384 529292 49390 529304
rect 71958 529292 71964 529304
rect 49384 529264 71964 529292
rect 49384 529252 49390 529264
rect 71958 529252 71964 529264
rect 72016 529252 72022 529304
rect 46566 529184 46572 529236
rect 46624 529224 46630 529236
rect 77110 529224 77116 529236
rect 46624 529196 77116 529224
rect 46624 529184 46630 529196
rect 77110 529184 77116 529196
rect 77168 529184 77174 529236
rect 106918 528612 106924 528624
rect 106246 528584 106924 528612
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 106246 528544 106274 528584
rect 106918 528572 106924 528584
rect 106976 528612 106982 528624
rect 116210 528612 116216 528624
rect 106976 528584 116216 528612
rect 106976 528572 106982 528584
rect 116210 528572 116216 528584
rect 116268 528572 116274 528624
rect 3200 528516 106274 528544
rect 3200 528504 3206 528516
rect 39758 525784 39764 525836
rect 39816 525824 39822 525836
rect 39816 525796 64874 525824
rect 39816 525784 39822 525796
rect 64846 525756 64874 525796
rect 68922 525756 68928 525768
rect 64846 525728 68928 525756
rect 68922 525716 68928 525728
rect 68980 525756 68986 525768
rect 579798 525756 579804 525768
rect 68980 525728 579804 525756
rect 68980 525716 68986 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 58618 512184 58624 512236
rect 58676 512224 58682 512236
rect 59170 512224 59176 512236
rect 58676 512196 59176 512224
rect 58676 512184 58682 512196
rect 59170 512184 59176 512196
rect 59228 512184 59234 512236
rect 59170 511980 59176 512032
rect 59228 512020 59234 512032
rect 59228 511992 68968 512020
rect 59228 511980 59234 511992
rect 68940 511952 68968 511992
rect 580166 511952 580172 511964
rect 68940 511924 580172 511952
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 84194 500216 84200 500268
rect 84252 500256 84258 500268
rect 117498 500256 117504 500268
rect 84252 500228 117504 500256
rect 84252 500216 84258 500228
rect 117498 500216 117504 500228
rect 117556 500216 117562 500268
rect 96430 497632 96436 497684
rect 96488 497672 96494 497684
rect 118878 497672 118884 497684
rect 96488 497644 118884 497672
rect 96488 497632 96494 497644
rect 118878 497632 118884 497644
rect 118936 497632 118942 497684
rect 57606 497564 57612 497616
rect 57664 497604 57670 497616
rect 77754 497604 77760 497616
rect 57664 497576 77760 497604
rect 57664 497564 57670 497576
rect 77754 497564 77760 497576
rect 77812 497564 77818 497616
rect 86770 497564 86776 497616
rect 86828 497604 86834 497616
rect 117590 497604 117596 497616
rect 86828 497576 117596 497604
rect 86828 497564 86834 497576
rect 117590 497564 117596 497576
rect 117648 497564 117654 497616
rect 45370 497496 45376 497548
rect 45428 497536 45434 497548
rect 72602 497536 72608 497548
rect 45428 497508 72608 497536
rect 45428 497496 45434 497508
rect 72602 497496 72608 497508
rect 72660 497496 72666 497548
rect 91278 497536 91284 497548
rect 84166 497508 91284 497536
rect 4798 497428 4804 497480
rect 4856 497468 4862 497480
rect 84166 497468 84194 497508
rect 91278 497496 91284 497508
rect 91336 497536 91342 497548
rect 124214 497536 124220 497548
rect 91336 497508 124220 497536
rect 91336 497496 91342 497508
rect 124214 497496 124220 497508
rect 124272 497536 124278 497548
rect 135254 497536 135260 497548
rect 124272 497508 135260 497536
rect 124272 497496 124278 497508
rect 135254 497496 135260 497508
rect 135312 497496 135318 497548
rect 4856 497440 84194 497468
rect 4856 497428 4862 497440
rect 92566 497428 92572 497480
rect 92624 497468 92630 497480
rect 133230 497468 133236 497480
rect 92624 497440 133236 497468
rect 92624 497428 92630 497440
rect 133230 497428 133236 497440
rect 133288 497468 133294 497480
rect 138014 497468 138020 497480
rect 133288 497440 138020 497468
rect 133288 497428 133294 497440
rect 138014 497428 138020 497440
rect 138072 497428 138078 497480
rect 118786 496748 118792 496800
rect 118844 496788 118850 496800
rect 119062 496788 119068 496800
rect 118844 496760 119068 496788
rect 118844 496748 118850 496760
rect 119062 496748 119068 496760
rect 119120 496748 119126 496800
rect 56226 496204 56232 496256
rect 56284 496244 56290 496256
rect 81434 496244 81440 496256
rect 56284 496216 81440 496244
rect 56284 496204 56290 496216
rect 81434 496204 81440 496216
rect 81492 496204 81498 496256
rect 89622 496136 89628 496188
rect 89680 496176 89686 496188
rect 123110 496176 123116 496188
rect 89680 496148 123116 496176
rect 89680 496136 89686 496148
rect 123110 496136 123116 496148
rect 123168 496176 123174 496188
rect 124214 496176 124220 496188
rect 123168 496148 124220 496176
rect 123168 496136 123174 496148
rect 124214 496136 124220 496148
rect 124272 496136 124278 496188
rect 56318 496068 56324 496120
rect 56376 496108 56382 496120
rect 75822 496108 75828 496120
rect 56376 496080 75828 496108
rect 56376 496068 56382 496080
rect 75822 496068 75828 496080
rect 75880 496108 75886 496120
rect 81434 496108 81440 496120
rect 75880 496080 81440 496108
rect 75880 496068 75886 496080
rect 81434 496068 81440 496080
rect 81492 496068 81498 496120
rect 88058 496068 88064 496120
rect 88116 496108 88122 496120
rect 127066 496108 127072 496120
rect 88116 496080 127072 496108
rect 88116 496068 88122 496080
rect 127066 496068 127072 496080
rect 127124 496108 127130 496120
rect 133874 496108 133880 496120
rect 127124 496080 133880 496108
rect 127124 496068 127130 496080
rect 133874 496068 133880 496080
rect 133932 496068 133938 496120
rect 81434 495456 81440 495508
rect 81492 495496 81498 495508
rect 110414 495496 110420 495508
rect 81492 495468 110420 495496
rect 81492 495456 81498 495468
rect 110414 495456 110420 495468
rect 110472 495456 110478 495508
rect 52086 494844 52092 494896
rect 52144 494884 52150 494896
rect 73246 494884 73252 494896
rect 52144 494856 73252 494884
rect 52144 494844 52150 494856
rect 73246 494844 73252 494856
rect 73304 494844 73310 494896
rect 98638 494844 98644 494896
rect 98696 494884 98702 494896
rect 112070 494884 112076 494896
rect 98696 494856 112076 494884
rect 98696 494844 98702 494856
rect 112070 494844 112076 494856
rect 112128 494844 112134 494896
rect 118786 494884 118792 494896
rect 113146 494856 118792 494884
rect 49510 494776 49516 494828
rect 49568 494816 49574 494828
rect 74718 494816 74724 494828
rect 49568 494788 74724 494816
rect 49568 494776 49574 494788
rect 74718 494776 74724 494788
rect 74776 494816 74782 494828
rect 76098 494816 76104 494828
rect 74776 494788 76104 494816
rect 74776 494776 74782 494788
rect 76098 494776 76104 494788
rect 76156 494776 76162 494828
rect 82906 494776 82912 494828
rect 82964 494816 82970 494828
rect 113146 494816 113174 494856
rect 118786 494844 118792 494856
rect 118844 494844 118850 494896
rect 123202 494816 123208 494828
rect 82964 494788 113174 494816
rect 116872 494788 123208 494816
rect 82964 494776 82970 494788
rect 3510 494708 3516 494760
rect 3568 494748 3574 494760
rect 82814 494748 82820 494760
rect 3568 494720 82820 494748
rect 3568 494708 3574 494720
rect 82814 494708 82820 494720
rect 82872 494708 82878 494760
rect 97718 494708 97724 494760
rect 97776 494748 97782 494760
rect 102134 494748 102140 494760
rect 97776 494720 102140 494748
rect 97776 494708 97782 494720
rect 102134 494708 102140 494720
rect 102192 494708 102198 494760
rect 114554 494748 114560 494760
rect 109006 494720 114560 494748
rect 95786 494640 95792 494692
rect 95844 494680 95850 494692
rect 109006 494680 109034 494720
rect 114554 494708 114560 494720
rect 114612 494748 114618 494760
rect 116872 494748 116900 494788
rect 123202 494776 123208 494788
rect 123260 494776 123266 494828
rect 114612 494720 116900 494748
rect 114612 494708 114618 494720
rect 118786 494708 118792 494760
rect 118844 494748 118850 494760
rect 118970 494748 118976 494760
rect 118844 494720 118976 494748
rect 118844 494708 118850 494720
rect 118970 494708 118976 494720
rect 119028 494748 119034 494760
rect 130010 494748 130016 494760
rect 119028 494720 130016 494748
rect 119028 494708 119034 494720
rect 130010 494708 130016 494720
rect 130068 494708 130074 494760
rect 95844 494652 109034 494680
rect 95844 494640 95850 494652
rect 85482 494368 85488 494420
rect 85540 494408 85546 494420
rect 89622 494408 89628 494420
rect 85540 494380 89628 494408
rect 85540 494368 85546 494380
rect 89622 494368 89628 494380
rect 89680 494368 89686 494420
rect 80974 494096 80980 494148
rect 81032 494136 81038 494148
rect 121454 494136 121460 494148
rect 81032 494108 121460 494136
rect 81032 494096 81038 494108
rect 121454 494096 121460 494108
rect 121512 494096 121518 494148
rect 41230 494028 41236 494080
rect 41288 494068 41294 494080
rect 74534 494068 74540 494080
rect 41288 494040 74540 494068
rect 41288 494028 41294 494040
rect 74534 494028 74540 494040
rect 74592 494028 74598 494080
rect 76650 494028 76656 494080
rect 76708 494068 76714 494080
rect 120350 494068 120356 494080
rect 76708 494040 120356 494068
rect 76708 494028 76714 494040
rect 120350 494028 120356 494040
rect 120408 494028 120414 494080
rect 82814 493960 82820 494012
rect 82872 494000 82878 494012
rect 83550 494000 83556 494012
rect 82872 493972 83556 494000
rect 82872 493960 82878 493972
rect 83550 493960 83556 493972
rect 83608 494000 83614 494012
rect 124306 494000 124312 494012
rect 83608 493972 124312 494000
rect 83608 493960 83614 493972
rect 124306 493960 124312 493972
rect 124364 494000 124370 494012
rect 130102 494000 130108 494012
rect 124364 493972 130108 494000
rect 124364 493960 124370 493972
rect 130102 493960 130108 493972
rect 130160 493960 130166 494012
rect 129734 493892 129740 493944
rect 129792 493932 129798 493944
rect 131206 493932 131212 493944
rect 129792 493904 131212 493932
rect 129792 493892 129798 493904
rect 131206 493892 131212 493904
rect 131264 493892 131270 493944
rect 90266 493416 90272 493468
rect 90324 493456 90330 493468
rect 110690 493456 110696 493468
rect 90324 493428 110696 493456
rect 90324 493416 90330 493428
rect 110690 493416 110696 493428
rect 110748 493416 110754 493468
rect 54754 493348 54760 493400
rect 54812 493388 54818 493400
rect 59262 493388 59268 493400
rect 54812 493360 59268 493388
rect 54812 493348 54818 493360
rect 59262 493348 59268 493360
rect 59320 493388 59326 493400
rect 68002 493388 68008 493400
rect 59320 493360 68008 493388
rect 59320 493348 59326 493360
rect 68002 493348 68008 493360
rect 68060 493348 68066 493400
rect 91922 493348 91928 493400
rect 91980 493388 91986 493400
rect 95142 493388 95148 493400
rect 91980 493360 95148 493388
rect 91980 493348 91986 493360
rect 95142 493348 95148 493360
rect 95200 493388 95206 493400
rect 116026 493388 116032 493400
rect 95200 493360 116032 493388
rect 95200 493348 95206 493360
rect 116026 493348 116032 493360
rect 116084 493348 116090 493400
rect 43990 493280 43996 493332
rect 44048 493320 44054 493332
rect 50798 493320 50804 493332
rect 44048 493292 50804 493320
rect 44048 493280 44054 493292
rect 50798 493280 50804 493292
rect 50856 493320 50862 493332
rect 70302 493320 70308 493332
rect 50856 493292 70308 493320
rect 50856 493280 50862 493292
rect 70302 493280 70308 493292
rect 70360 493280 70366 493332
rect 93210 493280 93216 493332
rect 93268 493320 93274 493332
rect 129734 493320 129740 493332
rect 93268 493292 129740 493320
rect 93268 493280 93274 493292
rect 129734 493280 129740 493292
rect 129792 493280 129798 493332
rect 57698 492872 57704 492924
rect 57756 492912 57762 492924
rect 74994 492912 75000 492924
rect 57756 492884 75000 492912
rect 57756 492872 57762 492884
rect 74994 492872 75000 492884
rect 75052 492872 75058 492924
rect 52086 492844 52092 492856
rect 51460 492816 52092 492844
rect 46842 492600 46848 492652
rect 46900 492640 46906 492652
rect 51460 492640 51488 492816
rect 52086 492804 52092 492816
rect 52144 492844 52150 492856
rect 79318 492844 79324 492856
rect 52144 492816 79324 492844
rect 52144 492804 52150 492816
rect 79318 492804 79324 492816
rect 79376 492804 79382 492856
rect 59262 492736 59268 492788
rect 59320 492776 59326 492788
rect 90266 492776 90272 492788
rect 59320 492748 90272 492776
rect 59320 492736 59326 492748
rect 90266 492736 90272 492748
rect 90324 492736 90330 492788
rect 92474 492736 92480 492788
rect 92532 492776 92538 492788
rect 93762 492776 93768 492788
rect 92532 492748 93768 492776
rect 92532 492736 92538 492748
rect 93762 492736 93768 492748
rect 93820 492776 93826 492788
rect 114554 492776 114560 492788
rect 93820 492748 114560 492776
rect 93820 492736 93826 492748
rect 114554 492736 114560 492748
rect 114612 492736 114618 492788
rect 54938 492668 54944 492720
rect 54996 492708 55002 492720
rect 580350 492708 580356 492720
rect 54996 492680 56640 492708
rect 54996 492668 55002 492680
rect 46900 492612 51488 492640
rect 56612 492640 56640 492680
rect 64846 492680 580356 492708
rect 57238 492640 57244 492652
rect 56612 492612 57244 492640
rect 46900 492600 46906 492612
rect 57238 492600 57244 492612
rect 57296 492640 57302 492652
rect 64846 492640 64874 492680
rect 580350 492668 580356 492680
rect 580408 492668 580414 492720
rect 57296 492612 64874 492640
rect 57296 492600 57302 492612
rect 87414 492600 87420 492652
rect 87472 492640 87478 492652
rect 92474 492640 92480 492652
rect 87472 492612 92480 492640
rect 87472 492600 87478 492612
rect 92474 492600 92480 492612
rect 92532 492600 92538 492652
rect 46658 492464 46664 492516
rect 46716 492504 46722 492516
rect 48038 492504 48044 492516
rect 46716 492476 48044 492504
rect 46716 492464 46722 492476
rect 48038 492464 48044 492476
rect 48096 492464 48102 492516
rect 93302 492124 93308 492176
rect 93360 492164 93366 492176
rect 102226 492164 102232 492176
rect 93360 492136 102232 492164
rect 93360 492124 93366 492136
rect 102226 492124 102232 492136
rect 102284 492124 102290 492176
rect 53282 492056 53288 492108
rect 53340 492096 53346 492108
rect 54478 492096 54484 492108
rect 53340 492068 54484 492096
rect 53340 492056 53346 492068
rect 54478 492056 54484 492068
rect 54536 492096 54542 492108
rect 70026 492096 70032 492108
rect 54536 492068 70032 492096
rect 54536 492056 54542 492068
rect 70026 492056 70032 492068
rect 70084 492056 70090 492108
rect 97902 492056 97908 492108
rect 97960 492096 97966 492108
rect 111058 492096 111064 492108
rect 97960 492068 111064 492096
rect 97960 492056 97966 492068
rect 111058 492056 111064 492068
rect 111116 492056 111122 492108
rect 53466 491988 53472 492040
rect 53524 492028 53530 492040
rect 55122 492028 55128 492040
rect 53524 492000 55128 492028
rect 53524 491988 53530 492000
rect 55122 491988 55128 492000
rect 55180 492028 55186 492040
rect 72234 492028 72240 492040
rect 55180 492000 72240 492028
rect 55180 491988 55186 492000
rect 72234 491988 72240 492000
rect 72292 491988 72298 492040
rect 97074 491988 97080 492040
rect 97132 492028 97138 492040
rect 116302 492028 116308 492040
rect 97132 492000 116308 492028
rect 97132 491988 97138 492000
rect 116302 491988 116308 492000
rect 116360 492028 116366 492040
rect 116360 492000 122834 492028
rect 116360 491988 116366 492000
rect 48038 491920 48044 491972
rect 48096 491960 48102 491972
rect 78030 491960 78036 491972
rect 48096 491932 78036 491960
rect 48096 491920 48102 491932
rect 78030 491920 78036 491932
rect 78088 491920 78094 491972
rect 81618 491920 81624 491972
rect 81676 491960 81682 491972
rect 82998 491960 83004 491972
rect 81676 491932 83004 491960
rect 81676 491920 81682 491932
rect 82998 491920 83004 491932
rect 83056 491960 83062 491972
rect 113450 491960 113456 491972
rect 83056 491932 113456 491960
rect 83056 491920 83062 491932
rect 113450 491920 113456 491932
rect 113508 491920 113514 491972
rect 122806 491960 122834 492000
rect 143534 491960 143540 491972
rect 122806 491932 143540 491960
rect 143534 491920 143540 491932
rect 143592 491920 143598 491972
rect 96430 491784 96436 491836
rect 96488 491824 96494 491836
rect 97902 491824 97908 491836
rect 96488 491796 97908 491824
rect 96488 491784 96494 491796
rect 97902 491784 97908 491796
rect 97960 491784 97966 491836
rect 68002 491648 68008 491700
rect 68060 491688 68066 491700
rect 71130 491688 71136 491700
rect 68060 491660 71136 491688
rect 68060 491648 68066 491660
rect 71130 491648 71136 491660
rect 71188 491648 71194 491700
rect 86402 491580 86408 491632
rect 86460 491620 86466 491632
rect 100662 491620 100668 491632
rect 86460 491592 100668 491620
rect 86460 491580 86466 491592
rect 100662 491580 100668 491592
rect 100720 491580 100726 491632
rect 82262 491512 82268 491564
rect 82320 491552 82326 491564
rect 109126 491552 109132 491564
rect 82320 491524 109132 491552
rect 82320 491512 82326 491524
rect 109126 491512 109132 491524
rect 109184 491512 109190 491564
rect 52178 491444 52184 491496
rect 52236 491484 52242 491496
rect 71774 491484 71780 491496
rect 52236 491456 71780 491484
rect 52236 491444 52242 491456
rect 71774 491444 71780 491456
rect 71832 491444 71838 491496
rect 89990 491376 89996 491428
rect 90048 491416 90054 491428
rect 92842 491416 92848 491428
rect 90048 491388 92848 491416
rect 90048 491376 90054 491388
rect 92842 491376 92848 491388
rect 92900 491376 92906 491428
rect 99650 491376 99656 491428
rect 99708 491416 99714 491428
rect 118786 491416 118792 491428
rect 99708 491388 118792 491416
rect 99708 491376 99714 491388
rect 118786 491376 118792 491388
rect 118844 491416 118850 491428
rect 119062 491416 119068 491428
rect 118844 491388 119068 491416
rect 118844 491376 118850 491388
rect 119062 491376 119068 491388
rect 119120 491376 119126 491428
rect 46750 491308 46756 491360
rect 46808 491348 46814 491360
rect 80054 491348 80060 491360
rect 46808 491320 80060 491348
rect 46808 491308 46814 491320
rect 80054 491308 80060 491320
rect 80112 491308 80118 491360
rect 100662 491240 100668 491292
rect 100720 491280 100726 491292
rect 125594 491280 125600 491292
rect 100720 491252 125600 491280
rect 100720 491240 100726 491252
rect 125594 491240 125600 491252
rect 125652 491240 125658 491292
rect 109126 491172 109132 491224
rect 109184 491212 109190 491224
rect 123110 491212 123116 491224
rect 109184 491184 123116 491212
rect 109184 491172 109190 491184
rect 123110 491172 123116 491184
rect 123168 491212 123174 491224
rect 124490 491212 124496 491224
rect 123168 491184 124496 491212
rect 123168 491172 123174 491184
rect 124490 491172 124496 491184
rect 124548 491212 124554 491224
rect 125502 491212 125508 491224
rect 124548 491184 125508 491212
rect 124548 491172 124554 491184
rect 125502 491172 125508 491184
rect 125560 491172 125566 491224
rect 101858 491104 101864 491156
rect 101916 491144 101922 491156
rect 109310 491144 109316 491156
rect 101916 491116 109316 491144
rect 101916 491104 101922 491116
rect 109310 491104 109316 491116
rect 109368 491104 109374 491156
rect 60366 490764 60372 490816
rect 60424 490804 60430 490816
rect 86126 490804 86132 490816
rect 60424 490776 86132 490804
rect 60424 490764 60430 490776
rect 86126 490764 86132 490776
rect 86184 490764 86190 490816
rect 54846 490696 54852 490748
rect 54904 490736 54910 490748
rect 83458 490736 83464 490748
rect 54904 490708 83464 490736
rect 54904 490696 54910 490708
rect 83458 490696 83464 490708
rect 83516 490696 83522 490748
rect 47946 490628 47952 490680
rect 48004 490668 48010 490680
rect 79042 490668 79048 490680
rect 48004 490640 79048 490668
rect 48004 490628 48010 490640
rect 79042 490628 79048 490640
rect 79100 490628 79106 490680
rect 88978 490628 88984 490680
rect 89036 490668 89042 490680
rect 101306 490668 101312 490680
rect 89036 490640 101312 490668
rect 89036 490628 89042 490640
rect 101306 490628 101312 490640
rect 101364 490628 101370 490680
rect 35802 490560 35808 490612
rect 35860 490600 35866 490612
rect 36998 490600 37004 490612
rect 35860 490572 37004 490600
rect 35860 490560 35866 490572
rect 36998 490560 37004 490572
rect 37056 490600 37062 490612
rect 69750 490600 69756 490612
rect 37056 490572 69756 490600
rect 37056 490560 37062 490572
rect 69750 490560 69756 490572
rect 69808 490560 69814 490612
rect 94130 490560 94136 490612
rect 94188 490600 94194 490612
rect 95050 490600 95056 490612
rect 94188 490572 95056 490600
rect 94188 490560 94194 490572
rect 95050 490560 95056 490572
rect 95108 490600 95114 490612
rect 109678 490600 109684 490612
rect 95108 490572 109684 490600
rect 95108 490560 95114 490572
rect 109678 490560 109684 490572
rect 109736 490560 109742 490612
rect 125502 490560 125508 490612
rect 125560 490600 125566 490612
rect 580258 490600 580264 490612
rect 125560 490572 580264 490600
rect 125560 490560 125566 490572
rect 580258 490560 580264 490572
rect 580316 490560 580322 490612
rect 125594 490288 125600 490340
rect 125652 490328 125658 490340
rect 127066 490328 127072 490340
rect 125652 490300 127072 490328
rect 125652 490288 125658 490300
rect 127066 490288 127072 490300
rect 127124 490288 127130 490340
rect 86954 489880 86960 489932
rect 87012 489920 87018 489932
rect 101858 489920 101864 489932
rect 87012 489892 101864 489920
rect 87012 489880 87018 489892
rect 101858 489880 101864 489892
rect 101916 489880 101922 489932
rect 118786 489880 118792 489932
rect 118844 489920 118850 489932
rect 124306 489920 124312 489932
rect 118844 489892 124312 489920
rect 118844 489880 118850 489892
rect 124306 489880 124312 489892
rect 124364 489880 124370 489932
rect 69842 489812 69848 489864
rect 69900 489852 69906 489864
rect 70854 489852 70860 489864
rect 69900 489824 70860 489852
rect 69900 489812 69906 489824
rect 70854 489812 70860 489824
rect 70912 489812 70918 489864
rect 98730 489812 98736 489864
rect 98788 489852 98794 489864
rect 99282 489852 99288 489864
rect 98788 489824 99288 489852
rect 98788 489812 98794 489824
rect 99282 489812 99288 489824
rect 99340 489812 99346 489864
rect 101306 489812 101312 489864
rect 101364 489852 101370 489864
rect 122834 489852 122840 489864
rect 101364 489824 122840 489852
rect 101364 489812 101370 489824
rect 122834 489812 122840 489824
rect 122892 489812 122898 489864
rect 104250 489744 104256 489796
rect 104308 489784 104314 489796
rect 118694 489784 118700 489796
rect 104308 489756 118700 489784
rect 104308 489744 104314 489756
rect 118694 489744 118700 489756
rect 118752 489744 118758 489796
rect 110322 489676 110328 489728
rect 110380 489716 110386 489728
rect 113174 489716 113180 489728
rect 110380 489688 113180 489716
rect 110380 489676 110386 489688
rect 113174 489676 113180 489688
rect 113232 489676 113238 489728
rect 103330 488452 103336 488504
rect 103388 488492 103394 488504
rect 117314 488492 117320 488504
rect 103388 488464 117320 488492
rect 103388 488452 103394 488464
rect 117314 488452 117320 488464
rect 117372 488452 117378 488504
rect 103422 488384 103428 488436
rect 103480 488424 103486 488436
rect 109034 488424 109040 488436
rect 103480 488396 109040 488424
rect 103480 488384 103486 488396
rect 109034 488384 109040 488396
rect 109092 488384 109098 488436
rect 114462 488384 114468 488436
rect 114520 488424 114526 488436
rect 123018 488424 123024 488436
rect 114520 488396 123024 488424
rect 114520 488384 114526 488396
rect 123018 488384 123024 488396
rect 123076 488384 123082 488436
rect 53558 487840 53564 487892
rect 53616 487880 53622 487892
rect 59170 487880 59176 487892
rect 53616 487852 59176 487880
rect 53616 487840 53622 487852
rect 59170 487840 59176 487852
rect 59228 487840 59234 487892
rect 109034 487840 109040 487892
rect 109092 487880 109098 487892
rect 116118 487880 116124 487892
rect 109092 487852 116124 487880
rect 109092 487840 109098 487852
rect 116118 487840 116124 487852
rect 116176 487840 116182 487892
rect 117314 487840 117320 487892
rect 117372 487880 117378 487892
rect 125686 487880 125692 487892
rect 117372 487852 125692 487880
rect 117372 487840 117378 487852
rect 125686 487840 125692 487852
rect 125744 487840 125750 487892
rect 56502 487772 56508 487824
rect 56560 487812 56566 487824
rect 67634 487812 67640 487824
rect 56560 487784 67640 487812
rect 56560 487772 56566 487784
rect 67634 487772 67640 487784
rect 67692 487772 67698 487824
rect 103514 487772 103520 487824
rect 103572 487812 103578 487824
rect 134058 487812 134064 487824
rect 103572 487784 134064 487812
rect 103572 487772 103578 487784
rect 134058 487772 134064 487784
rect 134116 487812 134122 487824
rect 145006 487812 145012 487824
rect 134116 487784 145012 487812
rect 134116 487772 134122 487784
rect 145006 487772 145012 487784
rect 145064 487772 145070 487824
rect 59170 487160 59176 487212
rect 59228 487200 59234 487212
rect 67726 487200 67732 487212
rect 59228 487172 67732 487200
rect 59228 487160 59234 487172
rect 67726 487160 67732 487172
rect 67784 487160 67790 487212
rect 67634 485840 67640 485852
rect 35866 485812 67640 485840
rect 34238 485732 34244 485784
rect 34296 485772 34302 485784
rect 35158 485772 35164 485784
rect 34296 485744 35164 485772
rect 34296 485732 34302 485744
rect 35158 485732 35164 485744
rect 35216 485772 35222 485784
rect 35866 485772 35894 485812
rect 67634 485800 67640 485812
rect 67692 485800 67698 485852
rect 35216 485744 35894 485772
rect 35216 485732 35222 485744
rect 102318 485052 102324 485104
rect 102376 485092 102382 485104
rect 112162 485092 112168 485104
rect 102376 485064 112168 485092
rect 102376 485052 102382 485064
rect 112162 485052 112168 485064
rect 112220 485052 112226 485104
rect 65886 484576 65892 484628
rect 65944 484616 65950 484628
rect 68738 484616 68744 484628
rect 65944 484588 68744 484616
rect 65944 484576 65950 484588
rect 68738 484576 68744 484588
rect 68796 484576 68802 484628
rect 67634 484412 67640 484424
rect 57900 484384 67640 484412
rect 55030 484304 55036 484356
rect 55088 484344 55094 484356
rect 57330 484344 57336 484356
rect 55088 484316 57336 484344
rect 55088 484304 55094 484316
rect 57330 484304 57336 484316
rect 57388 484344 57394 484356
rect 57900 484344 57928 484384
rect 67634 484372 67640 484384
rect 67692 484372 67698 484424
rect 113082 484372 113088 484424
rect 113140 484412 113146 484424
rect 128446 484412 128452 484424
rect 113140 484384 128452 484412
rect 113140 484372 113146 484384
rect 128446 484372 128452 484384
rect 128504 484372 128510 484424
rect 57388 484316 57928 484344
rect 57388 484304 57394 484316
rect 102318 483624 102324 483676
rect 102376 483664 102382 483676
rect 125594 483664 125600 483676
rect 102376 483636 125600 483664
rect 102376 483624 102382 483636
rect 125594 483624 125600 483636
rect 125652 483664 125658 483676
rect 126238 483664 126244 483676
rect 125652 483636 126244 483664
rect 125652 483624 125658 483636
rect 126238 483624 126244 483636
rect 126296 483624 126302 483676
rect 67634 483052 67640 483064
rect 64846 483024 67640 483052
rect 35618 482944 35624 482996
rect 35676 482984 35682 482996
rect 64138 482984 64144 482996
rect 35676 482956 64144 482984
rect 35676 482944 35682 482956
rect 64138 482944 64144 482956
rect 64196 482984 64202 482996
rect 64846 482984 64874 483024
rect 67634 483012 67640 483024
rect 67692 483012 67698 483064
rect 146478 483052 146484 483064
rect 132466 483024 146484 483052
rect 64196 482956 64874 482984
rect 64196 482944 64202 482956
rect 102410 482944 102416 482996
rect 102468 482984 102474 482996
rect 131758 482984 131764 482996
rect 102468 482956 131764 482984
rect 102468 482944 102474 482956
rect 131758 482944 131764 482956
rect 131816 482984 131822 482996
rect 132466 482984 132494 483024
rect 146478 483012 146484 483024
rect 146536 483012 146542 483064
rect 131816 482956 132494 482984
rect 131816 482944 131822 482956
rect 43806 482876 43812 482928
rect 43864 482916 43870 482928
rect 68094 482916 68100 482928
rect 43864 482888 68100 482916
rect 43864 482876 43870 482888
rect 68094 482876 68100 482888
rect 68152 482876 68158 482928
rect 102318 482876 102324 482928
rect 102376 482916 102382 482928
rect 106366 482916 106372 482928
rect 102376 482888 106372 482916
rect 102376 482876 102382 482888
rect 106366 482876 106372 482888
rect 106424 482916 106430 482928
rect 107470 482916 107476 482928
rect 106424 482888 107476 482916
rect 106424 482876 106430 482888
rect 107470 482876 107476 482888
rect 107528 482876 107534 482928
rect 107470 482264 107476 482316
rect 107528 482304 107534 482316
rect 118786 482304 118792 482316
rect 107528 482276 118792 482304
rect 107528 482264 107534 482276
rect 118786 482264 118792 482276
rect 118844 482264 118850 482316
rect 102410 481584 102416 481636
rect 102468 481624 102474 481636
rect 113358 481624 113364 481636
rect 102468 481596 113364 481624
rect 102468 481584 102474 481596
rect 113358 481584 113364 481596
rect 113416 481624 113422 481636
rect 120166 481624 120172 481636
rect 113416 481596 120172 481624
rect 113416 481584 113422 481596
rect 120166 481584 120172 481596
rect 120224 481584 120230 481636
rect 102318 481516 102324 481568
rect 102376 481556 102382 481568
rect 110506 481556 110512 481568
rect 102376 481528 110512 481556
rect 102376 481516 102382 481528
rect 110506 481516 110512 481528
rect 110564 481556 110570 481568
rect 111702 481556 111708 481568
rect 110564 481528 111708 481556
rect 110564 481516 110570 481528
rect 111702 481516 111708 481528
rect 111760 481516 111766 481568
rect 111702 480904 111708 480956
rect 111760 480944 111766 480956
rect 118694 480944 118700 480956
rect 111760 480916 118700 480944
rect 111760 480904 111766 480916
rect 118694 480904 118700 480916
rect 118752 480904 118758 480956
rect 55030 480224 55036 480276
rect 55088 480264 55094 480276
rect 58618 480264 58624 480276
rect 55088 480236 58624 480264
rect 55088 480224 55094 480236
rect 58618 480224 58624 480236
rect 58676 480224 58682 480276
rect 68554 480264 68560 480276
rect 67606 480236 68560 480264
rect 39850 480156 39856 480208
rect 39908 480196 39914 480208
rect 67606 480196 67634 480236
rect 68554 480224 68560 480236
rect 68612 480224 68618 480276
rect 39908 480168 67634 480196
rect 39908 480156 39914 480168
rect 102318 480156 102324 480208
rect 102376 480196 102382 480208
rect 128354 480196 128360 480208
rect 102376 480168 128360 480196
rect 102376 480156 102382 480168
rect 128354 480156 128360 480168
rect 128412 480156 128418 480208
rect 58618 480088 58624 480140
rect 58676 480128 58682 480140
rect 67634 480128 67640 480140
rect 58676 480100 67640 480128
rect 58676 480088 58682 480100
rect 67634 480088 67640 480100
rect 67692 480088 67698 480140
rect 63218 480020 63224 480072
rect 63276 480060 63282 480072
rect 67726 480060 67732 480072
rect 63276 480032 67732 480060
rect 63276 480020 63282 480032
rect 67726 480020 67732 480032
rect 67784 480020 67790 480072
rect 128354 479476 128360 479528
rect 128412 479516 128418 479528
rect 151906 479516 151912 479528
rect 128412 479488 151912 479516
rect 128412 479476 128418 479488
rect 151906 479476 151912 479488
rect 151964 479476 151970 479528
rect 61746 478864 61752 478916
rect 61804 478904 61810 478916
rect 63218 478904 63224 478916
rect 61804 478876 63224 478904
rect 61804 478864 61810 478876
rect 63218 478864 63224 478876
rect 63276 478864 63282 478916
rect 111702 478252 111708 478304
rect 111760 478292 111766 478304
rect 116026 478292 116032 478304
rect 111760 478264 116032 478292
rect 111760 478252 111766 478264
rect 116026 478252 116032 478264
rect 116084 478252 116090 478304
rect 107470 477572 107476 477624
rect 107528 477612 107534 477624
rect 107838 477612 107844 477624
rect 107528 477584 107844 477612
rect 107528 477572 107534 477584
rect 107838 477572 107844 477584
rect 107896 477572 107902 477624
rect 102410 477504 102416 477556
rect 102468 477544 102474 477556
rect 116026 477544 116032 477556
rect 102468 477516 116032 477544
rect 102468 477504 102474 477516
rect 116026 477504 116032 477516
rect 116084 477504 116090 477556
rect 100662 477436 100668 477488
rect 100720 477476 100726 477488
rect 114646 477476 114652 477488
rect 100720 477448 114652 477476
rect 100720 477436 100726 477448
rect 114646 477436 114652 477448
rect 114704 477436 114710 477488
rect 108390 476144 108396 476196
rect 108448 476184 108454 476196
rect 109218 476184 109224 476196
rect 108448 476156 109224 476184
rect 108448 476144 108454 476156
rect 109218 476144 109224 476156
rect 109276 476144 109282 476196
rect 39666 476076 39672 476128
rect 39724 476116 39730 476128
rect 67634 476116 67640 476128
rect 39724 476088 67640 476116
rect 39724 476076 39730 476088
rect 67634 476076 67640 476088
rect 67692 476076 67698 476128
rect 102318 476076 102324 476128
rect 102376 476116 102382 476128
rect 116026 476116 116032 476128
rect 102376 476088 116032 476116
rect 102376 476076 102382 476088
rect 116026 476076 116032 476088
rect 116084 476116 116090 476128
rect 116084 476088 117912 476116
rect 116084 476076 116090 476088
rect 102410 476008 102416 476060
rect 102468 476048 102474 476060
rect 117406 476048 117412 476060
rect 102468 476020 117412 476048
rect 102468 476008 102474 476020
rect 117406 476008 117412 476020
rect 117464 476048 117470 476060
rect 117774 476048 117780 476060
rect 117464 476020 117780 476048
rect 117464 476008 117470 476020
rect 117774 476008 117780 476020
rect 117832 476008 117838 476060
rect 117884 476048 117912 476088
rect 120074 476048 120080 476060
rect 117884 476020 120080 476048
rect 120074 476008 120080 476020
rect 120132 476008 120138 476060
rect 102318 475940 102324 475992
rect 102376 475980 102382 475992
rect 115934 475980 115940 475992
rect 102376 475952 115940 475980
rect 102376 475940 102382 475952
rect 115934 475940 115940 475952
rect 115992 475940 115998 475992
rect 99742 475668 99748 475720
rect 99800 475708 99806 475720
rect 100754 475708 100760 475720
rect 99800 475680 100760 475708
rect 99800 475668 99806 475680
rect 100754 475668 100760 475680
rect 100812 475668 100818 475720
rect 53374 475328 53380 475380
rect 53432 475368 53438 475380
rect 53742 475368 53748 475380
rect 53432 475340 53748 475368
rect 53432 475328 53438 475340
rect 53742 475328 53748 475340
rect 53800 475368 53806 475380
rect 67634 475368 67640 475380
rect 53800 475340 67640 475368
rect 53800 475328 53806 475340
rect 67634 475328 67640 475340
rect 67692 475328 67698 475380
rect 117774 475328 117780 475380
rect 117832 475368 117838 475380
rect 132494 475368 132500 475380
rect 117832 475340 132500 475368
rect 117832 475328 117838 475340
rect 132494 475328 132500 475340
rect 132552 475328 132558 475380
rect 64690 474988 64696 475040
rect 64748 475028 64754 475040
rect 67634 475028 67640 475040
rect 64748 475000 67640 475028
rect 64748 474988 64754 475000
rect 67634 474988 67640 475000
rect 67692 474988 67698 475040
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 7558 474756 7564 474768
rect 3476 474728 7564 474756
rect 3476 474716 3482 474728
rect 7558 474716 7564 474728
rect 7616 474716 7622 474768
rect 107378 474716 107384 474768
rect 107436 474756 107442 474768
rect 107746 474756 107752 474768
rect 107436 474728 107752 474756
rect 107436 474716 107442 474728
rect 107746 474716 107752 474728
rect 107804 474716 107810 474768
rect 102318 474648 102324 474700
rect 102376 474688 102382 474700
rect 125870 474688 125876 474700
rect 102376 474660 125876 474688
rect 102376 474648 102382 474660
rect 125870 474648 125876 474660
rect 125928 474688 125934 474700
rect 128354 474688 128360 474700
rect 125928 474660 128360 474688
rect 125928 474648 125934 474660
rect 128354 474648 128360 474660
rect 128412 474648 128418 474700
rect 61838 474308 61844 474360
rect 61896 474348 61902 474360
rect 67634 474348 67640 474360
rect 61896 474320 67640 474348
rect 61896 474308 61902 474320
rect 67634 474308 67640 474320
rect 67692 474308 67698 474360
rect 102318 472744 102324 472796
rect 102376 472784 102382 472796
rect 131114 472784 131120 472796
rect 102376 472756 131120 472784
rect 102376 472744 102382 472756
rect 131114 472744 131120 472756
rect 131172 472744 131178 472796
rect 103422 472676 103428 472728
rect 103480 472716 103486 472728
rect 135162 472716 135168 472728
rect 103480 472688 135168 472716
rect 103480 472676 103486 472688
rect 135162 472676 135168 472688
rect 135220 472676 135226 472728
rect 102318 472608 102324 472660
rect 102376 472648 102382 472660
rect 136818 472648 136824 472660
rect 102376 472620 136824 472648
rect 102376 472608 102382 472620
rect 136818 472608 136824 472620
rect 136876 472648 136882 472660
rect 140866 472648 140872 472660
rect 136876 472620 140872 472648
rect 136876 472608 136882 472620
rect 140866 472608 140872 472620
rect 140924 472608 140930 472660
rect 105538 472200 105544 472252
rect 105596 472240 105602 472252
rect 110598 472240 110604 472252
rect 105596 472212 110604 472240
rect 105596 472200 105602 472212
rect 110598 472200 110604 472212
rect 110656 472200 110662 472252
rect 58986 471996 58992 472048
rect 59044 472036 59050 472048
rect 66162 472036 66168 472048
rect 59044 472008 66168 472036
rect 59044 471996 59050 472008
rect 66162 471996 66168 472008
rect 66220 472036 66226 472048
rect 67634 472036 67640 472048
rect 66220 472008 67640 472036
rect 66220 471996 66226 472008
rect 67634 471996 67640 472008
rect 67692 471996 67698 472048
rect 67450 471928 67456 471980
rect 67508 471968 67514 471980
rect 67726 471968 67732 471980
rect 67508 471940 67732 471968
rect 67508 471928 67514 471940
rect 67726 471928 67732 471940
rect 67784 471928 67790 471980
rect 102410 471928 102416 471980
rect 102468 471968 102474 471980
rect 107378 471968 107384 471980
rect 102468 471940 107384 471968
rect 102468 471928 102474 471940
rect 107378 471928 107384 471940
rect 107436 471928 107442 471980
rect 135162 471248 135168 471300
rect 135220 471288 135226 471300
rect 147766 471288 147772 471300
rect 135220 471260 147772 471288
rect 135220 471248 135226 471260
rect 147766 471248 147772 471260
rect 147824 471248 147830 471300
rect 107378 470976 107384 471028
rect 107436 471016 107442 471028
rect 108298 471016 108304 471028
rect 107436 470988 108304 471016
rect 107436 470976 107442 470988
rect 108298 470976 108304 470988
rect 108356 470976 108362 471028
rect 30282 470568 30288 470620
rect 30340 470608 30346 470620
rect 67634 470608 67640 470620
rect 30340 470580 38654 470608
rect 30340 470568 30346 470580
rect 38626 470540 38654 470580
rect 60706 470580 67640 470608
rect 39298 470540 39304 470552
rect 38626 470512 39304 470540
rect 39298 470500 39304 470512
rect 39356 470540 39362 470552
rect 60706 470540 60734 470580
rect 67634 470568 67640 470580
rect 67692 470568 67698 470620
rect 102778 470568 102784 470620
rect 102836 470608 102842 470620
rect 139486 470608 139492 470620
rect 102836 470580 139492 470608
rect 102836 470568 102842 470580
rect 139486 470568 139492 470580
rect 139544 470568 139550 470620
rect 147766 470568 147772 470620
rect 147824 470608 147830 470620
rect 580166 470608 580172 470620
rect 147824 470580 580172 470608
rect 147824 470568 147830 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 39356 470512 60734 470540
rect 39356 470500 39362 470512
rect 64782 470500 64788 470552
rect 64840 470540 64846 470552
rect 66898 470540 66904 470552
rect 64840 470512 66904 470540
rect 64840 470500 64846 470512
rect 66898 470500 66904 470512
rect 66956 470540 66962 470552
rect 67726 470540 67732 470552
rect 66956 470512 67732 470540
rect 66956 470500 66962 470512
rect 67726 470500 67732 470512
rect 67784 470500 67790 470552
rect 42518 469820 42524 469872
rect 42576 469860 42582 469872
rect 67174 469860 67180 469872
rect 42576 469832 67180 469860
rect 42576 469820 42582 469832
rect 67174 469820 67180 469832
rect 67232 469860 67238 469872
rect 67634 469860 67640 469872
rect 67232 469832 67640 469860
rect 67232 469820 67238 469832
rect 67634 469820 67640 469832
rect 67692 469820 67698 469872
rect 107010 469820 107016 469872
rect 107068 469860 107074 469872
rect 121638 469860 121644 469872
rect 107068 469832 121644 469860
rect 107068 469820 107074 469832
rect 121638 469820 121644 469832
rect 121696 469820 121702 469872
rect 102318 469140 102324 469192
rect 102376 469180 102382 469192
rect 120258 469180 120264 469192
rect 102376 469152 120264 469180
rect 102376 469140 102382 469152
rect 120258 469140 120264 469152
rect 120316 469140 120322 469192
rect 120258 468528 120264 468580
rect 120316 468568 120322 468580
rect 129918 468568 129924 468580
rect 120316 468540 129924 468568
rect 120316 468528 120322 468540
rect 129918 468528 129924 468540
rect 129976 468528 129982 468580
rect 103514 468460 103520 468512
rect 103572 468500 103578 468512
rect 138106 468500 138112 468512
rect 103572 468472 138112 468500
rect 103572 468460 103578 468472
rect 138106 468460 138112 468472
rect 138164 468500 138170 468512
rect 147674 468500 147680 468512
rect 138164 468472 147680 468500
rect 138164 468460 138170 468472
rect 147674 468460 147680 468472
rect 147732 468460 147738 468512
rect 64782 468120 64788 468172
rect 64840 468160 64846 468172
rect 66070 468160 66076 468172
rect 64840 468132 66076 468160
rect 64840 468120 64846 468132
rect 66070 468120 66076 468132
rect 66128 468160 66134 468172
rect 67634 468160 67640 468172
rect 66128 468132 67640 468160
rect 66128 468120 66134 468132
rect 67634 468120 67640 468132
rect 67692 468120 67698 468172
rect 119982 467780 119988 467832
rect 120040 467820 120046 467832
rect 123018 467820 123024 467832
rect 120040 467792 123024 467820
rect 120040 467780 120046 467792
rect 123018 467780 123024 467792
rect 123076 467780 123082 467832
rect 102778 466420 102784 466472
rect 102836 466460 102842 466472
rect 102836 466432 117268 466460
rect 102836 466420 102842 466432
rect 117240 466404 117268 466432
rect 102318 466352 102324 466404
rect 102376 466392 102382 466404
rect 111886 466392 111892 466404
rect 102376 466364 111892 466392
rect 102376 466352 102382 466364
rect 111886 466352 111892 466364
rect 111944 466392 111950 466404
rect 112346 466392 112352 466404
rect 111944 466364 112352 466392
rect 111944 466352 111950 466364
rect 112346 466352 112352 466364
rect 112404 466352 112410 466404
rect 117222 466392 117228 466404
rect 117135 466364 117228 466392
rect 117222 466352 117228 466364
rect 117280 466392 117286 466404
rect 128630 466392 128636 466404
rect 117280 466364 128636 466392
rect 117280 466352 117286 466364
rect 128630 466352 128636 466364
rect 128688 466352 128694 466404
rect 49602 465672 49608 465724
rect 49660 465712 49666 465724
rect 67634 465712 67640 465724
rect 49660 465684 67640 465712
rect 49660 465672 49666 465684
rect 67634 465672 67640 465684
rect 67692 465672 67698 465724
rect 112346 465672 112352 465724
rect 112404 465712 112410 465724
rect 119338 465712 119344 465724
rect 112404 465684 119344 465712
rect 112404 465672 112410 465684
rect 119338 465672 119344 465684
rect 119396 465672 119402 465724
rect 66162 465400 66168 465452
rect 66220 465440 66226 465452
rect 67634 465440 67640 465452
rect 66220 465412 67640 465440
rect 66220 465400 66226 465412
rect 67634 465400 67640 465412
rect 67692 465400 67698 465452
rect 142246 465100 142252 465112
rect 107580 465072 142252 465100
rect 48038 464992 48044 465044
rect 48096 465032 48102 465044
rect 49602 465032 49608 465044
rect 48096 465004 49608 465032
rect 48096 464992 48102 465004
rect 49602 464992 49608 465004
rect 49660 464992 49666 465044
rect 60458 464992 60464 465044
rect 60516 465032 60522 465044
rect 61930 465032 61936 465044
rect 60516 465004 61936 465032
rect 60516 464992 60522 465004
rect 61930 464992 61936 465004
rect 61988 465032 61994 465044
rect 67726 465032 67732 465044
rect 61988 465004 67732 465032
rect 61988 464992 61994 465004
rect 67726 464992 67732 465004
rect 67784 464992 67790 465044
rect 102318 464992 102324 465044
rect 102376 465032 102382 465044
rect 107470 465032 107476 465044
rect 102376 465004 107476 465032
rect 102376 464992 102382 465004
rect 107470 464992 107476 465004
rect 107528 465032 107534 465044
rect 107580 465032 107608 465072
rect 142246 465060 142252 465072
rect 142304 465060 142310 465112
rect 107528 465004 107608 465032
rect 107528 464992 107534 465004
rect 47854 464720 47860 464772
rect 47912 464760 47918 464772
rect 48130 464760 48136 464772
rect 47912 464732 48136 464760
rect 47912 464720 47918 464732
rect 48130 464720 48136 464732
rect 48188 464720 48194 464772
rect 47854 464312 47860 464364
rect 47912 464352 47918 464364
rect 67634 464352 67640 464364
rect 47912 464324 67640 464352
rect 47912 464312 47918 464324
rect 67634 464312 67640 464324
rect 67692 464312 67698 464364
rect 102410 463700 102416 463752
rect 102468 463740 102474 463752
rect 113082 463740 113088 463752
rect 102468 463712 113088 463740
rect 102468 463700 102474 463712
rect 113082 463700 113088 463712
rect 113140 463700 113146 463752
rect 136818 463740 136824 463752
rect 115860 463712 136824 463740
rect 51994 463632 52000 463684
rect 52052 463672 52058 463684
rect 52270 463672 52276 463684
rect 52052 463644 52276 463672
rect 52052 463632 52058 463644
rect 52270 463632 52276 463644
rect 52328 463632 52334 463684
rect 102318 463632 102324 463684
rect 102376 463672 102382 463684
rect 115198 463672 115204 463684
rect 102376 463644 115204 463672
rect 102376 463632 102382 463644
rect 115198 463632 115204 463644
rect 115256 463672 115262 463684
rect 115860 463672 115888 463712
rect 136818 463700 136824 463712
rect 136876 463700 136882 463752
rect 115256 463644 115888 463672
rect 115256 463632 115262 463644
rect 51994 462952 52000 463004
rect 52052 462992 52058 463004
rect 67634 462992 67640 463004
rect 52052 462964 67640 462992
rect 52052 462952 52058 462964
rect 67634 462952 67640 462964
rect 67692 462952 67698 463004
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 22738 462380 22744 462392
rect 3292 462352 22744 462380
rect 3292 462340 3298 462352
rect 22738 462340 22744 462352
rect 22796 462340 22802 462392
rect 133966 462380 133972 462392
rect 107580 462352 133972 462380
rect 102318 462272 102324 462324
rect 102376 462312 102382 462324
rect 107580 462312 107608 462352
rect 133966 462340 133972 462352
rect 134024 462340 134030 462392
rect 102376 462284 107608 462312
rect 102376 462272 102382 462284
rect 102318 460912 102324 460964
rect 102376 460952 102382 460964
rect 114646 460952 114652 460964
rect 102376 460924 114652 460952
rect 102376 460912 102382 460924
rect 114646 460912 114652 460924
rect 114704 460912 114710 460964
rect 50982 460232 50988 460284
rect 51040 460272 51046 460284
rect 67634 460272 67640 460284
rect 51040 460244 67640 460272
rect 51040 460232 51046 460244
rect 67634 460232 67640 460244
rect 67692 460232 67698 460284
rect 115474 460232 115480 460284
rect 115532 460272 115538 460284
rect 116210 460272 116216 460284
rect 115532 460244 116216 460272
rect 115532 460232 115538 460244
rect 116210 460232 116216 460244
rect 116268 460272 116274 460284
rect 126974 460272 126980 460284
rect 116268 460244 126980 460272
rect 116268 460232 116274 460244
rect 126974 460232 126980 460244
rect 127032 460232 127038 460284
rect 44450 460164 44456 460216
rect 44508 460204 44514 460216
rect 45462 460204 45468 460216
rect 44508 460176 45468 460204
rect 44508 460164 44514 460176
rect 45462 460164 45468 460176
rect 45520 460204 45526 460216
rect 67726 460204 67732 460216
rect 45520 460176 67732 460204
rect 45520 460164 45526 460176
rect 67726 460164 67732 460176
rect 67784 460164 67790 460216
rect 102318 460164 102324 460216
rect 102376 460204 102382 460216
rect 102376 460176 103514 460204
rect 102376 460164 102382 460176
rect 103486 460136 103514 460176
rect 106182 460136 106188 460148
rect 103486 460108 106188 460136
rect 106182 460096 106188 460108
rect 106240 460136 106246 460148
rect 115290 460136 115296 460148
rect 106240 460108 115296 460136
rect 106240 460096 106246 460108
rect 115290 460096 115296 460108
rect 115348 460096 115354 460148
rect 50798 459620 50804 459672
rect 50856 459660 50862 459672
rect 50982 459660 50988 459672
rect 50856 459632 50988 459660
rect 50856 459620 50862 459632
rect 50982 459620 50988 459632
rect 51040 459620 51046 459672
rect 45462 459552 45468 459604
rect 45520 459592 45526 459604
rect 62758 459592 62764 459604
rect 45520 459564 62764 459592
rect 45520 459552 45526 459564
rect 62758 459552 62764 459564
rect 62816 459552 62822 459604
rect 102870 459552 102876 459604
rect 102928 459592 102934 459604
rect 102928 459564 106228 459592
rect 102928 459552 102934 459564
rect 62776 459524 62804 459552
rect 106200 459536 106228 459564
rect 67634 459524 67640 459536
rect 62776 459496 67640 459524
rect 67634 459484 67640 459496
rect 67692 459484 67698 459536
rect 106182 459524 106188 459536
rect 106095 459496 106188 459524
rect 106182 459484 106188 459496
rect 106240 459524 106246 459536
rect 136634 459524 136640 459536
rect 106240 459496 136640 459524
rect 106240 459484 106246 459496
rect 136634 459484 136640 459496
rect 136692 459484 136698 459536
rect 102318 459416 102324 459468
rect 102376 459456 102382 459468
rect 115474 459456 115480 459468
rect 102376 459428 115480 459456
rect 102376 459416 102382 459428
rect 115474 459416 115480 459428
rect 115532 459416 115538 459468
rect 107746 458872 107752 458924
rect 107804 458912 107810 458924
rect 142338 458912 142344 458924
rect 107804 458884 142344 458912
rect 107804 458872 107810 458884
rect 142338 458872 142344 458884
rect 142396 458912 142402 458924
rect 146386 458912 146392 458924
rect 142396 458884 146392 458912
rect 142396 458872 142402 458884
rect 146386 458872 146392 458884
rect 146444 458872 146450 458924
rect 34146 458804 34152 458856
rect 34204 458844 34210 458856
rect 67266 458844 67272 458856
rect 34204 458816 67272 458844
rect 34204 458804 34210 458816
rect 67266 458804 67272 458816
rect 67324 458804 67330 458856
rect 103514 458804 103520 458856
rect 103572 458844 103578 458856
rect 140958 458844 140964 458856
rect 103572 458816 140964 458844
rect 103572 458804 103578 458816
rect 140958 458804 140964 458816
rect 141016 458844 141022 458856
rect 149146 458844 149152 458856
rect 141016 458816 149152 458844
rect 141016 458804 141022 458816
rect 149146 458804 149152 458816
rect 149204 458804 149210 458856
rect 36906 458192 36912 458244
rect 36964 458232 36970 458244
rect 44450 458232 44456 458244
rect 36964 458204 44456 458232
rect 36964 458192 36970 458204
rect 44450 458192 44456 458204
rect 44508 458192 44514 458244
rect 102410 458192 102416 458244
rect 102468 458232 102474 458244
rect 115198 458232 115204 458244
rect 102468 458204 115204 458232
rect 102468 458192 102474 458204
rect 115198 458192 115204 458204
rect 115256 458192 115262 458244
rect 53650 458124 53656 458176
rect 53708 458164 53714 458176
rect 68094 458164 68100 458176
rect 53708 458136 68100 458164
rect 53708 458124 53714 458136
rect 68094 458124 68100 458136
rect 68152 458124 68158 458176
rect 108482 458124 108488 458176
rect 108540 458164 108546 458176
rect 114830 458164 114836 458176
rect 108540 458136 114836 458164
rect 108540 458124 108546 458136
rect 114830 458124 114836 458136
rect 114888 458124 114894 458176
rect 43898 457444 43904 457496
rect 43956 457484 43962 457496
rect 67634 457484 67640 457496
rect 43956 457456 67640 457484
rect 43956 457444 43962 457456
rect 67634 457444 67640 457456
rect 67692 457444 67698 457496
rect 103514 457104 103520 457156
rect 103572 457144 103578 457156
rect 107746 457144 107752 457156
rect 103572 457116 107752 457144
rect 103572 457104 103578 457116
rect 107746 457104 107752 457116
rect 107804 457104 107810 457156
rect 102226 455472 102232 455524
rect 102284 455512 102290 455524
rect 105538 455512 105544 455524
rect 102284 455484 105544 455512
rect 102284 455472 102290 455484
rect 105538 455472 105544 455484
rect 105596 455472 105602 455524
rect 67634 455444 67640 455456
rect 40696 455416 67640 455444
rect 40696 455388 40724 455416
rect 67634 455404 67640 455416
rect 67692 455404 67698 455456
rect 102410 455404 102416 455456
rect 102468 455444 102474 455456
rect 102468 455416 132494 455444
rect 102468 455404 102474 455416
rect 35710 455336 35716 455388
rect 35768 455376 35774 455388
rect 40678 455376 40684 455388
rect 35768 455348 40684 455376
rect 35768 455336 35774 455348
rect 40678 455336 40684 455348
rect 40736 455336 40742 455388
rect 102226 455336 102232 455388
rect 102284 455376 102290 455388
rect 107562 455376 107568 455388
rect 102284 455348 107568 455376
rect 102284 455336 102290 455348
rect 107562 455336 107568 455348
rect 107620 455336 107626 455388
rect 132466 455376 132494 455416
rect 133782 455376 133788 455388
rect 132466 455348 133788 455376
rect 133782 455336 133788 455348
rect 133840 455376 133846 455388
rect 139394 455376 139400 455388
rect 133840 455348 139400 455376
rect 133840 455336 133846 455348
rect 139394 455336 139400 455348
rect 139452 455336 139458 455388
rect 49602 454656 49608 454708
rect 49660 454696 49666 454708
rect 54938 454696 54944 454708
rect 49660 454668 54944 454696
rect 49660 454656 49666 454668
rect 54938 454656 54944 454668
rect 54996 454696 55002 454708
rect 67726 454696 67732 454708
rect 54996 454668 67732 454696
rect 54996 454656 55002 454668
rect 67726 454656 67732 454668
rect 67784 454656 67790 454708
rect 48222 454044 48228 454096
rect 48280 454084 48286 454096
rect 55122 454084 55128 454096
rect 48280 454056 55128 454084
rect 48280 454044 48286 454056
rect 55122 454044 55128 454056
rect 55180 454084 55186 454096
rect 67634 454084 67640 454096
rect 55180 454056 67640 454084
rect 55180 454044 55186 454056
rect 67634 454044 67640 454056
rect 67692 454044 67698 454096
rect 102226 453976 102232 454028
rect 102284 454016 102290 454028
rect 124398 454016 124404 454028
rect 102284 453988 124404 454016
rect 102284 453976 102290 453988
rect 124398 453976 124404 453988
rect 124456 454016 124462 454028
rect 129826 454016 129832 454028
rect 124456 453988 129832 454016
rect 124456 453976 124462 453988
rect 129826 453976 129832 453988
rect 129884 453976 129890 454028
rect 102226 453364 102232 453416
rect 102284 453404 102290 453416
rect 106090 453404 106096 453416
rect 102284 453376 106096 453404
rect 102284 453364 102290 453376
rect 106090 453364 106096 453376
rect 106148 453364 106154 453416
rect 50890 453296 50896 453348
rect 50948 453336 50954 453348
rect 67634 453336 67640 453348
rect 50948 453308 67640 453336
rect 50948 453296 50954 453308
rect 67634 453296 67640 453308
rect 67692 453296 67698 453348
rect 34238 452616 34244 452668
rect 34296 452656 34302 452668
rect 67726 452656 67732 452668
rect 34296 452628 67732 452656
rect 34296 452616 34302 452628
rect 67726 452616 67732 452628
rect 67784 452656 67790 452668
rect 68278 452656 68284 452668
rect 67784 452628 68284 452656
rect 67784 452616 67790 452628
rect 68278 452616 68284 452628
rect 68336 452616 68342 452668
rect 102226 452548 102232 452600
rect 102284 452588 102290 452600
rect 136726 452588 136732 452600
rect 102284 452560 136732 452588
rect 102284 452548 102290 452560
rect 136726 452548 136732 452560
rect 136784 452588 136790 452600
rect 137094 452588 137100 452600
rect 136784 452560 137100 452588
rect 136784 452548 136790 452560
rect 137094 452548 137100 452560
rect 137152 452548 137158 452600
rect 42702 451868 42708 451920
rect 42760 451908 42766 451920
rect 66990 451908 66996 451920
rect 42760 451880 66996 451908
rect 42760 451868 42766 451880
rect 66990 451868 66996 451880
rect 67048 451868 67054 451920
rect 103514 451868 103520 451920
rect 103572 451908 103578 451920
rect 142154 451908 142160 451920
rect 103572 451880 142160 451908
rect 103572 451868 103578 451880
rect 142154 451868 142160 451880
rect 142212 451908 142218 451920
rect 150526 451908 150532 451920
rect 142212 451880 150532 451908
rect 142212 451868 142218 451880
rect 150526 451868 150532 451880
rect 150584 451868 150590 451920
rect 137094 451256 137100 451308
rect 137152 451296 137158 451308
rect 142338 451296 142344 451308
rect 137152 451268 142344 451296
rect 137152 451256 137158 451268
rect 142338 451256 142344 451268
rect 142396 451256 142402 451308
rect 100846 450576 100852 450628
rect 100904 450616 100910 450628
rect 105814 450616 105820 450628
rect 100904 450588 105820 450616
rect 100904 450576 100910 450588
rect 105814 450576 105820 450588
rect 105872 450616 105878 450628
rect 120074 450616 120080 450628
rect 105872 450588 120080 450616
rect 105872 450576 105878 450588
rect 120074 450576 120080 450588
rect 120132 450576 120138 450628
rect 107562 450508 107568 450560
rect 107620 450548 107626 450560
rect 140774 450548 140780 450560
rect 107620 450520 140780 450548
rect 107620 450508 107626 450520
rect 140774 450508 140780 450520
rect 140832 450508 140838 450560
rect 62758 449936 62764 449948
rect 62132 449908 62764 449936
rect 44082 449828 44088 449880
rect 44140 449868 44146 449880
rect 62132 449868 62160 449908
rect 62758 449896 62764 449908
rect 62816 449936 62822 449948
rect 67634 449936 67640 449948
rect 62816 449908 67640 449936
rect 62816 449896 62822 449908
rect 67634 449896 67640 449908
rect 67692 449896 67698 449948
rect 140774 449896 140780 449948
rect 140832 449936 140838 449948
rect 143626 449936 143632 449948
rect 140832 449908 143632 449936
rect 140832 449896 140838 449908
rect 143626 449896 143632 449908
rect 143684 449896 143690 449948
rect 44140 449840 62160 449868
rect 44140 449828 44146 449840
rect 102410 449828 102416 449880
rect 102468 449868 102474 449880
rect 107562 449868 107568 449880
rect 102468 449840 107568 449868
rect 102468 449828 102474 449840
rect 107562 449828 107568 449840
rect 107620 449828 107626 449880
rect 63402 449216 63408 449268
rect 63460 449256 63466 449268
rect 67726 449256 67732 449268
rect 63460 449228 67732 449256
rect 63460 449216 63466 449228
rect 67726 449216 67732 449228
rect 67784 449216 67790 449268
rect 102134 449216 102140 449268
rect 102192 449256 102198 449268
rect 107470 449256 107476 449268
rect 102192 449228 107476 449256
rect 102192 449216 102198 449228
rect 107470 449216 107476 449228
rect 107528 449216 107534 449268
rect 41138 449148 41144 449200
rect 41196 449188 41202 449200
rect 67634 449188 67640 449200
rect 41196 449160 67640 449188
rect 41196 449148 41202 449160
rect 67634 449148 67640 449160
rect 67692 449148 67698 449200
rect 106182 449148 106188 449200
rect 106240 449188 106246 449200
rect 134150 449188 134156 449200
rect 106240 449160 134156 449188
rect 106240 449148 106246 449160
rect 134150 449148 134156 449160
rect 134208 449188 134214 449200
rect 140774 449188 140780 449200
rect 134208 449160 140780 449188
rect 134208 449148 134214 449160
rect 140774 449148 140780 449160
rect 140832 449148 140838 449200
rect 107378 448604 107384 448656
rect 107436 448644 107442 448656
rect 107436 448616 113174 448644
rect 107436 448604 107442 448616
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 46198 448576 46204 448588
rect 3200 448548 46204 448576
rect 3200 448536 3206 448548
rect 46198 448536 46204 448548
rect 46256 448536 46262 448588
rect 106918 448536 106924 448588
rect 106976 448576 106982 448588
rect 107470 448576 107476 448588
rect 106976 448548 107476 448576
rect 106976 448536 106982 448548
rect 107470 448536 107476 448548
rect 107528 448536 107534 448588
rect 113146 448576 113174 448616
rect 144914 448576 144920 448588
rect 113146 448548 144920 448576
rect 144914 448536 144920 448548
rect 144972 448536 144978 448588
rect 61930 448468 61936 448520
rect 61988 448508 61994 448520
rect 63310 448508 63316 448520
rect 61988 448480 63316 448508
rect 61988 448468 61994 448480
rect 63310 448468 63316 448480
rect 63368 448508 63374 448520
rect 67634 448508 67640 448520
rect 63368 448480 67640 448508
rect 63368 448468 63374 448480
rect 67634 448468 67640 448480
rect 67692 448468 67698 448520
rect 102134 448468 102140 448520
rect 102192 448508 102198 448520
rect 106182 448508 106188 448520
rect 102192 448480 106188 448508
rect 102192 448468 102198 448480
rect 106182 448468 106188 448480
rect 106240 448468 106246 448520
rect 102410 448400 102416 448452
rect 102468 448440 102474 448452
rect 107378 448440 107384 448452
rect 102468 448412 107384 448440
rect 102468 448400 102474 448412
rect 107378 448400 107384 448412
rect 107436 448400 107442 448452
rect 41138 447924 41144 447976
rect 41196 447964 41202 447976
rect 42058 447964 42064 447976
rect 41196 447936 42064 447964
rect 41196 447924 41202 447936
rect 42058 447924 42064 447936
rect 42116 447924 42122 447976
rect 100018 447856 100024 447908
rect 100076 447896 100082 447908
rect 112070 447896 112076 447908
rect 100076 447868 112076 447896
rect 100076 447856 100082 447868
rect 112070 447856 112076 447868
rect 112128 447856 112134 447908
rect 105722 447788 105728 447840
rect 105780 447828 105786 447840
rect 118878 447828 118884 447840
rect 105780 447800 118884 447828
rect 105780 447788 105786 447800
rect 118878 447788 118884 447800
rect 118936 447788 118942 447840
rect 60642 445884 60648 445936
rect 60700 445924 60706 445936
rect 64506 445924 64512 445936
rect 60700 445896 64512 445924
rect 60700 445884 60706 445896
rect 64506 445884 64512 445896
rect 64564 445924 64570 445936
rect 67634 445924 67640 445936
rect 64564 445896 67640 445924
rect 64564 445884 64570 445896
rect 67634 445884 67640 445896
rect 67692 445884 67698 445936
rect 102134 445816 102140 445868
rect 102192 445856 102198 445868
rect 105538 445856 105544 445868
rect 102192 445828 105544 445856
rect 102192 445816 102198 445828
rect 105538 445816 105544 445828
rect 105596 445816 105602 445868
rect 65518 445788 65524 445800
rect 64846 445760 65524 445788
rect 37182 445680 37188 445732
rect 37240 445720 37246 445732
rect 64846 445720 64874 445760
rect 65518 445748 65524 445760
rect 65576 445788 65582 445800
rect 67726 445788 67732 445800
rect 65576 445760 67732 445788
rect 65576 445748 65582 445760
rect 67726 445748 67732 445760
rect 67784 445748 67790 445800
rect 37240 445692 64874 445720
rect 37240 445680 37246 445692
rect 133138 445176 133144 445188
rect 122806 445148 133144 445176
rect 103514 445068 103520 445120
rect 103572 445108 103578 445120
rect 122806 445108 122834 445148
rect 133138 445136 133144 445148
rect 133196 445176 133202 445188
rect 134058 445176 134064 445188
rect 133196 445148 134064 445176
rect 133196 445136 133202 445148
rect 134058 445136 134064 445148
rect 134116 445136 134122 445188
rect 103572 445080 122834 445108
rect 103572 445068 103578 445080
rect 38562 445000 38568 445052
rect 38620 445040 38626 445052
rect 67634 445040 67640 445052
rect 38620 445012 67640 445040
rect 38620 445000 38626 445012
rect 67634 445000 67640 445012
rect 67692 445000 67698 445052
rect 102594 445000 102600 445052
rect 102652 445040 102658 445052
rect 132586 445040 132592 445052
rect 102652 445012 132592 445040
rect 102652 445000 102658 445012
rect 132586 445000 132592 445012
rect 132644 445040 132650 445052
rect 136726 445040 136732 445052
rect 132644 445012 136732 445040
rect 132644 445000 132650 445012
rect 136726 445000 136732 445012
rect 136784 445000 136790 445052
rect 49418 444320 49424 444372
rect 49476 444360 49482 444372
rect 67634 444360 67640 444372
rect 49476 444332 67640 444360
rect 49476 444320 49482 444332
rect 67634 444320 67640 444332
rect 67692 444320 67698 444372
rect 45186 443640 45192 443692
rect 45244 443680 45250 443692
rect 49418 443680 49424 443692
rect 45244 443652 49424 443680
rect 45244 443640 45250 443652
rect 49418 443640 49424 443652
rect 49476 443640 49482 443692
rect 106090 443640 106096 443692
rect 106148 443680 106154 443692
rect 117406 443680 117412 443692
rect 106148 443652 117412 443680
rect 106148 443640 106154 443652
rect 117406 443640 117412 443652
rect 117464 443640 117470 443692
rect 34330 443028 34336 443080
rect 34388 443068 34394 443080
rect 36998 443068 37004 443080
rect 34388 443040 37004 443068
rect 34388 443028 34394 443040
rect 36998 443028 37004 443040
rect 37056 443068 37062 443080
rect 37056 443040 45554 443068
rect 37056 443028 37062 443040
rect 35710 442960 35716 443012
rect 35768 443000 35774 443012
rect 38562 443000 38568 443012
rect 35768 442972 38568 443000
rect 35768 442960 35774 442972
rect 38562 442960 38568 442972
rect 38620 442960 38626 443012
rect 45526 443000 45554 443040
rect 67726 443000 67732 443012
rect 45526 442972 67732 443000
rect 67726 442960 67732 442972
rect 67784 442960 67790 443012
rect 39758 442892 39764 442944
rect 39816 442932 39822 442944
rect 67634 442932 67640 442944
rect 39816 442904 67640 442932
rect 39816 442892 39822 442904
rect 67634 442892 67640 442904
rect 67692 442892 67698 442944
rect 102870 442824 102876 442876
rect 102928 442864 102934 442876
rect 127158 442864 127164 442876
rect 102928 442836 127164 442864
rect 102928 442824 102934 442836
rect 127158 442824 127164 442836
rect 127216 442864 127222 442876
rect 127434 442864 127440 442876
rect 127216 442836 127440 442864
rect 127216 442824 127222 442836
rect 127434 442824 127440 442836
rect 127492 442824 127498 442876
rect 38562 442280 38568 442332
rect 38620 442320 38626 442332
rect 39758 442320 39764 442332
rect 38620 442292 39764 442320
rect 38620 442280 38626 442292
rect 39758 442280 39764 442292
rect 39816 442280 39822 442332
rect 127434 442212 127440 442264
rect 127492 442252 127498 442264
rect 143810 442252 143816 442264
rect 127492 442224 143816 442252
rect 127492 442212 127498 442224
rect 143810 442212 143816 442224
rect 143868 442212 143874 442264
rect 103330 441600 103336 441652
rect 103388 441640 103394 441652
rect 139578 441640 139584 441652
rect 103388 441612 139584 441640
rect 103388 441600 103394 441612
rect 139578 441600 139584 441612
rect 139636 441600 139642 441652
rect 45370 440852 45376 440904
rect 45428 440892 45434 440904
rect 117590 440892 117596 440904
rect 45428 440864 64874 440892
rect 45428 440852 45434 440864
rect 64846 440756 64874 440864
rect 93826 440864 117596 440892
rect 64846 440728 72372 440756
rect 72344 440700 72372 440728
rect 69842 440648 69848 440700
rect 69900 440688 69906 440700
rect 70394 440688 70400 440700
rect 69900 440660 70400 440688
rect 69900 440648 69906 440660
rect 70394 440648 70400 440660
rect 70452 440648 70458 440700
rect 72326 440648 72332 440700
rect 72384 440648 72390 440700
rect 87690 440648 87696 440700
rect 87748 440688 87754 440700
rect 88426 440688 88432 440700
rect 87748 440660 88432 440688
rect 87748 440648 87754 440660
rect 88426 440648 88432 440660
rect 88484 440688 88490 440700
rect 93826 440688 93854 440864
rect 117590 440852 117596 440864
rect 117648 440852 117654 440904
rect 88484 440660 93854 440688
rect 88484 440648 88490 440660
rect 62022 440308 62028 440360
rect 62080 440348 62086 440360
rect 67542 440348 67548 440360
rect 62080 440320 67548 440348
rect 62080 440308 62086 440320
rect 67542 440308 67548 440320
rect 67600 440348 67606 440360
rect 67726 440348 67732 440360
rect 67600 440320 67732 440348
rect 67600 440308 67606 440320
rect 67726 440308 67732 440320
rect 67784 440308 67790 440360
rect 65978 440240 65984 440292
rect 66036 440280 66042 440292
rect 71130 440280 71136 440292
rect 66036 440252 71136 440280
rect 66036 440240 66042 440252
rect 71130 440240 71136 440252
rect 71188 440240 71194 440292
rect 102870 440240 102876 440292
rect 102928 440280 102934 440292
rect 138106 440280 138112 440292
rect 102928 440252 138112 440280
rect 102928 440240 102934 440252
rect 138106 440240 138112 440252
rect 138164 440240 138170 440292
rect 97442 440172 97448 440224
rect 97500 440212 97506 440224
rect 98638 440212 98644 440224
rect 97500 440184 98644 440212
rect 97500 440172 97506 440184
rect 98638 440172 98644 440184
rect 98696 440212 98702 440224
rect 105722 440212 105728 440224
rect 98696 440184 105728 440212
rect 98696 440172 98702 440184
rect 105722 440172 105728 440184
rect 105780 440172 105786 440224
rect 57606 439492 57612 439544
rect 57664 439532 57670 439544
rect 76006 439532 76012 439544
rect 57664 439504 76012 439532
rect 57664 439492 57670 439504
rect 76006 439492 76012 439504
rect 76064 439532 76070 439544
rect 77754 439532 77760 439544
rect 76064 439504 77760 439532
rect 76064 439492 76070 439504
rect 77754 439492 77760 439504
rect 77812 439492 77818 439544
rect 56226 439356 56232 439408
rect 56284 439396 56290 439408
rect 57238 439396 57244 439408
rect 56284 439368 57244 439396
rect 56284 439356 56290 439368
rect 57238 439356 57244 439368
rect 57296 439356 57302 439408
rect 121914 439288 121920 439340
rect 121972 439328 121978 439340
rect 122926 439328 122932 439340
rect 121972 439300 122932 439328
rect 121972 439288 121978 439300
rect 122926 439288 122932 439300
rect 122984 439288 122990 439340
rect 7558 439152 7564 439204
rect 7616 439192 7622 439204
rect 96430 439192 96436 439204
rect 7616 439164 96436 439192
rect 7616 439152 7622 439164
rect 96430 439152 96436 439164
rect 96488 439152 96494 439204
rect 57238 439084 57244 439136
rect 57296 439124 57302 439136
rect 80606 439124 80612 439136
rect 57296 439096 80612 439124
rect 57296 439084 57302 439096
rect 80606 439084 80612 439096
rect 80664 439084 80670 439136
rect 103054 439084 103060 439136
rect 103112 439124 103118 439136
rect 136910 439124 136916 439136
rect 103112 439096 136916 439124
rect 103112 439084 103118 439096
rect 136910 439084 136916 439096
rect 136968 439084 136974 439136
rect 56410 439016 56416 439068
rect 56468 439056 56474 439068
rect 74626 439056 74632 439068
rect 56468 439028 74632 439056
rect 56468 439016 56474 439028
rect 74626 439016 74632 439028
rect 74684 439056 74690 439068
rect 75822 439056 75828 439068
rect 74684 439028 75828 439056
rect 74684 439016 74690 439028
rect 75822 439016 75828 439028
rect 75880 439016 75886 439068
rect 97718 439016 97724 439068
rect 97776 439056 97782 439068
rect 108390 439056 108396 439068
rect 97776 439028 108396 439056
rect 97776 439016 97782 439028
rect 108390 439016 108396 439028
rect 108448 439016 108454 439068
rect 41322 438948 41328 439000
rect 41380 438988 41386 439000
rect 73890 438988 73896 439000
rect 41380 438960 73896 438988
rect 41380 438948 41386 438960
rect 73890 438948 73896 438960
rect 73948 438948 73954 439000
rect 88702 438948 88708 439000
rect 88760 438988 88766 439000
rect 121546 438988 121552 439000
rect 88760 438960 121552 438988
rect 88760 438948 88766 438960
rect 121546 438948 121552 438960
rect 121604 438948 121610 439000
rect 72970 438880 72976 438932
rect 73028 438920 73034 438932
rect 73430 438920 73436 438932
rect 73028 438892 73436 438920
rect 73028 438880 73034 438892
rect 73430 438880 73436 438892
rect 73488 438880 73494 438932
rect 93854 438880 93860 438932
rect 93912 438920 93918 438932
rect 95142 438920 95148 438932
rect 93912 438892 95148 438920
rect 93912 438880 93918 438892
rect 95142 438880 95148 438892
rect 95200 438920 95206 438932
rect 95200 438892 96568 438920
rect 95200 438880 95206 438892
rect 22738 438812 22744 438864
rect 22796 438852 22802 438864
rect 50706 438852 50712 438864
rect 22796 438824 50712 438852
rect 22796 438812 22802 438824
rect 50706 438812 50712 438824
rect 50764 438812 50770 438864
rect 96540 438852 96568 438892
rect 96614 438880 96620 438932
rect 96672 438920 96678 438932
rect 97718 438920 97724 438932
rect 96672 438892 97724 438920
rect 96672 438880 96678 438892
rect 97718 438880 97724 438892
rect 97776 438880 97782 438932
rect 108482 438920 108488 438932
rect 97828 438892 108488 438920
rect 97828 438852 97856 438892
rect 108482 438880 108488 438892
rect 108540 438880 108546 438932
rect 96540 438824 97856 438852
rect 99650 438812 99656 438864
rect 99708 438852 99714 438864
rect 121914 438852 121920 438864
rect 99708 438824 121920 438852
rect 99708 438812 99714 438824
rect 121914 438812 121920 438824
rect 121972 438852 121978 438864
rect 122190 438852 122196 438864
rect 121972 438824 122196 438852
rect 121972 438812 121978 438824
rect 122190 438812 122196 438824
rect 122248 438812 122254 438864
rect 45278 438744 45284 438796
rect 45336 438784 45342 438796
rect 78398 438784 78404 438796
rect 45336 438756 78404 438784
rect 45336 438744 45342 438756
rect 78398 438744 78404 438756
rect 78456 438744 78462 438796
rect 99006 438744 99012 438796
rect 99064 438784 99070 438796
rect 128538 438784 128544 438796
rect 99064 438756 128544 438784
rect 99064 438744 99070 438756
rect 128538 438744 128544 438756
rect 128596 438744 128602 438796
rect 46566 438676 46572 438728
rect 46624 438716 46630 438728
rect 77110 438716 77116 438728
rect 46624 438688 77116 438716
rect 46624 438676 46630 438688
rect 77110 438676 77116 438688
rect 77168 438676 77174 438728
rect 96430 438676 96436 438728
rect 96488 438716 96494 438728
rect 121730 438716 121736 438728
rect 96488 438688 121736 438716
rect 96488 438676 96494 438688
rect 121730 438676 121736 438688
rect 121788 438676 121794 438728
rect 59078 438608 59084 438660
rect 59136 438648 59142 438660
rect 70026 438648 70032 438660
rect 59136 438620 70032 438648
rect 59136 438608 59142 438620
rect 70026 438608 70032 438620
rect 70084 438608 70090 438660
rect 93210 438608 93216 438660
rect 93268 438648 93274 438660
rect 93762 438648 93768 438660
rect 93268 438620 93768 438648
rect 93268 438608 93274 438620
rect 93762 438608 93768 438620
rect 93820 438648 93826 438660
rect 107010 438648 107016 438660
rect 93820 438620 107016 438648
rect 93820 438608 93826 438620
rect 107010 438608 107016 438620
rect 107068 438608 107074 438660
rect 46198 438540 46204 438592
rect 46256 438580 46262 438592
rect 99742 438580 99748 438592
rect 46256 438552 99748 438580
rect 46256 438540 46262 438552
rect 99742 438540 99748 438552
rect 99800 438540 99806 438592
rect 93670 438472 93676 438524
rect 93728 438512 93734 438524
rect 102318 438512 102324 438524
rect 93728 438484 102324 438512
rect 93728 438472 93734 438484
rect 102318 438472 102324 438484
rect 102376 438472 102382 438524
rect 69382 438336 69388 438388
rect 69440 438376 69446 438388
rect 71866 438376 71872 438388
rect 69440 438348 71872 438376
rect 69440 438336 69446 438348
rect 71866 438336 71872 438348
rect 71924 438336 71930 438388
rect 98362 438268 98368 438320
rect 98420 438308 98426 438320
rect 99282 438308 99288 438320
rect 98420 438280 99288 438308
rect 98420 438268 98426 438280
rect 99282 438268 99288 438280
rect 99340 438308 99346 438320
rect 102226 438308 102232 438320
rect 99340 438280 102232 438308
rect 99340 438268 99346 438280
rect 102226 438268 102232 438280
rect 102284 438268 102290 438320
rect 65886 438200 65892 438252
rect 65944 438240 65950 438252
rect 75178 438240 75184 438252
rect 65944 438212 75184 438240
rect 65944 438200 65950 438212
rect 75178 438200 75184 438212
rect 75236 438200 75242 438252
rect 50706 438132 50712 438184
rect 50764 438172 50770 438184
rect 52178 438172 52184 438184
rect 50764 438144 52184 438172
rect 50764 438132 50770 438144
rect 52178 438132 52184 438144
rect 52236 438172 52242 438184
rect 83550 438172 83556 438184
rect 52236 438144 83556 438172
rect 52236 438132 52242 438144
rect 83550 438132 83556 438144
rect 83608 438132 83614 438184
rect 69290 437860 69296 437912
rect 69348 437900 69354 437912
rect 70026 437900 70032 437912
rect 69348 437872 70032 437900
rect 69348 437860 69354 437872
rect 70026 437860 70032 437872
rect 70084 437860 70090 437912
rect 91094 437588 91100 437640
rect 91152 437628 91158 437640
rect 92566 437628 92572 437640
rect 91152 437600 92572 437628
rect 91152 437588 91158 437600
rect 92566 437588 92572 437600
rect 92624 437588 92630 437640
rect 78398 437520 78404 437572
rect 78456 437560 78462 437572
rect 80698 437560 80704 437572
rect 78456 437532 80704 437560
rect 78456 437520 78462 437532
rect 80698 437520 80704 437532
rect 80756 437520 80762 437572
rect 46566 437452 46572 437504
rect 46624 437492 46630 437504
rect 46750 437492 46756 437504
rect 46624 437464 46756 437492
rect 46624 437452 46630 437464
rect 46750 437452 46756 437464
rect 46808 437452 46814 437504
rect 79042 437452 79048 437504
rect 79100 437492 79106 437504
rect 80054 437492 80060 437504
rect 79100 437464 80060 437492
rect 79100 437452 79106 437464
rect 80054 437452 80060 437464
rect 80112 437452 80118 437504
rect 83642 437452 83648 437504
rect 83700 437492 83706 437504
rect 84838 437492 84844 437504
rect 83700 437464 84844 437492
rect 83700 437452 83706 437464
rect 84838 437452 84844 437464
rect 84896 437452 84902 437504
rect 85022 437452 85028 437504
rect 85080 437492 85086 437504
rect 86770 437492 86776 437504
rect 85080 437464 86776 437492
rect 85080 437452 85086 437464
rect 86770 437452 86776 437464
rect 86828 437452 86834 437504
rect 57514 437384 57520 437436
rect 57572 437424 57578 437436
rect 91738 437424 91744 437436
rect 57572 437396 91744 437424
rect 57572 437384 57578 437396
rect 91738 437384 91744 437396
rect 91796 437384 91802 437436
rect 94498 437384 94504 437436
rect 94556 437424 94562 437436
rect 125778 437424 125784 437436
rect 94556 437396 125784 437424
rect 94556 437384 94562 437396
rect 125778 437384 125784 437396
rect 125836 437384 125842 437436
rect 42610 437316 42616 437368
rect 42668 437356 42674 437368
rect 73338 437356 73344 437368
rect 42668 437328 73344 437356
rect 42668 437316 42674 437328
rect 73338 437316 73344 437328
rect 73396 437316 73402 437368
rect 86218 437316 86224 437368
rect 86276 437356 86282 437368
rect 100018 437356 100024 437368
rect 86276 437328 100024 437356
rect 86276 437316 86282 437328
rect 100018 437316 100024 437328
rect 100076 437316 100082 437368
rect 52362 437248 52368 437300
rect 52420 437288 52426 437300
rect 82906 437288 82912 437300
rect 52420 437260 82912 437288
rect 52420 437248 52426 437260
rect 82906 437248 82912 437260
rect 82964 437248 82970 437300
rect 64138 436704 64144 436756
rect 64196 436744 64202 436756
rect 75270 436744 75276 436756
rect 64196 436716 75276 436744
rect 64196 436704 64202 436716
rect 75270 436704 75276 436716
rect 75328 436704 75334 436756
rect 47946 436024 47952 436076
rect 48004 436064 48010 436076
rect 80054 436064 80060 436076
rect 48004 436036 80060 436064
rect 48004 436024 48010 436036
rect 80054 436024 80060 436036
rect 80112 436024 80118 436076
rect 88242 436024 88248 436076
rect 88300 436064 88306 436076
rect 111794 436064 111800 436076
rect 88300 436036 111800 436064
rect 88300 436024 88306 436036
rect 111794 436024 111800 436036
rect 111852 436024 111858 436076
rect 54846 435956 54852 436008
rect 54904 435996 54910 436008
rect 83090 435996 83096 436008
rect 54904 435968 83096 435996
rect 54904 435956 54910 435968
rect 83090 435956 83096 435968
rect 83148 435996 83154 436008
rect 83642 435996 83648 436008
rect 83148 435968 83648 435996
rect 83148 435956 83154 435968
rect 83642 435956 83648 435968
rect 83700 435956 83706 436008
rect 60366 435888 60372 435940
rect 60424 435928 60430 435940
rect 84194 435928 84200 435940
rect 60424 435900 84200 435928
rect 60424 435888 60430 435900
rect 84194 435888 84200 435900
rect 84252 435928 84258 435940
rect 85022 435928 85028 435940
rect 84252 435900 85028 435928
rect 84252 435888 84258 435900
rect 85022 435888 85028 435900
rect 85080 435888 85086 435940
rect 38470 434664 38476 434716
rect 38528 434704 38534 434716
rect 71314 434704 71320 434716
rect 38528 434676 71320 434704
rect 38528 434664 38534 434676
rect 71314 434664 71320 434676
rect 71372 434664 71378 434716
rect 48958 433984 48964 434036
rect 49016 434024 49022 434036
rect 76466 434024 76472 434036
rect 49016 433996 76472 434024
rect 49016 433984 49022 433996
rect 76466 433984 76472 433996
rect 76524 433984 76530 434036
rect 80698 431196 80704 431248
rect 80756 431236 80762 431248
rect 580166 431236 580172 431248
rect 80756 431208 580172 431236
rect 80756 431196 80762 431208
rect 580166 431196 580172 431208
rect 580224 431196 580230 431248
rect 3418 429836 3424 429888
rect 3476 429876 3482 429888
rect 100846 429876 100852 429888
rect 3476 429848 100852 429876
rect 3476 429836 3482 429848
rect 100846 429836 100852 429848
rect 100904 429836 100910 429888
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 48130 422328 48136 422340
rect 3568 422300 48136 422328
rect 3568 422288 3574 422300
rect 48130 422288 48136 422300
rect 48188 422328 48194 422340
rect 48188 422300 100524 422328
rect 48188 422288 48194 422300
rect 100496 422260 100524 422300
rect 100662 422260 100668 422272
rect 100496 422232 100668 422260
rect 100662 422220 100668 422232
rect 100720 422260 100726 422272
rect 124306 422260 124312 422272
rect 100720 422232 124312 422260
rect 100720 422220 100726 422232
rect 124306 422220 124312 422232
rect 124364 422220 124370 422272
rect 66990 419432 66996 419484
rect 67048 419472 67054 419484
rect 67358 419472 67364 419484
rect 67048 419444 67364 419472
rect 67048 419432 67054 419444
rect 67358 419432 67364 419444
rect 67416 419472 67422 419484
rect 580166 419472 580172 419484
rect 67416 419444 580172 419472
rect 67416 419432 67422 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 56410 418752 56416 418804
rect 56468 418792 56474 418804
rect 67358 418792 67364 418804
rect 56468 418764 67364 418792
rect 56468 418752 56474 418764
rect 67358 418752 67364 418764
rect 67416 418752 67422 418804
rect 91830 404336 91836 404388
rect 91888 404376 91894 404388
rect 580166 404376 580172 404388
rect 91888 404348 580172 404376
rect 91888 404336 91894 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 108298 402364 108304 402416
rect 108356 402404 108362 402416
rect 117590 402404 117596 402416
rect 108356 402376 117596 402404
rect 108356 402364 108362 402376
rect 117590 402364 117596 402376
rect 117648 402364 117654 402416
rect 96614 402296 96620 402348
rect 96672 402336 96678 402348
rect 127158 402336 127164 402348
rect 96672 402308 127164 402336
rect 96672 402296 96678 402308
rect 127158 402296 127164 402308
rect 127216 402296 127222 402348
rect 88242 402228 88248 402280
rect 88300 402268 88306 402280
rect 124306 402268 124312 402280
rect 88300 402240 124312 402268
rect 88300 402228 88306 402240
rect 124306 402228 124312 402240
rect 124364 402228 124370 402280
rect 108850 401616 108856 401668
rect 108908 401656 108914 401668
rect 113450 401656 113456 401668
rect 108908 401628 113456 401656
rect 108908 401616 108914 401628
rect 113450 401616 113456 401628
rect 113508 401616 113514 401668
rect 74626 400188 74632 400240
rect 74684 400228 74690 400240
rect 75270 400228 75276 400240
rect 74684 400200 75276 400228
rect 74684 400188 74690 400200
rect 75270 400188 75276 400200
rect 75328 400228 75334 400240
rect 162118 400228 162124 400240
rect 75328 400200 162124 400228
rect 75328 400188 75334 400200
rect 162118 400188 162124 400200
rect 162176 400188 162182 400240
rect 104158 399508 104164 399560
rect 104216 399548 104222 399560
rect 138198 399548 138204 399560
rect 104216 399520 138204 399548
rect 104216 399508 104222 399520
rect 138198 399508 138204 399520
rect 138256 399508 138262 399560
rect 35158 399440 35164 399492
rect 35216 399480 35222 399492
rect 75914 399480 75920 399492
rect 35216 399452 75920 399480
rect 35216 399440 35222 399452
rect 75914 399440 75920 399452
rect 75972 399440 75978 399492
rect 98638 399440 98644 399492
rect 98696 399480 98702 399492
rect 135346 399480 135352 399492
rect 98696 399452 135352 399480
rect 98696 399440 98702 399452
rect 135346 399440 135352 399452
rect 135404 399440 135410 399492
rect 99374 398216 99380 398268
rect 99432 398256 99438 398268
rect 118878 398256 118884 398268
rect 99432 398228 118884 398256
rect 99432 398216 99438 398228
rect 118878 398216 118884 398228
rect 118936 398216 118942 398268
rect 89622 398148 89628 398200
rect 89680 398188 89686 398200
rect 122098 398188 122104 398200
rect 89680 398160 122104 398188
rect 89680 398148 89686 398160
rect 122098 398148 122104 398160
rect 122156 398148 122162 398200
rect 50982 398080 50988 398132
rect 51040 398120 51046 398132
rect 99374 398120 99380 398132
rect 51040 398092 99380 398120
rect 51040 398080 51046 398092
rect 99374 398080 99380 398092
rect 99432 398080 99438 398132
rect 106918 398080 106924 398132
rect 106976 398120 106982 398132
rect 141050 398120 141056 398132
rect 106976 398092 141056 398120
rect 106976 398080 106982 398092
rect 141050 398080 141056 398092
rect 141108 398080 141114 398132
rect 92474 397536 92480 397588
rect 92532 397576 92538 397588
rect 92658 397576 92664 397588
rect 92532 397548 92664 397576
rect 92532 397536 92538 397548
rect 92658 397536 92664 397548
rect 92716 397576 92722 397588
rect 220078 397576 220084 397588
rect 92716 397548 220084 397576
rect 92716 397536 92722 397548
rect 220078 397536 220084 397548
rect 220136 397536 220142 397588
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 50982 397508 50988 397520
rect 3476 397480 50988 397508
rect 3476 397468 3482 397480
rect 50982 397468 50988 397480
rect 51040 397468 51046 397520
rect 65978 397468 65984 397520
rect 66036 397508 66042 397520
rect 269758 397508 269764 397520
rect 66036 397480 269764 397508
rect 66036 397468 66042 397480
rect 269758 397468 269764 397480
rect 269816 397468 269822 397520
rect 46566 396856 46572 396908
rect 46624 396896 46630 396908
rect 80054 396896 80060 396908
rect 46624 396868 80060 396896
rect 46624 396856 46630 396868
rect 80054 396856 80060 396868
rect 80112 396856 80118 396908
rect 105630 396856 105636 396908
rect 105688 396896 105694 396908
rect 131298 396896 131304 396908
rect 105688 396868 131304 396896
rect 105688 396856 105694 396868
rect 131298 396856 131304 396868
rect 131356 396856 131362 396908
rect 53558 396788 53564 396840
rect 53616 396828 53622 396840
rect 80698 396828 80704 396840
rect 53616 396800 80704 396828
rect 53616 396788 53622 396800
rect 80698 396788 80704 396800
rect 80756 396788 80762 396840
rect 91738 396788 91744 396840
rect 91796 396828 91802 396840
rect 127250 396828 127256 396840
rect 91796 396800 127256 396828
rect 91796 396788 91802 396800
rect 127250 396788 127256 396800
rect 127308 396788 127314 396840
rect 46658 396720 46664 396772
rect 46716 396760 46722 396772
rect 91922 396760 91928 396772
rect 46716 396732 91928 396760
rect 46716 396720 46722 396732
rect 91922 396720 91928 396732
rect 91980 396720 91986 396772
rect 93854 396720 93860 396772
rect 93912 396760 93918 396772
rect 123110 396760 123116 396772
rect 93912 396732 123116 396760
rect 93912 396720 93918 396732
rect 123110 396720 123116 396732
rect 123168 396720 123174 396772
rect 53466 396040 53472 396092
rect 53524 396080 53530 396092
rect 54478 396080 54484 396092
rect 53524 396052 54484 396080
rect 53524 396040 53530 396052
rect 54478 396040 54484 396052
rect 54536 396080 54542 396092
rect 84194 396080 84200 396092
rect 54536 396052 84200 396080
rect 54536 396040 54542 396052
rect 84194 396040 84200 396052
rect 84252 396040 84258 396092
rect 85114 396040 85120 396092
rect 85172 396080 85178 396092
rect 166258 396080 166264 396092
rect 85172 396052 166264 396080
rect 85172 396040 85178 396052
rect 166258 396040 166264 396052
rect 166316 396040 166322 396092
rect 49510 395292 49516 395344
rect 49568 395332 49574 395344
rect 88334 395332 88340 395344
rect 49568 395304 88340 395332
rect 49568 395292 49574 395304
rect 88334 395292 88340 395304
rect 88392 395292 88398 395344
rect 97902 395292 97908 395344
rect 97960 395332 97966 395344
rect 121638 395332 121644 395344
rect 97960 395304 121644 395332
rect 97960 395292 97966 395304
rect 121638 395292 121644 395304
rect 121696 395332 121702 395344
rect 317414 395332 317420 395344
rect 121696 395304 317420 395332
rect 121696 395292 121702 395304
rect 317414 395292 317420 395304
rect 317472 395292 317478 395344
rect 70394 394952 70400 395004
rect 70452 394992 70458 395004
rect 71130 394992 71136 395004
rect 70452 394964 71136 394992
rect 70452 394952 70458 394964
rect 71130 394952 71136 394964
rect 71188 394952 71194 395004
rect 39758 394884 39764 394936
rect 39816 394924 39822 394936
rect 103698 394924 103704 394936
rect 39816 394896 103704 394924
rect 39816 394884 39822 394896
rect 103698 394884 103704 394896
rect 103756 394924 103762 394936
rect 104250 394924 104256 394936
rect 103756 394896 104256 394924
rect 103756 394884 103762 394896
rect 104250 394884 104256 394896
rect 104308 394884 104314 394936
rect 66070 394816 66076 394868
rect 66128 394856 66134 394868
rect 142154 394856 142160 394868
rect 66128 394828 142160 394856
rect 66128 394816 66134 394828
rect 142154 394816 142160 394828
rect 142212 394816 142218 394868
rect 88334 394748 88340 394800
rect 88392 394788 88398 394800
rect 170398 394788 170404 394800
rect 88392 394760 170404 394788
rect 88392 394748 88398 394760
rect 170398 394748 170404 394760
rect 170456 394748 170462 394800
rect 71130 394680 71136 394732
rect 71188 394720 71194 394732
rect 214558 394720 214564 394732
rect 71188 394692 214564 394720
rect 71188 394680 71194 394692
rect 214558 394680 214564 394692
rect 214616 394680 214622 394732
rect 77938 394612 77944 394664
rect 77996 394652 78002 394664
rect 91830 394652 91836 394664
rect 77996 394624 91836 394652
rect 77996 394612 78002 394624
rect 91830 394612 91836 394624
rect 91888 394612 91894 394664
rect 47854 394136 47860 394188
rect 47912 394176 47918 394188
rect 56226 394176 56232 394188
rect 47912 394148 56232 394176
rect 47912 394136 47918 394148
rect 56226 394136 56232 394148
rect 56284 394176 56290 394188
rect 66070 394176 66076 394188
rect 56284 394148 66076 394176
rect 56284 394136 56290 394148
rect 66070 394136 66076 394148
rect 66128 394136 66134 394188
rect 52086 394068 52092 394120
rect 52144 394108 52150 394120
rect 82906 394108 82912 394120
rect 52144 394080 82912 394108
rect 52144 394068 52150 394080
rect 82906 394068 82912 394080
rect 82964 394068 82970 394120
rect 47946 394000 47952 394052
rect 48004 394040 48010 394052
rect 79318 394040 79324 394052
rect 48004 394012 79324 394040
rect 48004 394000 48010 394012
rect 79318 394000 79324 394012
rect 79376 394000 79382 394052
rect 43990 393932 43996 393984
rect 44048 393972 44054 393984
rect 81434 393972 81440 393984
rect 44048 393944 81440 393972
rect 44048 393932 44054 393944
rect 81434 393932 81440 393944
rect 81492 393932 81498 393984
rect 87690 393932 87696 393984
rect 87748 393972 87754 393984
rect 110414 393972 110420 393984
rect 87748 393944 110420 393972
rect 87748 393932 87754 393944
rect 110414 393932 110420 393944
rect 110472 393932 110478 393984
rect 43990 393456 43996 393508
rect 44048 393496 44054 393508
rect 101398 393496 101404 393508
rect 44048 393468 101404 393496
rect 44048 393456 44054 393468
rect 101398 393456 101404 393468
rect 101456 393456 101462 393508
rect 81434 393388 81440 393440
rect 81492 393428 81498 393440
rect 151998 393428 152004 393440
rect 81492 393400 152004 393428
rect 81492 393388 81498 393400
rect 151998 393388 152004 393400
rect 152056 393388 152062 393440
rect 75914 393320 75920 393372
rect 75972 393360 75978 393372
rect 159358 393360 159364 393372
rect 75972 393332 159364 393360
rect 75972 393320 75978 393332
rect 159358 393320 159364 393332
rect 159416 393320 159422 393372
rect 110414 392776 110420 392828
rect 110472 392816 110478 392828
rect 123202 392816 123208 392828
rect 110472 392788 123208 392816
rect 110472 392776 110478 392788
rect 123202 392776 123208 392788
rect 123260 392776 123266 392828
rect 96522 392708 96528 392760
rect 96580 392748 96586 392760
rect 125870 392748 125876 392760
rect 96580 392720 125876 392748
rect 96580 392708 96586 392720
rect 125870 392708 125876 392720
rect 125928 392708 125934 392760
rect 57698 392640 57704 392692
rect 57756 392680 57762 392692
rect 88426 392680 88432 392692
rect 57756 392652 88432 392680
rect 57756 392640 57762 392652
rect 88426 392640 88432 392652
rect 88484 392640 88490 392692
rect 96246 392640 96252 392692
rect 96304 392680 96310 392692
rect 130010 392680 130016 392692
rect 96304 392652 130016 392680
rect 96304 392640 96310 392652
rect 130010 392640 130016 392652
rect 130068 392680 130074 392692
rect 140958 392680 140964 392692
rect 130068 392652 140964 392680
rect 130068 392640 130074 392652
rect 140958 392640 140964 392652
rect 141016 392640 141022 392692
rect 45278 392572 45284 392624
rect 45336 392612 45342 392624
rect 78674 392612 78680 392624
rect 45336 392584 78680 392612
rect 45336 392572 45342 392584
rect 78674 392572 78680 392584
rect 78732 392572 78738 392624
rect 99282 392572 99288 392624
rect 99340 392612 99346 392624
rect 135438 392612 135444 392624
rect 99340 392584 135444 392612
rect 99340 392572 99346 392584
rect 135438 392572 135444 392584
rect 135496 392572 135502 392624
rect 113082 392436 113088 392488
rect 113140 392476 113146 392488
rect 114554 392476 114560 392488
rect 113140 392448 114560 392476
rect 113140 392436 113146 392448
rect 114554 392436 114560 392448
rect 114612 392436 114618 392488
rect 46842 392028 46848 392080
rect 46900 392068 46906 392080
rect 92934 392068 92940 392080
rect 46900 392040 92940 392068
rect 46900 392028 46906 392040
rect 92934 392028 92940 392040
rect 92992 392028 92998 392080
rect 52270 391960 52276 392012
rect 52328 392000 52334 392012
rect 110414 392000 110420 392012
rect 52328 391972 110420 392000
rect 52328 391960 52334 391972
rect 110414 391960 110420 391972
rect 110472 392000 110478 392012
rect 110966 392000 110972 392012
rect 110472 391972 110972 392000
rect 110472 391960 110478 391972
rect 110966 391960 110972 391972
rect 111024 391960 111030 392012
rect 111058 391960 111064 392012
rect 111116 392000 111122 392012
rect 112070 392000 112076 392012
rect 111116 391972 112076 392000
rect 111116 391960 111122 391972
rect 112070 391960 112076 391972
rect 112128 391960 112134 392012
rect 113818 391960 113824 392012
rect 113876 392000 113882 392012
rect 177298 392000 177304 392012
rect 113876 391972 177304 392000
rect 113876 391960 113882 391972
rect 177298 391960 177304 391972
rect 177356 391960 177362 392012
rect 60550 391484 60556 391536
rect 60608 391524 60614 391536
rect 82814 391524 82820 391536
rect 60608 391496 82820 391524
rect 60608 391484 60614 391496
rect 82814 391484 82820 391496
rect 82872 391484 82878 391536
rect 54754 391348 54760 391400
rect 54812 391388 54818 391400
rect 82814 391388 82820 391400
rect 54812 391360 82820 391388
rect 54812 391348 54818 391360
rect 82814 391348 82820 391360
rect 82872 391348 82878 391400
rect 100662 391348 100668 391400
rect 100720 391388 100726 391400
rect 115382 391388 115388 391400
rect 100720 391360 115388 391388
rect 100720 391348 100726 391360
rect 115382 391348 115388 391360
rect 115440 391348 115446 391400
rect 60366 391280 60372 391332
rect 60424 391320 60430 391332
rect 94498 391320 94504 391332
rect 60424 391292 94504 391320
rect 60424 391280 60430 391292
rect 94498 391280 94504 391292
rect 94556 391280 94562 391332
rect 102042 391280 102048 391332
rect 102100 391320 102106 391332
rect 120350 391320 120356 391332
rect 102100 391292 120356 391320
rect 102100 391280 102106 391292
rect 120350 391280 120356 391292
rect 120408 391280 120414 391332
rect 41230 391212 41236 391264
rect 41288 391252 41294 391264
rect 85942 391252 85948 391264
rect 41288 391224 85948 391252
rect 41288 391212 41294 391224
rect 85942 391212 85948 391224
rect 86000 391212 86006 391264
rect 94130 391212 94136 391264
rect 94188 391252 94194 391264
rect 121454 391252 121460 391264
rect 94188 391224 121460 391252
rect 94188 391212 94194 391224
rect 121454 391212 121460 391224
rect 121512 391252 121518 391264
rect 147858 391252 147864 391264
rect 121512 391224 147864 391252
rect 121512 391212 121518 391224
rect 147858 391212 147864 391224
rect 147916 391212 147922 391264
rect 119338 390668 119344 390720
rect 119396 390708 119402 390720
rect 124214 390708 124220 390720
rect 119396 390680 124220 390708
rect 119396 390668 119402 390680
rect 124214 390668 124220 390680
rect 124272 390668 124278 390720
rect 82906 390600 82912 390652
rect 82964 390640 82970 390652
rect 83642 390640 83648 390652
rect 82964 390612 83648 390640
rect 82964 390600 82970 390612
rect 83642 390600 83648 390612
rect 83700 390640 83706 390652
rect 139394 390640 139400 390652
rect 83700 390612 139400 390640
rect 83700 390600 83706 390612
rect 139394 390600 139400 390612
rect 139452 390600 139458 390652
rect 82814 390532 82820 390584
rect 82872 390572 82878 390584
rect 82998 390572 83004 390584
rect 82872 390544 83004 390572
rect 82872 390532 82878 390544
rect 82998 390532 83004 390544
rect 83056 390572 83062 390584
rect 143718 390572 143724 390584
rect 83056 390544 143724 390572
rect 83056 390532 83062 390544
rect 143718 390532 143724 390544
rect 143776 390532 143782 390584
rect 124122 389988 124128 390040
rect 124180 390028 124186 390040
rect 135254 390028 135260 390040
rect 124180 390000 135260 390028
rect 124180 389988 124186 390000
rect 135254 389988 135260 390000
rect 135312 389988 135318 390040
rect 97442 389920 97448 389972
rect 97500 389960 97506 389972
rect 130102 389960 130108 389972
rect 97500 389932 130108 389960
rect 97500 389920 97506 389932
rect 130102 389920 130108 389932
rect 130160 389960 130166 389972
rect 146294 389960 146300 389972
rect 130160 389932 146300 389960
rect 130160 389920 130166 389932
rect 146294 389920 146300 389932
rect 146352 389920 146358 389972
rect 53650 389852 53656 389904
rect 53708 389892 53714 389904
rect 59262 389892 59268 389904
rect 53708 389864 59268 389892
rect 53708 389852 53714 389864
rect 59262 389852 59268 389864
rect 59320 389892 59326 389904
rect 104526 389892 104532 389904
rect 59320 389864 104532 389892
rect 59320 389852 59326 389864
rect 104526 389852 104532 389864
rect 104584 389852 104590 389904
rect 108942 389852 108948 389904
rect 109000 389892 109006 389904
rect 131206 389892 131212 389904
rect 109000 389864 131212 389892
rect 109000 389852 109006 389864
rect 131206 389852 131212 389864
rect 131264 389892 131270 389904
rect 134150 389892 134156 389904
rect 131264 389864 134156 389892
rect 131264 389852 131270 389864
rect 134150 389852 134156 389864
rect 134208 389852 134214 389904
rect 49050 389784 49056 389836
rect 49108 389824 49114 389836
rect 119338 389824 119344 389836
rect 49108 389796 119344 389824
rect 49108 389784 49114 389796
rect 119338 389784 119344 389796
rect 119396 389784 119402 389836
rect 106274 389240 106280 389292
rect 106332 389280 106338 389292
rect 122834 389280 122840 389292
rect 106332 389252 122840 389280
rect 106332 389240 106338 389252
rect 122834 389240 122840 389252
rect 122892 389280 122898 389292
rect 124122 389280 124128 389292
rect 122892 389252 124128 389280
rect 122892 389240 122898 389252
rect 124122 389240 124128 389252
rect 124180 389240 124186 389292
rect 39850 389172 39856 389224
rect 39908 389212 39914 389224
rect 71774 389212 71780 389224
rect 39908 389184 71780 389212
rect 39908 389172 39914 389184
rect 71774 389172 71780 389184
rect 71832 389172 71838 389224
rect 114370 389172 114376 389224
rect 114428 389212 114434 389224
rect 142430 389212 142436 389224
rect 114428 389184 142436 389212
rect 114428 389172 114434 389184
rect 142430 389172 142436 389184
rect 142488 389172 142494 389224
rect 101398 389104 101404 389156
rect 101456 389144 101462 389156
rect 103606 389144 103612 389156
rect 101456 389116 103612 389144
rect 101456 389104 101462 389116
rect 103606 389104 103612 389116
rect 103664 389104 103670 389156
rect 120626 389104 120632 389156
rect 120684 389144 120690 389156
rect 127066 389144 127072 389156
rect 120684 389116 127072 389144
rect 120684 389104 120690 389116
rect 127066 389104 127072 389116
rect 127124 389104 127130 389156
rect 71866 388832 71872 388884
rect 71924 388872 71930 388884
rect 72326 388872 72332 388884
rect 71924 388844 72332 388872
rect 71924 388832 71930 388844
rect 72326 388832 72332 388844
rect 72384 388832 72390 388884
rect 101858 388492 101864 388544
rect 101916 388532 101922 388544
rect 113082 388532 113088 388544
rect 101916 388504 113088 388532
rect 101916 388492 101922 388504
rect 113082 388492 113088 388504
rect 113140 388532 113146 388544
rect 122282 388532 122288 388544
rect 113140 388504 122288 388532
rect 113140 388492 113146 388504
rect 122282 388492 122288 388504
rect 122340 388492 122346 388544
rect 57330 388424 57336 388476
rect 57388 388464 57394 388476
rect 75822 388464 75828 388476
rect 57388 388436 75828 388464
rect 57388 388424 57394 388436
rect 75822 388424 75828 388436
rect 75880 388424 75886 388476
rect 107010 388424 107016 388476
rect 107068 388464 107074 388476
rect 111702 388464 111708 388476
rect 107068 388436 111708 388464
rect 107068 388424 107074 388436
rect 111702 388424 111708 388436
rect 111760 388464 111766 388476
rect 124950 388464 124956 388476
rect 111760 388436 124956 388464
rect 111760 388424 111766 388436
rect 124950 388424 124956 388436
rect 125008 388424 125014 388476
rect 55030 388084 55036 388136
rect 55088 388124 55094 388136
rect 69750 388124 69756 388136
rect 55088 388096 69756 388124
rect 55088 388084 55094 388096
rect 69750 388084 69756 388096
rect 69808 388084 69814 388136
rect 75178 388084 75184 388136
rect 75236 388124 75242 388136
rect 75546 388124 75552 388136
rect 75236 388096 75552 388124
rect 75236 388084 75242 388096
rect 75546 388084 75552 388096
rect 75604 388124 75610 388136
rect 82446 388124 82452 388136
rect 75604 388096 82452 388124
rect 75604 388084 75610 388096
rect 82446 388084 82452 388096
rect 82504 388084 82510 388136
rect 109678 388084 109684 388136
rect 109736 388124 109742 388136
rect 119338 388124 119344 388136
rect 109736 388096 119344 388124
rect 109736 388084 109742 388096
rect 119338 388084 119344 388096
rect 119396 388084 119402 388136
rect 59170 388016 59176 388068
rect 59228 388056 59234 388068
rect 79318 388056 79324 388068
rect 59228 388028 79324 388056
rect 59228 388016 59234 388028
rect 79318 388016 79324 388028
rect 79376 388016 79382 388068
rect 100018 388016 100024 388068
rect 100076 388056 100082 388068
rect 120626 388056 120632 388068
rect 100076 388028 120632 388056
rect 100076 388016 100082 388028
rect 120626 388016 120632 388028
rect 120684 388016 120690 388068
rect 56502 387948 56508 388000
rect 56560 387988 56566 388000
rect 78030 387988 78036 388000
rect 56560 387960 78036 387988
rect 56560 387948 56566 387960
rect 78030 387948 78036 387960
rect 78088 387948 78094 388000
rect 91002 387948 91008 388000
rect 91060 387988 91066 388000
rect 121914 387988 121920 388000
rect 91060 387960 121920 387988
rect 91060 387948 91066 387960
rect 121914 387948 121920 387960
rect 121972 387948 121978 388000
rect 25498 387880 25504 387932
rect 25556 387920 25562 387932
rect 41230 387920 41236 387932
rect 25556 387892 41236 387920
rect 25556 387880 25562 387892
rect 41230 387880 41236 387892
rect 41288 387920 41294 387932
rect 72326 387920 72332 387932
rect 41288 387892 72332 387920
rect 41288 387880 41294 387892
rect 72326 387880 72332 387892
rect 72384 387880 72390 387932
rect 75822 387880 75828 387932
rect 75880 387920 75886 387932
rect 113082 387920 113088 387932
rect 75880 387892 113088 387920
rect 75880 387880 75886 387892
rect 113082 387880 113088 387892
rect 113140 387880 113146 387932
rect 35802 387812 35808 387864
rect 35860 387852 35866 387864
rect 80054 387852 80060 387864
rect 35860 387824 80060 387852
rect 35860 387812 35866 387824
rect 80054 387812 80060 387824
rect 80112 387812 80118 387864
rect 90266 387812 90272 387864
rect 90324 387852 90330 387864
rect 98822 387852 98828 387864
rect 90324 387824 98828 387852
rect 90324 387812 90330 387824
rect 98822 387812 98828 387824
rect 98880 387812 98886 387864
rect 112070 387812 112076 387864
rect 112128 387852 112134 387864
rect 188338 387852 188344 387864
rect 112128 387824 188344 387852
rect 112128 387812 112134 387824
rect 188338 387812 188344 387824
rect 188396 387812 188402 387864
rect 53742 387472 53748 387524
rect 53800 387512 53806 387524
rect 56502 387512 56508 387524
rect 53800 387484 56508 387512
rect 53800 387472 53806 387484
rect 56502 387472 56508 387484
rect 56560 387472 56566 387524
rect 113082 387268 113088 387320
rect 113140 387308 113146 387320
rect 132586 387308 132592 387320
rect 113140 387280 132592 387308
rect 113140 387268 113146 387280
rect 132586 387268 132592 387280
rect 132644 387268 132650 387320
rect 105538 387200 105544 387252
rect 105596 387240 105602 387252
rect 131206 387240 131212 387252
rect 105596 387212 131212 387240
rect 105596 387200 105602 387212
rect 131206 387200 131212 387212
rect 131264 387200 131270 387252
rect 57606 387132 57612 387184
rect 57664 387172 57670 387184
rect 74534 387172 74540 387184
rect 57664 387144 74540 387172
rect 57664 387132 57670 387144
rect 74534 387132 74540 387144
rect 74592 387132 74598 387184
rect 90910 387132 90916 387184
rect 90968 387172 90974 387184
rect 125778 387172 125784 387184
rect 90968 387144 125784 387172
rect 90968 387132 90974 387144
rect 125778 387132 125784 387144
rect 125836 387132 125842 387184
rect 128630 387132 128636 387184
rect 128688 387172 128694 387184
rect 143534 387172 143540 387184
rect 128688 387144 143540 387172
rect 128688 387132 128694 387144
rect 143534 387132 143540 387144
rect 143592 387132 143598 387184
rect 58894 387064 58900 387116
rect 58952 387104 58958 387116
rect 90358 387104 90364 387116
rect 58952 387076 90364 387104
rect 58952 387064 58958 387076
rect 90358 387064 90364 387076
rect 90416 387064 90422 387116
rect 94866 387064 94872 387116
rect 94924 387104 94930 387116
rect 108850 387104 108856 387116
rect 94924 387076 108856 387104
rect 94924 387064 94930 387076
rect 108850 387064 108856 387076
rect 108908 387104 108914 387116
rect 215938 387104 215944 387116
rect 108908 387076 215944 387104
rect 108908 387064 108914 387076
rect 215938 387064 215944 387076
rect 215996 387064 216002 387116
rect 52362 386452 52368 386504
rect 52420 386492 52426 386504
rect 53466 386492 53472 386504
rect 52420 386464 53472 386492
rect 52420 386452 52426 386464
rect 53466 386452 53472 386464
rect 53524 386492 53530 386504
rect 80606 386492 80612 386504
rect 53524 386464 80612 386492
rect 53524 386452 53530 386464
rect 80606 386452 80612 386464
rect 80664 386452 80670 386504
rect 112898 386452 112904 386504
rect 112956 386492 112962 386504
rect 128630 386492 128636 386504
rect 112956 386464 128636 386492
rect 112956 386452 112962 386464
rect 128630 386452 128636 386464
rect 128688 386452 128694 386504
rect 57882 386384 57888 386436
rect 57940 386424 57946 386436
rect 87046 386424 87052 386436
rect 57940 386396 87052 386424
rect 57940 386384 57946 386396
rect 87046 386384 87052 386396
rect 87104 386384 87110 386436
rect 110322 386384 110328 386436
rect 110380 386424 110386 386436
rect 136634 386424 136640 386436
rect 110380 386396 136640 386424
rect 110380 386384 110386 386396
rect 136634 386384 136640 386396
rect 136692 386384 136698 386436
rect 61746 386316 61752 386368
rect 61804 386356 61810 386368
rect 68830 386356 68836 386368
rect 61804 386328 68836 386356
rect 61804 386316 61810 386328
rect 68830 386316 68836 386328
rect 68888 386316 68894 386368
rect 135254 386316 135260 386368
rect 135312 386356 135318 386368
rect 138014 386356 138020 386368
rect 135312 386328 138020 386356
rect 135312 386316 135318 386328
rect 138014 386316 138020 386328
rect 138072 386316 138078 386368
rect 61654 385840 61660 385892
rect 61712 385880 61718 385892
rect 73430 385880 73436 385892
rect 61712 385852 73436 385880
rect 61712 385840 61718 385852
rect 73430 385840 73436 385852
rect 73488 385840 73494 385892
rect 70302 385772 70308 385824
rect 70360 385812 70366 385824
rect 83090 385812 83096 385824
rect 70360 385784 83096 385812
rect 70360 385772 70366 385784
rect 83090 385772 83096 385784
rect 83148 385772 83154 385824
rect 59078 385704 59084 385756
rect 59136 385744 59142 385756
rect 59136 385716 74534 385744
rect 59136 385704 59142 385716
rect 56318 385636 56324 385688
rect 56376 385676 56382 385688
rect 73430 385676 73436 385688
rect 56376 385648 73436 385676
rect 56376 385636 56382 385648
rect 73430 385636 73436 385648
rect 73488 385636 73494 385688
rect 74506 385608 74534 385716
rect 112990 385704 112996 385756
rect 113048 385744 113054 385756
rect 122926 385744 122932 385756
rect 113048 385716 122932 385744
rect 113048 385704 113054 385716
rect 122926 385704 122932 385716
rect 122984 385704 122990 385756
rect 82446 385636 82452 385688
rect 82504 385676 82510 385688
rect 303614 385676 303620 385688
rect 82504 385648 303620 385676
rect 82504 385636 82510 385648
rect 303614 385636 303620 385648
rect 303672 385636 303678 385688
rect 86310 385608 86316 385620
rect 74506 385580 86316 385608
rect 86310 385568 86316 385580
rect 86368 385568 86374 385620
rect 117314 385432 117320 385484
rect 117372 385472 117378 385484
rect 117682 385472 117688 385484
rect 117372 385444 117688 385472
rect 117372 385432 117378 385444
rect 117682 385432 117688 385444
rect 117740 385432 117746 385484
rect 77478 385336 77484 385348
rect 64846 385308 77484 385336
rect 56502 385024 56508 385076
rect 56560 385064 56566 385076
rect 64846 385064 64874 385308
rect 77478 385296 77484 385308
rect 77536 385296 77542 385348
rect 102594 385296 102600 385348
rect 102652 385336 102658 385348
rect 102652 385308 103514 385336
rect 102652 385296 102658 385308
rect 56560 385036 64874 385064
rect 103486 385064 103514 385308
rect 107562 385296 107568 385348
rect 107620 385336 107626 385348
rect 107620 385308 109034 385336
rect 107620 385296 107626 385308
rect 109006 385132 109034 385308
rect 135254 385132 135260 385144
rect 109006 385104 135260 385132
rect 135254 385092 135260 385104
rect 135312 385092 135318 385144
rect 133874 385064 133880 385076
rect 103486 385036 133880 385064
rect 56560 385024 56566 385036
rect 133874 385024 133880 385036
rect 133932 385064 133938 385076
rect 134610 385064 134616 385076
rect 133932 385036 134616 385064
rect 133932 385024 133938 385036
rect 134610 385024 134616 385036
rect 134668 385024 134674 385076
rect 117406 384888 117412 384940
rect 117464 384888 117470 384940
rect 118234 384888 118240 384940
rect 118292 384928 118298 384940
rect 121454 384928 121460 384940
rect 118292 384900 121460 384928
rect 118292 384888 118298 384900
rect 121454 384888 121460 384900
rect 121512 384888 121518 384940
rect 117424 384600 117452 384888
rect 117406 384548 117412 384600
rect 117464 384548 117470 384600
rect 34330 383664 34336 383716
rect 34388 383704 34394 383716
rect 68738 383704 68744 383716
rect 34388 383676 68744 383704
rect 34388 383664 34394 383676
rect 68738 383664 68744 383676
rect 68796 383664 68802 383716
rect 116670 383664 116676 383716
rect 116728 383704 116734 383716
rect 130010 383704 130016 383716
rect 116728 383676 130016 383704
rect 116728 383664 116734 383676
rect 130010 383664 130016 383676
rect 130068 383664 130074 383716
rect 116762 383596 116768 383648
rect 116820 383636 116826 383648
rect 125686 383636 125692 383648
rect 116820 383608 125692 383636
rect 116820 383596 116826 383608
rect 125686 383596 125692 383608
rect 125744 383596 125750 383648
rect 121454 382916 121460 382968
rect 121512 382956 121518 382968
rect 349246 382956 349252 382968
rect 121512 382928 349252 382956
rect 121512 382916 121518 382928
rect 349246 382916 349252 382928
rect 349304 382916 349310 382968
rect 44082 382236 44088 382288
rect 44140 382276 44146 382288
rect 67726 382276 67732 382288
rect 44140 382248 67732 382276
rect 44140 382236 44146 382248
rect 67726 382236 67732 382248
rect 67784 382236 67790 382288
rect 62022 382168 62028 382220
rect 62080 382208 62086 382220
rect 67634 382208 67640 382220
rect 62080 382180 67640 382208
rect 62080 382168 62086 382180
rect 67634 382168 67640 382180
rect 67692 382168 67698 382220
rect 117314 382168 117320 382220
rect 117372 382208 117378 382220
rect 145006 382208 145012 382220
rect 117372 382180 145012 382208
rect 117372 382168 117378 382180
rect 145006 382168 145012 382180
rect 145064 382168 145070 382220
rect 145006 381488 145012 381540
rect 145064 381528 145070 381540
rect 206278 381528 206284 381540
rect 145064 381500 206284 381528
rect 145064 381488 145070 381500
rect 206278 381488 206284 381500
rect 206336 381488 206342 381540
rect 64414 380808 64420 380860
rect 64472 380848 64478 380860
rect 67450 380848 67456 380860
rect 64472 380820 67456 380848
rect 64472 380808 64478 380820
rect 67450 380808 67456 380820
rect 67508 380808 67514 380860
rect 117314 380808 117320 380860
rect 117372 380848 117378 380860
rect 128446 380848 128452 380860
rect 117372 380820 128452 380848
rect 117372 380808 117378 380820
rect 128446 380808 128452 380820
rect 128504 380808 128510 380860
rect 64690 380740 64696 380792
rect 64748 380780 64754 380792
rect 68002 380780 68008 380792
rect 64748 380752 68008 380780
rect 64748 380740 64754 380752
rect 68002 380740 68008 380752
rect 68060 380740 68066 380792
rect 50706 380672 50712 380724
rect 50764 380712 50770 380724
rect 53374 380712 53380 380724
rect 50764 380684 53380 380712
rect 50764 380672 50770 380684
rect 53374 380672 53380 380684
rect 53432 380712 53438 380724
rect 67634 380712 67640 380724
rect 53432 380684 67640 380712
rect 53432 380672 53438 380684
rect 67634 380672 67640 380684
rect 67692 380672 67698 380724
rect 117682 380128 117688 380180
rect 117740 380168 117746 380180
rect 126238 380168 126244 380180
rect 117740 380140 126244 380168
rect 117740 380128 117746 380140
rect 126238 380128 126244 380140
rect 126296 380128 126302 380180
rect 128446 379516 128452 379568
rect 128504 379556 128510 379568
rect 129734 379556 129740 379568
rect 128504 379528 129740 379556
rect 128504 379516 128510 379528
rect 129734 379516 129740 379528
rect 129792 379516 129798 379568
rect 33042 378768 33048 378820
rect 33100 378808 33106 378820
rect 47854 378808 47860 378820
rect 33100 378780 47860 378808
rect 33100 378768 33106 378780
rect 47854 378768 47860 378780
rect 47912 378768 47918 378820
rect 60274 378768 60280 378820
rect 60332 378808 60338 378820
rect 70302 378808 70308 378820
rect 60332 378780 70308 378808
rect 60332 378768 60338 378780
rect 70302 378768 70308 378780
rect 70360 378768 70366 378820
rect 118602 378768 118608 378820
rect 118660 378808 118666 378820
rect 125686 378808 125692 378820
rect 118660 378780 125692 378808
rect 118660 378768 118666 378780
rect 125686 378768 125692 378780
rect 125744 378768 125750 378820
rect 47854 378156 47860 378208
rect 47912 378196 47918 378208
rect 48222 378196 48228 378208
rect 47912 378168 48228 378196
rect 47912 378156 47918 378168
rect 48222 378156 48228 378168
rect 48280 378196 48286 378208
rect 67634 378196 67640 378208
rect 48280 378168 67640 378196
rect 48280 378156 48286 378168
rect 67634 378156 67640 378168
rect 67692 378156 67698 378208
rect 124858 378156 124864 378208
rect 124916 378196 124922 378208
rect 580166 378196 580172 378208
rect 124916 378168 580172 378196
rect 124916 378156 124922 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 58986 377408 58992 377460
rect 59044 377448 59050 377460
rect 59170 377448 59176 377460
rect 59044 377420 59176 377448
rect 59044 377408 59050 377420
rect 59170 377408 59176 377420
rect 59228 377448 59234 377460
rect 67634 377448 67640 377460
rect 59228 377420 67640 377448
rect 59228 377408 59234 377420
rect 67634 377408 67640 377420
rect 67692 377408 67698 377460
rect 118602 377408 118608 377460
rect 118660 377448 118666 377460
rect 121454 377448 121460 377460
rect 118660 377420 121460 377448
rect 118660 377408 118666 377420
rect 121454 377408 121460 377420
rect 121512 377448 121518 377460
rect 146478 377448 146484 377460
rect 121512 377420 146484 377448
rect 121512 377408 121518 377420
rect 146478 377408 146484 377420
rect 146536 377408 146542 377460
rect 66070 376660 66076 376712
rect 66128 376700 66134 376712
rect 68370 376700 68376 376712
rect 66128 376672 68376 376700
rect 66128 376660 66134 376672
rect 68370 376660 68376 376672
rect 68428 376660 68434 376712
rect 118602 376048 118608 376100
rect 118660 376088 118666 376100
rect 128446 376088 128452 376100
rect 118660 376060 128452 376088
rect 118660 376048 118666 376060
rect 128446 376048 128452 376060
rect 128504 376048 128510 376100
rect 49510 375980 49516 376032
rect 49568 376020 49574 376032
rect 59170 376020 59176 376032
rect 49568 375992 59176 376020
rect 49568 375980 49574 375992
rect 59170 375980 59176 375992
rect 59228 375980 59234 376032
rect 118510 375980 118516 376032
rect 118568 376020 118574 376032
rect 120166 376020 120172 376032
rect 118568 375992 120172 376020
rect 118568 375980 118574 375992
rect 120166 375980 120172 375992
rect 120224 376020 120230 376032
rect 143534 376020 143540 376032
rect 120224 375992 143540 376020
rect 120224 375980 120230 375992
rect 143534 375980 143540 375992
rect 143592 375980 143598 376032
rect 64690 375300 64696 375352
rect 64748 375340 64754 375352
rect 66898 375340 66904 375352
rect 64748 375312 66904 375340
rect 64748 375300 64754 375312
rect 66898 375300 66904 375312
rect 66956 375340 66962 375352
rect 67634 375340 67640 375352
rect 66956 375312 67640 375340
rect 66956 375300 66962 375312
rect 67634 375300 67640 375312
rect 67692 375300 67698 375352
rect 118602 375300 118608 375352
rect 118660 375340 118666 375352
rect 151906 375340 151912 375352
rect 118660 375312 151912 375340
rect 118660 375300 118666 375312
rect 151906 375300 151912 375312
rect 151964 375340 151970 375352
rect 153102 375340 153108 375352
rect 151964 375312 153108 375340
rect 151964 375300 151970 375312
rect 153102 375300 153108 375312
rect 153160 375300 153166 375352
rect 153102 374620 153108 374672
rect 153160 374660 153166 374672
rect 202138 374660 202144 374672
rect 153160 374632 202144 374660
rect 153160 374620 153166 374632
rect 202138 374620 202144 374632
rect 202196 374620 202202 374672
rect 67726 374048 67732 374060
rect 67606 374020 67732 374048
rect 42518 373940 42524 373992
rect 42576 373980 42582 373992
rect 66898 373980 66904 373992
rect 42576 373952 66904 373980
rect 42576 373940 42582 373952
rect 66898 373940 66904 373952
rect 66956 373980 66962 373992
rect 67606 373980 67634 374020
rect 67726 374008 67732 374020
rect 67784 374008 67790 374060
rect 66956 373952 67634 373980
rect 66956 373940 66962 373952
rect 117498 373328 117504 373380
rect 117556 373368 117562 373380
rect 123846 373368 123852 373380
rect 117556 373340 123852 373368
rect 117556 373328 117562 373340
rect 123846 373328 123852 373340
rect 123904 373328 123910 373380
rect 118418 372580 118424 372632
rect 118476 372620 118482 372632
rect 222930 372620 222936 372632
rect 118476 372592 222936 372620
rect 118476 372580 118482 372592
rect 222930 372580 222936 372592
rect 222988 372580 222994 372632
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 49050 372552 49056 372564
rect 3292 372524 49056 372552
rect 3292 372512 3298 372524
rect 49050 372512 49056 372524
rect 49108 372512 49114 372564
rect 64782 372512 64788 372564
rect 64840 372552 64846 372564
rect 67634 372552 67640 372564
rect 64840 372524 67640 372552
rect 64840 372512 64846 372524
rect 67634 372512 67640 372524
rect 67692 372512 67698 372564
rect 119982 371900 119988 371952
rect 120040 371940 120046 371952
rect 122926 371940 122932 371952
rect 120040 371912 122932 371940
rect 120040 371900 120046 371912
rect 122926 371900 122932 371912
rect 122984 371900 122990 371952
rect 63218 371220 63224 371272
rect 63276 371260 63282 371272
rect 67450 371260 67456 371272
rect 63276 371232 67456 371260
rect 63276 371220 63282 371232
rect 67450 371220 67456 371232
rect 67508 371260 67514 371272
rect 67634 371260 67640 371272
rect 67508 371232 67640 371260
rect 67508 371220 67514 371232
rect 67634 371220 67640 371232
rect 67692 371220 67698 371272
rect 118602 371220 118608 371272
rect 118660 371260 118666 371272
rect 273990 371260 273996 371272
rect 118660 371232 273996 371260
rect 118660 371220 118666 371232
rect 273990 371220 273996 371232
rect 274048 371220 274054 371272
rect 56226 369792 56232 369844
rect 56284 369832 56290 369844
rect 67634 369832 67640 369844
rect 56284 369804 67640 369832
rect 56284 369792 56290 369804
rect 67634 369792 67640 369804
rect 67692 369792 67698 369844
rect 66162 369112 66168 369164
rect 66220 369152 66226 369164
rect 67726 369152 67732 369164
rect 66220 369124 67732 369152
rect 66220 369112 66226 369124
rect 67726 369112 67732 369124
rect 67784 369112 67790 369164
rect 118970 368500 118976 368552
rect 119028 368540 119034 368552
rect 127066 368540 127072 368552
rect 119028 368512 127072 368540
rect 119028 368500 119034 368512
rect 127066 368500 127072 368512
rect 127124 368500 127130 368552
rect 131666 368432 131672 368484
rect 131724 368472 131730 368484
rect 132494 368472 132500 368484
rect 131724 368444 132500 368472
rect 131724 368432 131730 368444
rect 132494 368432 132500 368444
rect 132552 368432 132558 368484
rect 51994 367752 52000 367804
rect 52052 367792 52058 367804
rect 61470 367792 61476 367804
rect 52052 367764 61476 367792
rect 52052 367752 52058 367764
rect 61470 367752 61476 367764
rect 61528 367752 61534 367804
rect 119338 367752 119344 367804
rect 119396 367792 119402 367804
rect 128354 367792 128360 367804
rect 119396 367764 128360 367792
rect 119396 367752 119402 367764
rect 128354 367752 128360 367764
rect 128412 367752 128418 367804
rect 118602 367208 118608 367260
rect 118660 367248 118666 367260
rect 119338 367248 119344 367260
rect 118660 367220 119344 367248
rect 118660 367208 118666 367220
rect 119338 367208 119344 367220
rect 119396 367208 119402 367260
rect 37182 367072 37188 367124
rect 37240 367112 37246 367124
rect 37240 367084 60412 367112
rect 37240 367072 37246 367084
rect 60384 367044 60412 367084
rect 60458 367072 60464 367124
rect 60516 367112 60522 367124
rect 63402 367112 63408 367124
rect 60516 367084 63408 367112
rect 60516 367072 60522 367084
rect 63402 367072 63408 367084
rect 63460 367112 63466 367124
rect 67634 367112 67640 367124
rect 63460 367084 67640 367112
rect 63460 367072 63466 367084
rect 67634 367072 67640 367084
rect 67692 367072 67698 367124
rect 118510 367072 118516 367124
rect 118568 367112 118574 367124
rect 131666 367112 131672 367124
rect 118568 367084 131672 367112
rect 118568 367072 118574 367084
rect 131666 367072 131672 367084
rect 131724 367072 131730 367124
rect 61378 367044 61384 367056
rect 60384 367016 61384 367044
rect 61378 367004 61384 367016
rect 61436 367044 61442 367056
rect 67726 367044 67732 367056
rect 61436 367016 67732 367044
rect 61436 367004 61442 367016
rect 67726 367004 67732 367016
rect 67784 367004 67790 367056
rect 118602 367004 118608 367056
rect 118660 367044 118666 367056
rect 131114 367044 131120 367056
rect 118660 367016 131120 367044
rect 118660 367004 118666 367016
rect 131114 367004 131120 367016
rect 131172 367004 131178 367056
rect 116026 366936 116032 366988
rect 116084 366976 116090 366988
rect 122926 366976 122932 366988
rect 116084 366948 122932 366976
rect 116084 366936 116090 366948
rect 122926 366936 122932 366948
rect 122984 366936 122990 366988
rect 61470 366324 61476 366376
rect 61528 366364 61534 366376
rect 67634 366364 67640 366376
rect 61528 366336 67640 366364
rect 61528 366324 61534 366336
rect 67634 366324 67640 366336
rect 67692 366324 67698 366376
rect 131114 365712 131120 365764
rect 131172 365752 131178 365764
rect 132494 365752 132500 365764
rect 131172 365724 132500 365752
rect 131172 365712 131178 365724
rect 132494 365712 132500 365724
rect 132552 365712 132558 365764
rect 118694 365100 118700 365152
rect 118752 365140 118758 365152
rect 140866 365140 140872 365152
rect 118752 365112 140872 365140
rect 118752 365100 118758 365112
rect 140866 365100 140872 365112
rect 140924 365100 140930 365152
rect 121546 365032 121552 365084
rect 121604 365072 121610 365084
rect 147766 365072 147772 365084
rect 121604 365044 147772 365072
rect 121604 365032 121610 365044
rect 147766 365032 147772 365044
rect 147824 365032 147830 365084
rect 122926 364964 122932 365016
rect 122984 365004 122990 365016
rect 580258 365004 580264 365016
rect 122984 364976 580264 365004
rect 122984 364964 122990 364976
rect 580258 364964 580264 364976
rect 580316 364964 580322 365016
rect 118602 364760 118608 364812
rect 118660 364800 118666 364812
rect 121546 364800 121552 364812
rect 118660 364772 121552 364800
rect 118660 364760 118666 364772
rect 121546 364760 121552 364772
rect 121604 364760 121610 364812
rect 50798 363672 50804 363724
rect 50856 363712 50862 363724
rect 67634 363712 67640 363724
rect 50856 363684 67640 363712
rect 50856 363672 50862 363684
rect 67634 363672 67640 363684
rect 67692 363672 67698 363724
rect 36906 363604 36912 363656
rect 36964 363644 36970 363656
rect 67726 363644 67732 363656
rect 36964 363616 67732 363644
rect 36964 363604 36970 363616
rect 67726 363604 67732 363616
rect 67784 363604 67790 363656
rect 36906 362924 36912 362976
rect 36964 362964 36970 362976
rect 37090 362964 37096 362976
rect 36964 362936 37096 362964
rect 36964 362924 36970 362936
rect 37090 362924 37096 362936
rect 37148 362924 37154 362976
rect 50614 362924 50620 362976
rect 50672 362964 50678 362976
rect 50798 362964 50804 362976
rect 50672 362936 50804 362964
rect 50672 362924 50678 362936
rect 50798 362924 50804 362936
rect 50856 362924 50862 362976
rect 117958 362856 117964 362908
rect 118016 362896 118022 362908
rect 151814 362896 151820 362908
rect 118016 362868 151820 362896
rect 118016 362856 118022 362868
rect 151814 362856 151820 362868
rect 151872 362896 151878 362908
rect 153102 362896 153108 362908
rect 151872 362868 153108 362896
rect 151872 362856 151878 362868
rect 153102 362856 153108 362868
rect 153160 362856 153166 362908
rect 34146 362176 34152 362228
rect 34204 362216 34210 362228
rect 60734 362216 60740 362228
rect 34204 362188 60740 362216
rect 34204 362176 34210 362188
rect 60734 362176 60740 362188
rect 60792 362176 60798 362228
rect 118602 362176 118608 362228
rect 118660 362216 118666 362228
rect 122098 362216 122104 362228
rect 118660 362188 122104 362216
rect 118660 362176 118666 362188
rect 122098 362176 122104 362188
rect 122156 362216 122162 362228
rect 139486 362216 139492 362228
rect 122156 362188 139492 362216
rect 122156 362176 122162 362188
rect 139486 362176 139492 362188
rect 139544 362176 139550 362228
rect 60734 361632 60740 361684
rect 60792 361672 60798 361684
rect 61746 361672 61752 361684
rect 60792 361644 61752 361672
rect 60792 361632 60798 361644
rect 61746 361632 61752 361644
rect 61804 361672 61810 361684
rect 67634 361672 67640 361684
rect 61804 361644 67640 361672
rect 61804 361632 61810 361644
rect 67634 361632 67640 361644
rect 67692 361632 67698 361684
rect 43806 361564 43812 361616
rect 43864 361604 43870 361616
rect 69198 361604 69204 361616
rect 43864 361576 69204 361604
rect 43864 361564 43870 361576
rect 69198 361564 69204 361576
rect 69256 361564 69262 361616
rect 43898 360816 43904 360868
rect 43956 360856 43962 360868
rect 59170 360856 59176 360868
rect 43956 360828 59176 360856
rect 43956 360816 43962 360828
rect 59170 360816 59176 360828
rect 59228 360816 59234 360868
rect 116670 360272 116676 360324
rect 116728 360312 116734 360324
rect 117222 360312 117228 360324
rect 116728 360284 117228 360312
rect 116728 360272 116734 360284
rect 117222 360272 117228 360284
rect 117280 360312 117286 360324
rect 117280 360284 122834 360312
rect 117280 360272 117286 360284
rect 65610 360244 65616 360256
rect 64846 360216 65616 360244
rect 45462 360136 45468 360188
rect 45520 360176 45526 360188
rect 64846 360176 64874 360216
rect 65610 360204 65616 360216
rect 65668 360244 65674 360256
rect 67634 360244 67640 360256
rect 65668 360216 67640 360244
rect 65668 360204 65674 360216
rect 67634 360204 67640 360216
rect 67692 360204 67698 360256
rect 118602 360204 118608 360256
rect 118660 360244 118666 360256
rect 120166 360244 120172 360256
rect 118660 360216 120172 360244
rect 118660 360204 118666 360216
rect 120166 360204 120172 360216
rect 120224 360204 120230 360256
rect 122806 360244 122834 360284
rect 132678 360244 132684 360256
rect 122806 360216 132684 360244
rect 132678 360204 132684 360216
rect 132736 360204 132742 360256
rect 45520 360148 64874 360176
rect 45520 360136 45526 360148
rect 118142 360136 118148 360188
rect 118200 360176 118206 360188
rect 147674 360176 147680 360188
rect 118200 360148 147680 360176
rect 118200 360136 118206 360148
rect 147674 360136 147680 360148
rect 147732 360136 147738 360188
rect 120166 360068 120172 360120
rect 120224 360108 120230 360120
rect 120718 360108 120724 360120
rect 120224 360080 120724 360108
rect 120224 360068 120230 360080
rect 120718 360068 120724 360080
rect 120776 360108 120782 360120
rect 129918 360108 129924 360120
rect 120776 360080 129924 360108
rect 120776 360068 120782 360080
rect 129918 360068 129924 360080
rect 129976 360068 129982 360120
rect 61470 359524 61476 359576
rect 61528 359564 61534 359576
rect 61838 359564 61844 359576
rect 61528 359536 61844 359564
rect 61528 359524 61534 359536
rect 61838 359524 61844 359536
rect 61896 359524 61902 359576
rect 59170 359456 59176 359508
rect 59228 359496 59234 359508
rect 67634 359496 67640 359508
rect 59228 359468 67640 359496
rect 59228 359456 59234 359468
rect 67634 359456 67640 359468
rect 67692 359456 67698 359508
rect 147674 359456 147680 359508
rect 147732 359496 147738 359508
rect 197998 359496 198004 359508
rect 147732 359468 198004 359496
rect 147732 359456 147738 359468
rect 197998 359456 198004 359468
rect 198056 359456 198062 359508
rect 118602 358436 118608 358488
rect 118660 358476 118666 358488
rect 124214 358476 124220 358488
rect 118660 358448 124220 358476
rect 118660 358436 118666 358448
rect 124214 358436 124220 358448
rect 124272 358436 124278 358488
rect 54846 358028 54852 358080
rect 54904 358068 54910 358080
rect 55122 358068 55128 358080
rect 54904 358040 55128 358068
rect 54904 358028 54910 358040
rect 55122 358028 55128 358040
rect 55180 358068 55186 358080
rect 67634 358068 67640 358080
rect 55180 358040 67640 358068
rect 55180 358028 55186 358040
rect 67634 358028 67640 358040
rect 67692 358028 67698 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 22738 357456 22744 357468
rect 3200 357428 22744 357456
rect 3200 357416 3206 357428
rect 22738 357416 22744 357428
rect 22796 357416 22802 357468
rect 62850 357456 62856 357468
rect 62132 357428 62856 357456
rect 40678 357348 40684 357400
rect 40736 357388 40742 357400
rect 62132 357388 62160 357428
rect 62850 357416 62856 357428
rect 62908 357456 62914 357468
rect 67726 357456 67732 357468
rect 62908 357428 67732 357456
rect 62908 357416 62914 357428
rect 67726 357416 67732 357428
rect 67784 357416 67790 357468
rect 40736 357360 62160 357388
rect 40736 357348 40742 357360
rect 115290 357348 115296 357400
rect 115348 357388 115354 357400
rect 117314 357388 117320 357400
rect 115348 357360 117320 357388
rect 115348 357348 115354 357360
rect 117314 357348 117320 357360
rect 117372 357348 117378 357400
rect 117682 357008 117688 357060
rect 117740 357048 117746 357060
rect 121638 357048 121644 357060
rect 117740 357020 121644 357048
rect 117740 357008 117746 357020
rect 121638 357008 121644 357020
rect 121696 357008 121702 357060
rect 122190 356736 122196 356788
rect 122248 356776 122254 356788
rect 128354 356776 128360 356788
rect 122248 356748 128360 356776
rect 122248 356736 122254 356748
rect 128354 356736 128360 356748
rect 128412 356736 128418 356788
rect 50890 356668 50896 356720
rect 50948 356708 50954 356720
rect 60642 356708 60648 356720
rect 50948 356680 60648 356708
rect 50948 356668 50954 356680
rect 60642 356668 60648 356680
rect 60700 356668 60706 356720
rect 124950 356668 124956 356720
rect 125008 356708 125014 356720
rect 325694 356708 325700 356720
rect 125008 356680 325700 356708
rect 125008 356668 125014 356680
rect 325694 356668 325700 356680
rect 325752 356668 325758 356720
rect 60642 356124 60648 356176
rect 60700 356164 60706 356176
rect 67726 356164 67732 356176
rect 60700 356136 67732 356164
rect 60700 356124 60706 356136
rect 67726 356124 67732 356136
rect 67784 356124 67790 356176
rect 34146 356056 34152 356108
rect 34204 356096 34210 356108
rect 69474 356096 69480 356108
rect 34204 356068 69480 356096
rect 34204 356056 34210 356068
rect 69474 356056 69480 356068
rect 69532 356056 69538 356108
rect 118602 355988 118608 356040
rect 118660 356028 118666 356040
rect 142246 356028 142252 356040
rect 118660 356000 142252 356028
rect 118660 355988 118666 356000
rect 142246 355988 142252 356000
rect 142304 356028 142310 356040
rect 143442 356028 143448 356040
rect 142304 356000 143448 356028
rect 142304 355988 142310 356000
rect 143442 355988 143448 356000
rect 143500 355988 143506 356040
rect 63494 355308 63500 355360
rect 63552 355348 63558 355360
rect 67634 355348 67640 355360
rect 63552 355320 67640 355348
rect 63552 355308 63558 355320
rect 67634 355308 67640 355320
rect 67692 355308 67698 355360
rect 143442 355308 143448 355360
rect 143500 355348 143506 355360
rect 233878 355348 233884 355360
rect 143500 355320 233884 355348
rect 143500 355308 143506 355320
rect 233878 355308 233884 355320
rect 233936 355308 233942 355360
rect 118602 354628 118608 354680
rect 118660 354668 118666 354680
rect 133966 354668 133972 354680
rect 118660 354640 133972 354668
rect 118660 354628 118666 354640
rect 133966 354628 133972 354640
rect 134024 354628 134030 354680
rect 121638 353948 121644 354000
rect 121696 353988 121702 354000
rect 324406 353988 324412 354000
rect 121696 353960 324412 353988
rect 121696 353948 121702 353960
rect 324406 353948 324412 353960
rect 324464 353948 324470 354000
rect 133966 353336 133972 353388
rect 134024 353376 134030 353388
rect 138014 353376 138020 353388
rect 134024 353348 138020 353376
rect 134024 353336 134030 353348
rect 138014 353336 138020 353348
rect 138072 353336 138078 353388
rect 67634 353308 67640 353320
rect 67376 353280 67640 353308
rect 56410 353200 56416 353252
rect 56468 353240 56474 353252
rect 66990 353240 66996 353252
rect 56468 353212 66996 353240
rect 56468 353200 56474 353212
rect 66990 353200 66996 353212
rect 67048 353240 67054 353252
rect 67376 353240 67404 353280
rect 67634 353268 67640 353280
rect 67692 353268 67698 353320
rect 118050 353268 118056 353320
rect 118108 353308 118114 353320
rect 133874 353308 133880 353320
rect 118108 353280 133880 353308
rect 118108 353268 118114 353280
rect 133874 353268 133880 353280
rect 133932 353308 133938 353320
rect 136818 353308 136824 353320
rect 133932 353280 136824 353308
rect 133932 353268 133938 353280
rect 136818 353268 136824 353280
rect 136876 353268 136882 353320
rect 67048 353212 67404 353240
rect 67048 353200 67054 353212
rect 11698 352520 11704 352572
rect 11756 352560 11762 352572
rect 34238 352560 34244 352572
rect 11756 352532 34244 352560
rect 11756 352520 11762 352532
rect 34238 352520 34244 352532
rect 34296 352560 34302 352572
rect 41414 352560 41420 352572
rect 34296 352532 41420 352560
rect 34296 352520 34302 352532
rect 41414 352520 41420 352532
rect 41472 352520 41478 352572
rect 62758 352520 62764 352572
rect 62816 352560 62822 352572
rect 67910 352560 67916 352572
rect 62816 352532 67916 352560
rect 62816 352520 62822 352532
rect 67910 352520 67916 352532
rect 67968 352520 67974 352572
rect 41414 351908 41420 351960
rect 41472 351948 41478 351960
rect 42702 351948 42708 351960
rect 41472 351920 42708 351948
rect 41472 351908 41478 351920
rect 42702 351908 42708 351920
rect 42760 351948 42766 351960
rect 67634 351948 67640 351960
rect 42760 351920 67640 351948
rect 42760 351908 42766 351920
rect 67634 351908 67640 351920
rect 67692 351908 67698 351960
rect 116578 351296 116584 351348
rect 116636 351336 116642 351348
rect 128446 351336 128452 351348
rect 116636 351308 128452 351336
rect 116636 351296 116642 351308
rect 128446 351296 128452 351308
rect 128504 351296 128510 351348
rect 118418 351228 118424 351280
rect 118476 351268 118482 351280
rect 204898 351268 204904 351280
rect 118476 351240 204904 351268
rect 118476 351228 118482 351240
rect 204898 351228 204904 351240
rect 204956 351228 204962 351280
rect 64598 351160 64604 351212
rect 64656 351200 64662 351212
rect 67726 351200 67732 351212
rect 64656 351172 67732 351200
rect 64656 351160 64662 351172
rect 67726 351160 67732 351172
rect 67784 351160 67790 351212
rect 118510 351160 118516 351212
rect 118568 351200 118574 351212
rect 271230 351200 271236 351212
rect 118568 351172 271236 351200
rect 118568 351160 118574 351172
rect 271230 351160 271236 351172
rect 271288 351160 271294 351212
rect 118602 349868 118608 349920
rect 118660 349908 118666 349920
rect 124398 349908 124404 349920
rect 118660 349880 124404 349908
rect 118660 349868 118666 349880
rect 124398 349868 124404 349880
rect 124456 349908 124462 349920
rect 126974 349908 126980 349920
rect 124456 349880 126980 349908
rect 124456 349868 124462 349880
rect 126974 349868 126980 349880
rect 127032 349868 127038 349920
rect 63310 349800 63316 349852
rect 63368 349840 63374 349852
rect 68002 349840 68008 349852
rect 63368 349812 68008 349840
rect 63368 349800 63374 349812
rect 68002 349800 68008 349812
rect 68060 349800 68066 349852
rect 126238 349800 126244 349852
rect 126296 349840 126302 349852
rect 314654 349840 314660 349852
rect 126296 349812 314660 349840
rect 126296 349800 126302 349812
rect 314654 349800 314660 349812
rect 314712 349800 314718 349852
rect 42058 349120 42064 349172
rect 42116 349160 42122 349172
rect 45462 349160 45468 349172
rect 42116 349132 45468 349160
rect 42116 349120 42122 349132
rect 45462 349120 45468 349132
rect 45520 349160 45526 349172
rect 67634 349160 67640 349172
rect 45520 349132 67640 349160
rect 45520 349120 45526 349132
rect 67634 349120 67640 349132
rect 67692 349120 67698 349172
rect 61930 348372 61936 348424
rect 61988 348412 61994 348424
rect 68830 348412 68836 348424
rect 61988 348384 68836 348412
rect 61988 348372 61994 348384
rect 68830 348372 68836 348384
rect 68888 348372 68894 348424
rect 118602 347828 118608 347880
rect 118660 347868 118666 347880
rect 140866 347868 140872 347880
rect 118660 347840 140872 347868
rect 118660 347828 118666 347840
rect 140866 347828 140872 347840
rect 140924 347828 140930 347880
rect 117774 347760 117780 347812
rect 117832 347800 117838 347812
rect 258718 347800 258724 347812
rect 117832 347772 258724 347800
rect 117832 347760 117838 347772
rect 258718 347760 258724 347772
rect 258776 347760 258782 347812
rect 117406 347692 117412 347744
rect 117464 347732 117470 347744
rect 133782 347732 133788 347744
rect 117464 347704 133788 347732
rect 117464 347692 117470 347704
rect 133782 347692 133788 347704
rect 133840 347692 133846 347744
rect 140866 347692 140872 347744
rect 140924 347732 140930 347744
rect 149238 347732 149244 347744
rect 140924 347704 149244 347732
rect 140924 347692 140930 347704
rect 149238 347692 149244 347704
rect 149296 347692 149302 347744
rect 133782 347080 133788 347132
rect 133840 347120 133846 347132
rect 191098 347120 191104 347132
rect 133840 347092 191104 347120
rect 133840 347080 133846 347092
rect 191098 347080 191104 347092
rect 191156 347080 191162 347132
rect 3326 347012 3332 347064
rect 3384 347052 3390 347064
rect 25498 347052 25504 347064
rect 3384 347024 25504 347052
rect 3384 347012 3390 347024
rect 25498 347012 25504 347024
rect 25556 347012 25562 347064
rect 64506 347012 64512 347064
rect 64564 347052 64570 347064
rect 68554 347052 68560 347064
rect 64564 347024 68560 347052
rect 64564 347012 64570 347024
rect 68554 347012 68560 347024
rect 68612 347012 68618 347064
rect 149238 347012 149244 347064
rect 149296 347052 149302 347064
rect 316126 347052 316132 347064
rect 149296 347024 316132 347052
rect 149296 347012 149302 347024
rect 316126 347012 316132 347024
rect 316184 347012 316190 347064
rect 65518 346400 65524 346452
rect 65576 346440 65582 346452
rect 67634 346440 67640 346452
rect 65576 346412 67640 346440
rect 65576 346400 65582 346412
rect 67634 346400 67640 346412
rect 67692 346400 67698 346452
rect 22738 346332 22744 346384
rect 22796 346372 22802 346384
rect 35710 346372 35716 346384
rect 22796 346344 35716 346372
rect 22796 346332 22802 346344
rect 35710 346332 35716 346344
rect 35768 346332 35774 346384
rect 118602 346332 118608 346384
rect 118660 346372 118666 346384
rect 146386 346372 146392 346384
rect 118660 346344 146392 346372
rect 118660 346332 118666 346344
rect 146386 346332 146392 346344
rect 146444 346372 146450 346384
rect 146754 346372 146760 346384
rect 146444 346344 146760 346372
rect 146444 346332 146450 346344
rect 146754 346332 146760 346344
rect 146812 346332 146818 346384
rect 35710 345652 35716 345704
rect 35768 345692 35774 345704
rect 63310 345692 63316 345704
rect 35768 345664 63316 345692
rect 35768 345652 35774 345664
rect 63310 345652 63316 345664
rect 63368 345652 63374 345704
rect 118326 345652 118332 345704
rect 118384 345692 118390 345704
rect 122926 345692 122932 345704
rect 118384 345664 122932 345692
rect 118384 345652 118390 345664
rect 122926 345652 122932 345664
rect 122984 345692 122990 345704
rect 131298 345692 131304 345704
rect 122984 345664 131304 345692
rect 122984 345652 122990 345664
rect 131298 345652 131304 345664
rect 131356 345652 131362 345704
rect 146754 345652 146760 345704
rect 146812 345692 146818 345704
rect 217226 345692 217232 345704
rect 146812 345664 217232 345692
rect 146812 345652 146818 345664
rect 217226 345652 217232 345664
rect 217284 345652 217290 345704
rect 63310 345040 63316 345092
rect 63368 345080 63374 345092
rect 67726 345080 67732 345092
rect 63368 345052 67732 345080
rect 63368 345040 63374 345052
rect 67726 345040 67732 345052
rect 67784 345040 67790 345092
rect 116670 345040 116676 345092
rect 116728 345080 116734 345092
rect 124306 345080 124312 345092
rect 116728 345052 124312 345080
rect 116728 345040 116734 345052
rect 124306 345040 124312 345052
rect 124364 345040 124370 345092
rect 66070 344972 66076 345024
rect 66128 345012 66134 345024
rect 67634 345012 67640 345024
rect 66128 344984 67640 345012
rect 66128 344972 66134 344984
rect 67634 344972 67640 344984
rect 67692 344972 67698 345024
rect 118602 344972 118608 345024
rect 118660 345012 118666 345024
rect 149054 345012 149060 345024
rect 118660 344984 149060 345012
rect 118660 344972 118666 344984
rect 149054 344972 149060 344984
rect 149112 344972 149118 345024
rect 149054 344292 149060 344344
rect 149112 344332 149118 344344
rect 331858 344332 331864 344344
rect 149112 344304 331864 344332
rect 149112 344292 149118 344304
rect 331858 344292 331864 344304
rect 331916 344292 331922 344344
rect 63494 343680 63500 343732
rect 63552 343720 63558 343732
rect 67726 343720 67732 343732
rect 63552 343692 67732 343720
rect 63552 343680 63558 343692
rect 67726 343680 67732 343692
rect 67784 343680 67790 343732
rect 45186 343612 45192 343664
rect 45244 343652 45250 343664
rect 47854 343652 47860 343664
rect 45244 343624 47860 343652
rect 45244 343612 45250 343624
rect 47854 343612 47860 343624
rect 47912 343652 47918 343664
rect 67634 343652 67640 343664
rect 47912 343624 67640 343652
rect 47912 343612 47918 343624
rect 67634 343612 67640 343624
rect 67692 343612 67698 343664
rect 118602 343544 118608 343596
rect 118660 343584 118666 343596
rect 150434 343584 150440 343596
rect 118660 343556 150440 343584
rect 118660 343544 118666 343556
rect 150434 343544 150440 343556
rect 150492 343544 150498 343596
rect 128722 342932 128728 342984
rect 128780 342972 128786 342984
rect 129826 342972 129832 342984
rect 128780 342944 129832 342972
rect 128780 342932 128786 342944
rect 129826 342932 129832 342944
rect 129884 342932 129890 342984
rect 36998 342864 37004 342916
rect 37056 342904 37062 342916
rect 41138 342904 41144 342916
rect 37056 342876 41144 342904
rect 37056 342864 37062 342876
rect 41138 342864 41144 342876
rect 41196 342904 41202 342916
rect 63494 342904 63500 342916
rect 41196 342876 63500 342904
rect 41196 342864 41202 342876
rect 63494 342864 63500 342876
rect 63552 342864 63558 342916
rect 150434 342864 150440 342916
rect 150492 342904 150498 342916
rect 282178 342904 282184 342916
rect 150492 342876 282184 342904
rect 150492 342864 150498 342876
rect 282178 342864 282184 342876
rect 282236 342864 282242 342916
rect 115290 342320 115296 342372
rect 115348 342360 115354 342372
rect 118786 342360 118792 342372
rect 115348 342332 118792 342360
rect 115348 342320 115354 342332
rect 118786 342320 118792 342332
rect 118844 342320 118850 342372
rect 118142 342252 118148 342304
rect 118200 342292 118206 342304
rect 128722 342292 128728 342304
rect 118200 342264 128728 342292
rect 118200 342252 118206 342264
rect 128722 342252 128728 342264
rect 128780 342252 128786 342304
rect 118602 341504 118608 341556
rect 118660 341544 118666 341556
rect 142338 341544 142344 341556
rect 118660 341516 142344 341544
rect 118660 341504 118666 341516
rect 142338 341504 142344 341516
rect 142396 341504 142402 341556
rect 65978 340932 65984 340944
rect 64846 340904 65984 340932
rect 38562 340824 38568 340876
rect 38620 340864 38626 340876
rect 64846 340864 64874 340904
rect 65978 340892 65984 340904
rect 66036 340932 66042 340944
rect 67634 340932 67640 340944
rect 66036 340904 67640 340932
rect 66036 340892 66042 340904
rect 67634 340892 67640 340904
rect 67692 340892 67698 340944
rect 118786 340932 118792 340944
rect 118699 340904 118792 340932
rect 38620 340836 64874 340864
rect 38620 340824 38626 340836
rect 118050 340824 118056 340876
rect 118108 340864 118114 340876
rect 118712 340864 118740 340904
rect 118786 340892 118792 340904
rect 118844 340932 118850 340944
rect 120074 340932 120080 340944
rect 118844 340904 120080 340932
rect 118844 340892 118850 340904
rect 120074 340892 120080 340904
rect 120132 340892 120138 340944
rect 140866 340892 140872 340944
rect 140924 340932 140930 340944
rect 580258 340932 580264 340944
rect 140924 340904 580264 340932
rect 140924 340892 140930 340904
rect 580258 340892 580264 340904
rect 580316 340892 580322 340944
rect 150526 340864 150532 340876
rect 118108 340836 118740 340864
rect 122806 340836 150532 340864
rect 118108 340824 118114 340836
rect 117774 340756 117780 340808
rect 117832 340796 117838 340808
rect 122806 340796 122834 340836
rect 150526 340824 150532 340836
rect 150584 340864 150590 340876
rect 151538 340864 151544 340876
rect 150584 340836 151544 340864
rect 150584 340824 150590 340836
rect 151538 340824 151544 340836
rect 151596 340824 151602 340876
rect 117832 340768 122834 340796
rect 117832 340756 117838 340768
rect 151538 340144 151544 340196
rect 151596 340184 151602 340196
rect 352558 340184 352564 340196
rect 151596 340156 352564 340184
rect 151596 340144 151602 340156
rect 352558 340144 352564 340156
rect 352616 340144 352622 340196
rect 113910 339600 113916 339652
rect 113968 339640 113974 339652
rect 115106 339640 115112 339652
rect 113968 339612 115112 339640
rect 113968 339600 113974 339612
rect 115106 339600 115112 339612
rect 115164 339640 115170 339652
rect 143626 339640 143632 339652
rect 115164 339612 143632 339640
rect 115164 339600 115170 339612
rect 143626 339600 143632 339612
rect 143684 339600 143690 339652
rect 61654 339532 61660 339584
rect 61712 339572 61718 339584
rect 73246 339572 73252 339584
rect 61712 339544 73252 339572
rect 61712 339532 61718 339544
rect 73246 339532 73252 339544
rect 73304 339532 73310 339584
rect 113818 339532 113824 339584
rect 113876 339572 113882 339584
rect 140774 339572 140780 339584
rect 113876 339544 140780 339572
rect 113876 339532 113882 339544
rect 140774 339532 140780 339544
rect 140832 339532 140838 339584
rect 48038 339464 48044 339516
rect 48096 339504 48102 339516
rect 71958 339504 71964 339516
rect 48096 339476 71964 339504
rect 48096 339464 48102 339476
rect 71958 339464 71964 339476
rect 72016 339464 72022 339516
rect 48958 339396 48964 339448
rect 49016 339436 49022 339448
rect 76650 339436 76656 339448
rect 49016 339408 76656 339436
rect 49016 339396 49022 339408
rect 76650 339396 76656 339408
rect 76708 339436 76714 339448
rect 77110 339436 77116 339448
rect 76708 339408 77116 339436
rect 76708 339396 76714 339408
rect 77110 339396 77116 339408
rect 77168 339396 77174 339448
rect 87414 339396 87420 339448
rect 87472 339436 87478 339448
rect 87598 339436 87604 339448
rect 87472 339408 87604 339436
rect 87472 339396 87478 339408
rect 87598 339396 87604 339408
rect 87656 339436 87662 339448
rect 580350 339436 580356 339448
rect 87656 339408 580356 339436
rect 87656 339396 87662 339408
rect 580350 339396 580356 339408
rect 580408 339396 580414 339448
rect 56318 339328 56324 339380
rect 56376 339368 56382 339380
rect 73890 339368 73896 339380
rect 56376 339340 73896 339368
rect 56376 339328 56382 339340
rect 73890 339328 73896 339340
rect 73948 339368 73954 339380
rect 74442 339368 74448 339380
rect 73948 339340 74448 339368
rect 73948 339328 73954 339340
rect 74442 339328 74448 339340
rect 74500 339368 74506 339380
rect 124858 339368 124864 339380
rect 74500 339340 124864 339368
rect 74500 339328 74506 339340
rect 124858 339328 124864 339340
rect 124916 339328 124922 339380
rect 58894 339260 58900 339312
rect 58952 339300 58958 339312
rect 93210 339300 93216 339312
rect 58952 339272 93216 339300
rect 58952 339260 58958 339272
rect 93210 339260 93216 339272
rect 93268 339260 93274 339312
rect 113174 339260 113180 339312
rect 113232 339300 113238 339312
rect 114002 339300 114008 339312
rect 113232 339272 114008 339300
rect 113232 339260 113238 339272
rect 114002 339260 114008 339272
rect 114060 339300 114066 339312
rect 144914 339300 144920 339312
rect 114060 339272 144920 339300
rect 114060 339260 114066 339272
rect 144914 339260 144920 339272
rect 144972 339260 144978 339312
rect 54938 339192 54944 339244
rect 54996 339232 55002 339244
rect 57238 339232 57244 339244
rect 54996 339204 57244 339232
rect 54996 339192 55002 339204
rect 57238 339192 57244 339204
rect 57296 339232 57302 339244
rect 82262 339232 82268 339244
rect 57296 339204 82268 339232
rect 57296 339192 57302 339204
rect 82262 339192 82268 339204
rect 82320 339192 82326 339244
rect 100294 339192 100300 339244
rect 100352 339232 100358 339244
rect 125594 339232 125600 339244
rect 100352 339204 125600 339232
rect 100352 339192 100358 339204
rect 125594 339192 125600 339204
rect 125652 339232 125658 339244
rect 125870 339232 125876 339244
rect 125652 339204 125876 339232
rect 125652 339192 125658 339204
rect 125870 339192 125876 339204
rect 125928 339192 125934 339244
rect 127158 339164 127164 339176
rect 103486 339136 127164 339164
rect 102226 339056 102232 339108
rect 102284 339096 102290 339108
rect 103330 339096 103336 339108
rect 102284 339068 103336 339096
rect 102284 339056 102290 339068
rect 103330 339056 103336 339068
rect 103388 339096 103394 339108
rect 103486 339096 103514 339136
rect 127158 339124 127164 339136
rect 127216 339124 127222 339176
rect 103388 339068 103514 339096
rect 103388 339056 103394 339068
rect 66070 338784 66076 338836
rect 66128 338824 66134 338836
rect 80698 338824 80704 338836
rect 66128 338796 80704 338824
rect 66128 338784 66134 338796
rect 80698 338784 80704 338796
rect 80756 338784 80762 338836
rect 62850 338716 62856 338768
rect 62908 338756 62914 338768
rect 97258 338756 97264 338768
rect 62908 338728 97264 338756
rect 62908 338716 62914 338728
rect 97258 338716 97264 338728
rect 97316 338716 97322 338768
rect 104158 338716 104164 338768
rect 104216 338756 104222 338768
rect 120718 338756 120724 338768
rect 104216 338728 120724 338756
rect 104216 338716 104222 338728
rect 120718 338716 120724 338728
rect 120776 338716 120782 338768
rect 91002 338104 91008 338156
rect 91060 338144 91066 338156
rect 91922 338144 91928 338156
rect 91060 338116 91928 338144
rect 91060 338104 91066 338116
rect 91922 338104 91928 338116
rect 91980 338104 91986 338156
rect 70026 338036 70032 338088
rect 70084 338076 70090 338088
rect 72970 338076 72976 338088
rect 70084 338048 72976 338076
rect 70084 338036 70090 338048
rect 72970 338036 72976 338048
rect 73028 338036 73034 338088
rect 75822 338036 75828 338088
rect 75880 338076 75886 338088
rect 79962 338076 79968 338088
rect 75880 338048 79968 338076
rect 75880 338036 75886 338048
rect 79962 338036 79968 338048
rect 80020 338036 80026 338088
rect 108022 338036 108028 338088
rect 108080 338076 108086 338088
rect 143810 338076 143816 338088
rect 108080 338048 143816 338076
rect 108080 338036 108086 338048
rect 143810 338036 143816 338048
rect 143868 338036 143874 338088
rect 47946 337968 47952 338020
rect 48004 338008 48010 338020
rect 83550 338008 83556 338020
rect 48004 337980 83556 338008
rect 48004 337968 48010 337980
rect 83550 337968 83556 337980
rect 83608 337968 83614 338020
rect 115750 337968 115756 338020
rect 115808 338008 115814 338020
rect 141050 338008 141056 338020
rect 115808 337980 141056 338008
rect 115808 337968 115814 337980
rect 141050 337968 141056 337980
rect 141108 338008 141114 338020
rect 141326 338008 141332 338020
rect 141108 337980 141332 338008
rect 141108 337968 141114 337980
rect 141326 337968 141332 337980
rect 141384 337968 141390 338020
rect 61378 337900 61384 337952
rect 61436 337940 61442 337952
rect 84194 337940 84200 337952
rect 61436 337912 84200 337940
rect 61436 337900 61442 337912
rect 84194 337900 84200 337912
rect 84252 337900 84258 337952
rect 97718 337900 97724 337952
rect 97776 337940 97782 337952
rect 128446 337940 128452 337952
rect 97776 337912 128452 337940
rect 97776 337900 97782 337912
rect 128446 337900 128452 337912
rect 128504 337900 128510 337952
rect 57606 337832 57612 337884
rect 57664 337872 57670 337884
rect 76466 337872 76472 337884
rect 57664 337844 76472 337872
rect 57664 337832 57670 337844
rect 76466 337832 76472 337844
rect 76524 337832 76530 337884
rect 95786 337832 95792 337884
rect 95844 337872 95850 337884
rect 125778 337872 125784 337884
rect 95844 337844 125784 337872
rect 95844 337832 95850 337844
rect 125778 337832 125784 337844
rect 125836 337872 125842 337884
rect 126882 337872 126888 337884
rect 125836 337844 126888 337872
rect 125836 337832 125842 337844
rect 126882 337832 126888 337844
rect 126940 337832 126946 337884
rect 86770 337764 86776 337816
rect 86828 337804 86834 337816
rect 120442 337804 120448 337816
rect 86828 337776 120448 337804
rect 86828 337764 86834 337776
rect 120442 337764 120448 337776
rect 120500 337764 120506 337816
rect 57882 337696 57888 337748
rect 57940 337736 57946 337748
rect 60366 337736 60372 337748
rect 57940 337708 60372 337736
rect 57940 337696 57946 337708
rect 60366 337696 60372 337708
rect 60424 337736 60430 337748
rect 98362 337736 98368 337748
rect 60424 337708 98368 337736
rect 60424 337696 60430 337708
rect 98362 337696 98368 337708
rect 98420 337696 98426 337748
rect 105538 337696 105544 337748
rect 105596 337736 105602 337748
rect 108022 337736 108028 337748
rect 105596 337708 108028 337736
rect 105596 337696 105602 337708
rect 108022 337696 108028 337708
rect 108080 337696 108086 337748
rect 80974 337628 80980 337680
rect 81032 337668 81038 337680
rect 81434 337668 81440 337680
rect 81032 337640 81440 337668
rect 81032 337628 81038 337640
rect 81434 337628 81440 337640
rect 81492 337628 81498 337680
rect 141326 337424 141332 337476
rect 141384 337464 141390 337476
rect 196618 337464 196624 337476
rect 141384 337436 196624 337464
rect 141384 337424 141390 337436
rect 196618 337424 196624 337436
rect 196676 337424 196682 337476
rect 66990 337356 66996 337408
rect 67048 337396 67054 337408
rect 77294 337396 77300 337408
rect 67048 337368 77300 337396
rect 67048 337356 67054 337368
rect 77294 337356 77300 337368
rect 77352 337356 77358 337408
rect 99650 337356 99656 337408
rect 99708 337396 99714 337408
rect 103422 337396 103428 337408
rect 99708 337368 103428 337396
rect 99708 337356 99714 337368
rect 103422 337356 103428 337368
rect 103480 337396 103486 337408
rect 123110 337396 123116 337408
rect 103480 337368 123116 337396
rect 103480 337356 103486 337368
rect 123110 337356 123116 337368
rect 123168 337356 123174 337408
rect 126882 337356 126888 337408
rect 126940 337396 126946 337408
rect 276658 337396 276664 337408
rect 126940 337368 276664 337396
rect 126940 337356 126946 337368
rect 276658 337356 276664 337368
rect 276716 337356 276722 337408
rect 102870 337220 102876 337272
rect 102928 337260 102934 337272
rect 104894 337260 104900 337272
rect 102928 337232 104900 337260
rect 102928 337220 102934 337232
rect 104894 337220 104900 337232
rect 104952 337220 104958 337272
rect 103514 337016 103520 337068
rect 103572 337056 103578 337068
rect 109126 337056 109132 337068
rect 103572 337028 109132 337056
rect 103572 337016 103578 337028
rect 109126 337016 109132 337028
rect 109184 337016 109190 337068
rect 92566 336812 92572 336864
rect 92624 336852 92630 336864
rect 95234 336852 95240 336864
rect 92624 336824 95240 336852
rect 92624 336812 92630 336824
rect 95234 336812 95240 336824
rect 95292 336812 95298 336864
rect 71958 336744 71964 336796
rect 72016 336784 72022 336796
rect 75178 336784 75184 336796
rect 72016 336756 75184 336784
rect 72016 336744 72022 336756
rect 75178 336744 75184 336756
rect 75236 336744 75242 336796
rect 81618 336744 81624 336796
rect 81676 336784 81682 336796
rect 100018 336784 100024 336796
rect 81676 336756 100024 336784
rect 81676 336744 81682 336756
rect 100018 336744 100024 336756
rect 100076 336744 100082 336796
rect 112438 336744 112444 336796
rect 112496 336784 112502 336796
rect 113818 336784 113824 336796
rect 112496 336756 113824 336784
rect 112496 336744 112502 336756
rect 113818 336744 113824 336756
rect 113876 336744 113882 336796
rect 128446 336744 128452 336796
rect 128504 336784 128510 336796
rect 180058 336784 180064 336796
rect 128504 336756 180064 336784
rect 128504 336744 128510 336756
rect 180058 336744 180064 336756
rect 180116 336744 180122 336796
rect 41322 336676 41328 336728
rect 41380 336716 41386 336728
rect 74534 336716 74540 336728
rect 41380 336688 74540 336716
rect 41380 336676 41386 336688
rect 74534 336676 74540 336688
rect 74592 336716 74598 336728
rect 75270 336716 75276 336728
rect 74592 336688 75276 336716
rect 74592 336676 74598 336688
rect 75270 336676 75276 336688
rect 75328 336676 75334 336728
rect 91278 336676 91284 336728
rect 91336 336716 91342 336728
rect 92382 336716 92388 336728
rect 91336 336688 92388 336716
rect 91336 336676 91342 336688
rect 92382 336676 92388 336688
rect 92440 336716 92446 336728
rect 92440 336688 93854 336716
rect 92440 336676 92446 336688
rect 46750 336608 46756 336660
rect 46808 336648 46814 336660
rect 78674 336648 78680 336660
rect 46808 336620 78680 336648
rect 46808 336608 46814 336620
rect 78674 336608 78680 336620
rect 78732 336608 78738 336660
rect 93826 336648 93854 336688
rect 107562 336676 107568 336728
rect 107620 336716 107626 336728
rect 139578 336716 139584 336728
rect 107620 336688 139584 336716
rect 107620 336676 107626 336688
rect 139578 336676 139584 336688
rect 139636 336676 139642 336728
rect 116670 336648 116676 336660
rect 93826 336620 116676 336648
rect 116670 336608 116676 336620
rect 116728 336608 116734 336660
rect 126974 336608 126980 336660
rect 127032 336648 127038 336660
rect 128538 336648 128544 336660
rect 127032 336620 128544 336648
rect 127032 336608 127038 336620
rect 128538 336608 128544 336620
rect 128596 336608 128602 336660
rect 59078 336540 59084 336592
rect 59136 336580 59142 336592
rect 88978 336580 88984 336592
rect 59136 336552 88984 336580
rect 59136 336540 59142 336552
rect 88978 336540 88984 336552
rect 89036 336540 89042 336592
rect 109862 336540 109868 336592
rect 109920 336580 109926 336592
rect 134058 336580 134064 336592
rect 109920 336552 134064 336580
rect 109920 336540 109926 336552
rect 134058 336540 134064 336552
rect 134116 336540 134122 336592
rect 53558 336472 53564 336524
rect 53616 336512 53622 336524
rect 79318 336512 79324 336524
rect 53616 336484 79324 336512
rect 53616 336472 53622 336484
rect 79318 336472 79324 336484
rect 79376 336472 79382 336524
rect 56410 336404 56416 336456
rect 56468 336444 56474 336456
rect 60550 336444 60556 336456
rect 56468 336416 60556 336444
rect 56468 336404 56474 336416
rect 60550 336404 60556 336416
rect 60608 336444 60614 336456
rect 84746 336444 84752 336456
rect 60608 336416 84752 336444
rect 60608 336404 60614 336416
rect 84746 336404 84752 336416
rect 84804 336404 84810 336456
rect 109126 335996 109132 336048
rect 109184 336036 109190 336048
rect 126974 336036 126980 336048
rect 109184 336008 126980 336036
rect 109184 335996 109190 336008
rect 126974 335996 126980 336008
rect 127032 335996 127038 336048
rect 45278 335248 45284 335300
rect 45336 335288 45342 335300
rect 81618 335288 81624 335300
rect 45336 335260 81624 335288
rect 45336 335248 45342 335260
rect 81618 335248 81624 335260
rect 81676 335248 81682 335300
rect 108298 335248 108304 335300
rect 108356 335288 108362 335300
rect 136726 335288 136732 335300
rect 108356 335260 136732 335288
rect 108356 335248 108362 335260
rect 136726 335248 136732 335260
rect 136784 335248 136790 335300
rect 42610 335180 42616 335232
rect 42668 335220 42674 335232
rect 70394 335220 70400 335232
rect 42668 335192 70400 335220
rect 42668 335180 42674 335192
rect 70394 335180 70400 335192
rect 70452 335180 70458 335232
rect 104802 335180 104808 335232
rect 104860 335220 104866 335232
rect 128354 335220 128360 335232
rect 104860 335192 128360 335220
rect 104860 335180 104866 335192
rect 128354 335180 128360 335192
rect 128412 335180 128418 335232
rect 60550 335112 60556 335164
rect 60608 335152 60614 335164
rect 87598 335152 87604 335164
rect 60608 335124 87604 335152
rect 60608 335112 60614 335124
rect 87598 335112 87604 335124
rect 87656 335112 87662 335164
rect 112530 335112 112536 335164
rect 112588 335152 112594 335164
rect 113082 335152 113088 335164
rect 112588 335124 113088 335152
rect 112588 335112 112594 335124
rect 113082 335112 113088 335124
rect 113140 335152 113146 335164
rect 131206 335152 131212 335164
rect 113140 335124 131212 335152
rect 113140 335112 113146 335124
rect 131206 335112 131212 335124
rect 131264 335112 131270 335164
rect 57606 334636 57612 334688
rect 57664 334676 57670 334688
rect 104802 334676 104808 334688
rect 57664 334648 104808 334676
rect 57664 334636 57670 334648
rect 104802 334636 104808 334648
rect 104860 334636 104866 334688
rect 62022 334568 62028 334620
rect 62080 334608 62086 334620
rect 109862 334608 109868 334620
rect 62080 334580 109868 334608
rect 62080 334568 62086 334580
rect 109862 334568 109868 334580
rect 109920 334568 109926 334620
rect 70394 333956 70400 334008
rect 70452 333996 70458 334008
rect 71038 333996 71044 334008
rect 70452 333968 71044 333996
rect 70452 333956 70458 333968
rect 71038 333956 71044 333968
rect 71096 333956 71102 334008
rect 46566 333888 46572 333940
rect 46624 333928 46630 333940
rect 81434 333928 81440 333940
rect 46624 333900 81440 333928
rect 46624 333888 46630 333900
rect 81434 333888 81440 333900
rect 81492 333888 81498 333940
rect 95142 333888 95148 333940
rect 95200 333928 95206 333940
rect 127250 333928 127256 333940
rect 95200 333900 127256 333928
rect 95200 333888 95206 333900
rect 127250 333888 127256 333900
rect 127308 333888 127314 333940
rect 52178 333820 52184 333872
rect 52236 333860 52242 333872
rect 86218 333860 86224 333872
rect 52236 333832 86224 333860
rect 52236 333820 52242 333832
rect 86218 333820 86224 333832
rect 86276 333820 86282 333872
rect 104894 333820 104900 333872
rect 104952 333860 104958 333872
rect 135438 333860 135444 333872
rect 104952 333832 135444 333860
rect 104952 333820 104958 333832
rect 135438 333820 135444 333832
rect 135496 333820 135502 333872
rect 107654 333276 107660 333328
rect 107712 333316 107718 333328
rect 128630 333316 128636 333328
rect 107712 333288 128636 333316
rect 107712 333276 107718 333288
rect 128630 333276 128636 333288
rect 128688 333276 128694 333328
rect 61746 333208 61752 333260
rect 61804 333248 61810 333260
rect 115198 333248 115204 333260
rect 61804 333220 115204 333248
rect 61804 333208 61810 333220
rect 115198 333208 115204 333220
rect 115256 333208 115262 333260
rect 135438 333208 135444 333260
rect 135496 333248 135502 333260
rect 293954 333248 293960 333260
rect 135496 333220 293960 333248
rect 135496 333208 135502 333220
rect 293954 333208 293960 333220
rect 294012 333208 294018 333260
rect 81434 332596 81440 332648
rect 81492 332636 81498 332648
rect 82078 332636 82084 332648
rect 81492 332608 82084 332636
rect 81492 332596 81498 332608
rect 82078 332596 82084 332608
rect 82136 332596 82142 332648
rect 94590 332596 94596 332648
rect 94648 332636 94654 332648
rect 95142 332636 95148 332648
rect 94648 332608 95148 332636
rect 94648 332596 94654 332608
rect 95142 332596 95148 332608
rect 95200 332596 95206 332648
rect 57698 332528 57704 332580
rect 57756 332568 57762 332580
rect 90358 332568 90364 332580
rect 57756 332540 90364 332568
rect 57756 332528 57762 332540
rect 90358 332528 90364 332540
rect 90416 332528 90422 332580
rect 94498 332528 94504 332580
rect 94556 332568 94562 332580
rect 125778 332568 125784 332580
rect 94556 332540 125784 332568
rect 94556 332528 94562 332540
rect 125778 332528 125784 332540
rect 125836 332568 125842 332580
rect 128446 332568 128452 332580
rect 125836 332540 128452 332568
rect 125836 332528 125842 332540
rect 128446 332528 128452 332540
rect 128504 332528 128510 332580
rect 63310 331916 63316 331968
rect 63368 331956 63374 331968
rect 97994 331956 98000 331968
rect 63368 331928 98000 331956
rect 63368 331916 63374 331928
rect 97994 331916 98000 331928
rect 98052 331916 98058 331968
rect 106274 331916 106280 331968
rect 106332 331956 106338 331968
rect 118694 331956 118700 331968
rect 106332 331928 118700 331956
rect 106332 331916 106338 331928
rect 118694 331916 118700 331928
rect 118752 331916 118758 331968
rect 67450 331848 67456 331900
rect 67508 331888 67514 331900
rect 338114 331888 338120 331900
rect 67508 331860 338120 331888
rect 67508 331848 67514 331860
rect 338114 331848 338120 331860
rect 338172 331848 338178 331900
rect 105446 331168 105452 331220
rect 105504 331208 105510 331220
rect 136910 331208 136916 331220
rect 105504 331180 136916 331208
rect 105504 331168 105510 331180
rect 136910 331168 136916 331180
rect 136968 331208 136974 331220
rect 137186 331208 137192 331220
rect 136968 331180 137192 331208
rect 136968 331168 136974 331180
rect 137186 331168 137192 331180
rect 137244 331168 137250 331220
rect 137186 330488 137192 330540
rect 137244 330528 137250 330540
rect 335998 330528 336004 330540
rect 137244 330500 336004 330528
rect 137244 330488 137250 330500
rect 335998 330488 336004 330500
rect 336056 330488 336062 330540
rect 110598 329740 110604 329792
rect 110656 329780 110662 329792
rect 133138 329780 133144 329792
rect 110656 329752 133144 329780
rect 110656 329740 110662 329752
rect 133138 329740 133144 329752
rect 133196 329780 133202 329792
rect 133782 329780 133788 329792
rect 133196 329752 133788 329780
rect 133196 329740 133202 329752
rect 133782 329740 133788 329752
rect 133840 329740 133846 329792
rect 79962 329060 79968 329112
rect 80020 329100 80026 329112
rect 342254 329100 342260 329112
rect 80020 329072 342260 329100
rect 80020 329060 80026 329072
rect 342254 329060 342260 329072
rect 342312 329060 342318 329112
rect 97074 328380 97080 328432
rect 97132 328420 97138 328432
rect 129826 328420 129832 328432
rect 97132 328392 129832 328420
rect 97132 328380 97138 328392
rect 129826 328380 129832 328392
rect 129884 328420 129890 328432
rect 130562 328420 130568 328432
rect 129884 328392 130568 328420
rect 129884 328380 129890 328392
rect 130562 328380 130568 328392
rect 130620 328380 130626 328432
rect 49602 327768 49608 327820
rect 49660 327808 49666 327820
rect 105538 327808 105544 327820
rect 49660 327780 105544 327808
rect 49660 327768 49666 327780
rect 105538 327768 105544 327780
rect 105596 327768 105602 327820
rect 106090 327768 106096 327820
rect 106148 327808 106154 327820
rect 114462 327808 114468 327820
rect 106148 327780 114468 327808
rect 106148 327768 106154 327780
rect 114462 327768 114468 327780
rect 114520 327808 114526 327820
rect 138106 327808 138112 327820
rect 114520 327780 138112 327808
rect 114520 327768 114526 327780
rect 138106 327768 138112 327780
rect 138164 327768 138170 327820
rect 68830 327700 68836 327752
rect 68888 327740 68894 327752
rect 251174 327740 251180 327752
rect 68888 327712 251180 327740
rect 68888 327700 68894 327712
rect 251174 327700 251180 327712
rect 251232 327700 251238 327752
rect 3418 327088 3424 327140
rect 3476 327128 3482 327140
rect 49602 327128 49608 327140
rect 3476 327100 49608 327128
rect 3476 327088 3482 327100
rect 49602 327088 49608 327100
rect 49660 327088 49666 327140
rect 130562 327088 130568 327140
rect 130620 327128 130626 327140
rect 333974 327128 333980 327140
rect 130620 327100 333980 327128
rect 130620 327088 130626 327100
rect 333974 327088 333980 327100
rect 334032 327088 334038 327140
rect 68646 326476 68652 326528
rect 68704 326516 68710 326528
rect 115382 326516 115388 326528
rect 68704 326488 115388 326516
rect 68704 326476 68710 326488
rect 115382 326476 115388 326488
rect 115440 326476 115446 326528
rect 106182 326408 106188 326460
rect 106240 326448 106246 326460
rect 116118 326448 116124 326460
rect 106240 326420 116124 326448
rect 106240 326408 106246 326420
rect 116118 326408 116124 326420
rect 116176 326408 116182 326460
rect 68922 326340 68928 326392
rect 68980 326380 68986 326392
rect 309778 326380 309784 326392
rect 68980 326352 309784 326380
rect 68980 326340 68986 326352
rect 309778 326340 309784 326352
rect 309836 326340 309842 326392
rect 72418 324980 72424 325032
rect 72476 325020 72482 325032
rect 108298 325020 108304 325032
rect 72476 324992 108304 325020
rect 72476 324980 72482 324992
rect 108298 324980 108304 324992
rect 108356 324980 108362 325032
rect 73338 324912 73344 324964
rect 73396 324952 73402 324964
rect 116026 324952 116032 324964
rect 73396 324924 116032 324952
rect 73396 324912 73402 324924
rect 116026 324912 116032 324924
rect 116084 324912 116090 324964
rect 91002 324232 91008 324284
rect 91060 324272 91066 324284
rect 124306 324272 124312 324284
rect 91060 324244 124312 324272
rect 91060 324232 91066 324244
rect 124306 324232 124312 324244
rect 124364 324272 124370 324284
rect 128538 324272 128544 324284
rect 124364 324244 128544 324272
rect 124364 324232 124370 324244
rect 128538 324232 128544 324244
rect 128596 324232 128602 324284
rect 86310 323552 86316 323604
rect 86368 323592 86374 323604
rect 113910 323592 113916 323604
rect 86368 323564 113916 323592
rect 86368 323552 86374 323564
rect 113910 323552 113916 323564
rect 113968 323552 113974 323604
rect 66898 322192 66904 322244
rect 66956 322232 66962 322244
rect 309134 322232 309140 322244
rect 66956 322204 309140 322232
rect 66956 322192 66962 322204
rect 309134 322192 309140 322204
rect 309192 322192 309198 322244
rect 93946 320832 93952 320884
rect 94004 320872 94010 320884
rect 125686 320872 125692 320884
rect 94004 320844 125692 320872
rect 94004 320832 94010 320844
rect 125686 320832 125692 320844
rect 125744 320832 125750 320884
rect 118050 320492 118056 320544
rect 118108 320532 118114 320544
rect 120258 320532 120264 320544
rect 118108 320504 120264 320532
rect 118108 320492 118114 320504
rect 120258 320492 120264 320504
rect 120316 320492 120322 320544
rect 100938 320084 100944 320136
rect 100996 320124 101002 320136
rect 135346 320124 135352 320136
rect 100996 320096 135352 320124
rect 100996 320084 101002 320096
rect 135346 320084 135352 320096
rect 135404 320124 135410 320136
rect 136542 320124 136548 320136
rect 135404 320096 136548 320124
rect 135404 320084 135410 320096
rect 136542 320084 136548 320096
rect 136600 320084 136606 320136
rect 111242 320016 111248 320068
rect 111300 320056 111306 320068
rect 138198 320056 138204 320068
rect 111300 320028 138204 320056
rect 111300 320016 111306 320028
rect 138198 320016 138204 320028
rect 138256 320056 138262 320068
rect 138658 320056 138664 320068
rect 138256 320028 138664 320056
rect 138256 320016 138262 320028
rect 138658 320016 138664 320028
rect 138716 320016 138722 320068
rect 94038 319472 94044 319524
rect 94096 319512 94102 319524
rect 112438 319512 112444 319524
rect 94096 319484 112444 319512
rect 94096 319472 94102 319484
rect 112438 319472 112444 319484
rect 112496 319472 112502 319524
rect 136542 319472 136548 319524
rect 136600 319512 136606 319524
rect 266998 319512 267004 319524
rect 136600 319484 267004 319512
rect 136600 319472 136606 319484
rect 266998 319472 267004 319484
rect 267056 319472 267062 319524
rect 75270 319404 75276 319456
rect 75328 319444 75334 319456
rect 114554 319444 114560 319456
rect 75328 319416 114560 319444
rect 75328 319404 75334 319416
rect 114554 319404 114560 319416
rect 114612 319404 114618 319456
rect 138658 319404 138664 319456
rect 138716 319444 138722 319456
rect 339494 319444 339500 319456
rect 138716 319416 339500 319444
rect 138716 319404 138722 319416
rect 339494 319404 339500 319416
rect 339552 319404 339558 319456
rect 101398 318248 101404 318300
rect 101456 318288 101462 318300
rect 127066 318288 127072 318300
rect 101456 318260 127072 318288
rect 101456 318248 101462 318260
rect 127066 318248 127072 318260
rect 127124 318248 127130 318300
rect 67542 318180 67548 318232
rect 67600 318220 67606 318232
rect 115290 318220 115296 318232
rect 67600 318192 115296 318220
rect 67600 318180 67606 318192
rect 115290 318180 115296 318192
rect 115348 318180 115354 318232
rect 75178 318112 75184 318164
rect 75236 318152 75242 318164
rect 311894 318152 311900 318164
rect 75236 318124 311900 318152
rect 75236 318112 75242 318124
rect 311894 318112 311900 318124
rect 311952 318112 311958 318164
rect 84838 318044 84844 318096
rect 84896 318084 84902 318096
rect 345014 318084 345020 318096
rect 84896 318056 345020 318084
rect 84896 318044 84902 318056
rect 345014 318044 345020 318056
rect 345072 318044 345078 318096
rect 93210 316752 93216 316804
rect 93268 316792 93274 316804
rect 113818 316792 113824 316804
rect 93268 316764 113824 316792
rect 93268 316752 93274 316764
rect 113818 316752 113824 316764
rect 113876 316752 113882 316804
rect 71130 316684 71136 316736
rect 71188 316724 71194 316736
rect 320174 316724 320180 316736
rect 71188 316696 320180 316724
rect 71188 316684 71194 316696
rect 320174 316684 320180 316696
rect 320232 316684 320238 316736
rect 151998 315936 152004 315988
rect 152056 315976 152062 315988
rect 580350 315976 580356 315988
rect 152056 315948 580356 315976
rect 152056 315936 152062 315948
rect 580350 315936 580356 315948
rect 580408 315936 580414 315988
rect 120718 315256 120724 315308
rect 120776 315296 120782 315308
rect 151998 315296 152004 315308
rect 120776 315268 152004 315296
rect 120776 315256 120782 315268
rect 151998 315256 152004 315268
rect 152056 315256 152062 315308
rect 57698 313964 57704 314016
rect 57756 314004 57762 314016
rect 118786 314004 118792 314016
rect 57756 313976 118792 314004
rect 57756 313964 57762 313976
rect 118786 313964 118792 313976
rect 118844 313964 118850 314016
rect 88978 313896 88984 313948
rect 89036 313936 89042 313948
rect 216030 313936 216036 313948
rect 89036 313908 216036 313936
rect 89036 313896 89042 313908
rect 216030 313896 216036 313908
rect 216088 313896 216094 313948
rect 91094 313284 91100 313336
rect 91152 313324 91158 313336
rect 121638 313324 121644 313336
rect 91152 313296 121644 313324
rect 91152 313284 91158 313296
rect 121638 313284 121644 313296
rect 121696 313324 121702 313336
rect 582558 313324 582564 313336
rect 121696 313296 582564 313324
rect 121696 313284 121702 313296
rect 582558 313284 582564 313296
rect 582616 313284 582622 313336
rect 80054 312604 80060 312656
rect 80112 312644 80118 312656
rect 91094 312644 91100 312656
rect 80112 312616 91100 312644
rect 80112 312604 80118 312616
rect 91094 312604 91100 312616
rect 91152 312604 91158 312656
rect 97258 312604 97264 312656
rect 97316 312644 97322 312656
rect 125778 312644 125784 312656
rect 97316 312616 125784 312644
rect 97316 312604 97322 312616
rect 125778 312604 125784 312616
rect 125836 312644 125842 312656
rect 126882 312644 126888 312656
rect 125836 312616 126888 312644
rect 125836 312604 125842 312616
rect 126882 312604 126888 312616
rect 126940 312604 126946 312656
rect 89070 312536 89076 312588
rect 89128 312576 89134 312588
rect 209038 312576 209044 312588
rect 89128 312548 209044 312576
rect 89128 312536 89134 312548
rect 209038 312536 209044 312548
rect 209096 312536 209102 312588
rect 126882 311856 126888 311908
rect 126940 311896 126946 311908
rect 579982 311896 579988 311908
rect 126940 311868 579988 311896
rect 126940 311856 126946 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 311788 3516 311840
rect 3568 311828 3574 311840
rect 50706 311828 50712 311840
rect 3568 311800 50712 311828
rect 3568 311788 3574 311800
rect 50706 311788 50712 311800
rect 50764 311788 50770 311840
rect 50706 311108 50712 311160
rect 50764 311148 50770 311160
rect 115934 311148 115940 311160
rect 50764 311120 115940 311148
rect 50764 311108 50770 311120
rect 115934 311108 115940 311120
rect 115992 311108 115998 311160
rect 74442 309816 74448 309868
rect 74500 309856 74506 309868
rect 119706 309856 119712 309868
rect 74500 309828 119712 309856
rect 74500 309816 74506 309828
rect 119706 309816 119712 309828
rect 119764 309816 119770 309868
rect 83458 309748 83464 309800
rect 83516 309788 83522 309800
rect 322198 309788 322204 309800
rect 83516 309760 322204 309788
rect 83516 309748 83522 309760
rect 322198 309748 322204 309760
rect 322256 309748 322262 309800
rect 88334 309136 88340 309188
rect 88392 309176 88398 309188
rect 280798 309176 280804 309188
rect 88392 309148 280804 309176
rect 88392 309136 88398 309148
rect 280798 309136 280804 309148
rect 280856 309136 280862 309188
rect 113082 308388 113088 308440
rect 113140 308428 113146 308440
rect 253934 308428 253940 308440
rect 113140 308400 253940 308428
rect 113140 308388 113146 308400
rect 253934 308388 253940 308400
rect 253992 308388 253998 308440
rect 74626 307912 74632 307964
rect 74684 307952 74690 307964
rect 145558 307952 145564 307964
rect 74684 307924 145564 307952
rect 74684 307912 74690 307924
rect 145558 307912 145564 307924
rect 145616 307912 145622 307964
rect 81434 307844 81440 307896
rect 81492 307884 81498 307896
rect 155218 307884 155224 307896
rect 81492 307856 155224 307884
rect 81492 307844 81498 307856
rect 155218 307844 155224 307856
rect 155276 307844 155282 307896
rect 78766 307776 78772 307828
rect 78824 307816 78830 307828
rect 226978 307816 226984 307828
rect 78824 307788 226984 307816
rect 78824 307776 78830 307788
rect 226978 307776 226984 307788
rect 227036 307776 227042 307828
rect 79318 307164 79324 307216
rect 79376 307204 79382 307216
rect 120074 307204 120080 307216
rect 79376 307176 120080 307204
rect 79376 307164 79382 307176
rect 120074 307164 120080 307176
rect 120132 307164 120138 307216
rect 65610 307096 65616 307148
rect 65668 307136 65674 307148
rect 213178 307136 213184 307148
rect 65668 307108 213184 307136
rect 65668 307096 65674 307108
rect 213178 307096 213184 307108
rect 213236 307096 213242 307148
rect 103330 307028 103336 307080
rect 103388 307068 103394 307080
rect 266354 307068 266360 307080
rect 103388 307040 266360 307068
rect 103388 307028 103394 307040
rect 266354 307028 266360 307040
rect 266412 307028 266418 307080
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 11698 306320 11704 306332
rect 3568 306292 11704 306320
rect 3568 306280 3574 306292
rect 11698 306280 11704 306292
rect 11756 306280 11762 306332
rect 71038 305668 71044 305720
rect 71096 305708 71102 305720
rect 186958 305708 186964 305720
rect 71096 305680 186964 305708
rect 71096 305668 71102 305680
rect 186958 305668 186964 305680
rect 187016 305668 187022 305720
rect 100018 305600 100024 305652
rect 100076 305640 100082 305652
rect 321554 305640 321560 305652
rect 100076 305612 321560 305640
rect 100076 305600 100082 305612
rect 321554 305600 321560 305612
rect 321612 305600 321618 305652
rect 89714 304988 89720 305040
rect 89772 305028 89778 305040
rect 171778 305028 171784 305040
rect 89772 305000 171784 305028
rect 89772 304988 89778 305000
rect 171778 304988 171784 305000
rect 171836 304988 171842 305040
rect 80698 304308 80704 304360
rect 80756 304348 80762 304360
rect 129826 304348 129832 304360
rect 80756 304320 129832 304348
rect 80756 304308 80762 304320
rect 129826 304308 129832 304320
rect 129884 304308 129890 304360
rect 48130 304240 48136 304292
rect 48188 304280 48194 304292
rect 71774 304280 71780 304292
rect 48188 304252 71780 304280
rect 48188 304240 48194 304252
rect 71774 304240 71780 304252
rect 71832 304240 71838 304292
rect 109678 304240 109684 304292
rect 109736 304280 109742 304292
rect 119338 304280 119344 304292
rect 109736 304252 119344 304280
rect 109736 304240 109742 304252
rect 119338 304240 119344 304252
rect 119396 304280 119402 304292
rect 582834 304280 582840 304292
rect 119396 304252 582840 304280
rect 119396 304240 119402 304252
rect 582834 304240 582840 304252
rect 582892 304240 582898 304292
rect 75914 303764 75920 303816
rect 75972 303804 75978 303816
rect 163498 303804 163504 303816
rect 75972 303776 163504 303804
rect 75972 303764 75978 303776
rect 163498 303764 163504 303776
rect 163556 303764 163562 303816
rect 66162 303696 66168 303748
rect 66220 303736 66226 303748
rect 169018 303736 169024 303748
rect 66220 303708 169024 303736
rect 66220 303696 66226 303708
rect 169018 303696 169024 303708
rect 169076 303696 169082 303748
rect 85574 303628 85580 303680
rect 85632 303668 85638 303680
rect 278038 303668 278044 303680
rect 85632 303640 278044 303668
rect 85632 303628 85638 303640
rect 278038 303628 278044 303640
rect 278096 303628 278102 303680
rect 65978 302880 65984 302932
rect 66036 302920 66042 302932
rect 131114 302920 131120 302932
rect 66036 302892 131120 302920
rect 66036 302880 66042 302892
rect 131114 302880 131120 302892
rect 131172 302880 131178 302932
rect 87506 302404 87512 302456
rect 87564 302444 87570 302456
rect 222838 302444 222844 302456
rect 87564 302416 222844 302444
rect 87564 302404 87570 302416
rect 222838 302404 222844 302416
rect 222896 302404 222902 302456
rect 85666 302336 85672 302388
rect 85724 302376 85730 302388
rect 231118 302376 231124 302388
rect 85724 302348 231124 302376
rect 85724 302336 85730 302348
rect 231118 302336 231124 302348
rect 231176 302336 231182 302388
rect 112438 302268 112444 302320
rect 112496 302308 112502 302320
rect 272518 302308 272524 302320
rect 112496 302280 272524 302308
rect 112496 302268 112502 302280
rect 272518 302268 272524 302280
rect 272576 302268 272582 302320
rect 71866 302200 71872 302252
rect 71924 302240 71930 302252
rect 309226 302240 309232 302252
rect 71924 302212 309232 302240
rect 71924 302200 71930 302212
rect 309226 302200 309232 302212
rect 309284 302200 309290 302252
rect 90358 301520 90364 301572
rect 90416 301560 90422 301572
rect 195238 301560 195244 301572
rect 90416 301532 195244 301560
rect 90416 301520 90422 301532
rect 195238 301520 195244 301532
rect 195296 301520 195302 301572
rect 71038 301452 71044 301504
rect 71096 301492 71102 301504
rect 134150 301492 134156 301504
rect 71096 301464 134156 301492
rect 71096 301452 71102 301464
rect 134150 301452 134156 301464
rect 134208 301492 134214 301504
rect 582650 301492 582656 301504
rect 134208 301464 582656 301492
rect 134208 301452 134214 301464
rect 582650 301452 582656 301464
rect 582708 301452 582714 301504
rect 84194 301044 84200 301096
rect 84252 301084 84258 301096
rect 180150 301084 180156 301096
rect 84252 301056 180156 301084
rect 84252 301044 84258 301056
rect 180150 301044 180156 301056
rect 180208 301044 180214 301096
rect 106918 300976 106924 301028
rect 106976 301016 106982 301028
rect 203518 301016 203524 301028
rect 106976 300988 203524 301016
rect 106976 300976 106982 300988
rect 203518 300976 203524 300988
rect 203576 300976 203582 301028
rect 74534 300908 74540 300960
rect 74592 300948 74598 300960
rect 240410 300948 240416 300960
rect 74592 300920 240416 300948
rect 74592 300908 74598 300920
rect 240410 300908 240416 300920
rect 240468 300908 240474 300960
rect 110966 300840 110972 300892
rect 111024 300880 111030 300892
rect 302326 300880 302332 300892
rect 111024 300852 302332 300880
rect 111024 300840 111030 300852
rect 302326 300840 302332 300852
rect 302384 300840 302390 300892
rect 93118 300296 93124 300348
rect 93176 300336 93182 300348
rect 125870 300336 125876 300348
rect 93176 300308 125876 300336
rect 93176 300296 93182 300308
rect 125870 300296 125876 300308
rect 125928 300296 125934 300348
rect 86218 300228 86224 300280
rect 86276 300268 86282 300280
rect 124306 300268 124312 300280
rect 86276 300240 124312 300268
rect 86276 300228 86282 300240
rect 124306 300228 124312 300240
rect 124364 300228 124370 300280
rect 61930 300160 61936 300212
rect 61988 300200 61994 300212
rect 116578 300200 116584 300212
rect 61988 300172 116584 300200
rect 61988 300160 61994 300172
rect 116578 300160 116584 300172
rect 116636 300160 116642 300212
rect 42702 300092 42708 300144
rect 42760 300132 42766 300144
rect 123110 300132 123116 300144
rect 42760 300104 123116 300132
rect 42760 300092 42766 300104
rect 123110 300092 123116 300104
rect 123168 300092 123174 300144
rect 81894 299548 81900 299600
rect 81952 299588 81958 299600
rect 198182 299588 198188 299600
rect 81952 299560 198188 299588
rect 81952 299548 81958 299560
rect 198182 299548 198188 299560
rect 198240 299548 198246 299600
rect 102134 299480 102140 299532
rect 102192 299520 102198 299532
rect 224218 299520 224224 299532
rect 102192 299492 224224 299520
rect 102192 299480 102198 299492
rect 224218 299480 224224 299492
rect 224276 299480 224282 299532
rect 61838 298732 61844 298784
rect 61896 298772 61902 298784
rect 127158 298772 127164 298784
rect 61896 298744 127164 298772
rect 61896 298732 61902 298744
rect 127158 298732 127164 298744
rect 127216 298732 127222 298784
rect 73246 298392 73252 298444
rect 73304 298432 73310 298444
rect 157978 298432 157984 298444
rect 73304 298404 157984 298432
rect 73304 298392 73310 298404
rect 157978 298392 157984 298404
rect 158036 298392 158042 298444
rect 82906 298324 82912 298376
rect 82964 298364 82970 298376
rect 178770 298364 178776 298376
rect 82964 298336 178776 298364
rect 82964 298324 82970 298336
rect 178770 298324 178776 298336
rect 178828 298324 178834 298376
rect 75178 298256 75184 298308
rect 75236 298296 75242 298308
rect 227070 298296 227076 298308
rect 75236 298268 227076 298296
rect 75236 298256 75242 298268
rect 227070 298256 227076 298268
rect 227128 298256 227134 298308
rect 102870 298188 102876 298240
rect 102928 298228 102934 298240
rect 262214 298228 262220 298240
rect 102928 298200 262220 298228
rect 102928 298188 102934 298200
rect 262214 298188 262220 298200
rect 262272 298188 262278 298240
rect 103422 298120 103428 298172
rect 103480 298160 103486 298172
rect 104802 298160 104808 298172
rect 103480 298132 104808 298160
rect 103480 298120 103486 298132
rect 104802 298120 104808 298132
rect 104860 298120 104866 298172
rect 106182 298120 106188 298172
rect 106240 298160 106246 298172
rect 582374 298160 582380 298172
rect 106240 298132 582380 298160
rect 106240 298120 106246 298132
rect 582374 298120 582380 298132
rect 582432 298120 582438 298172
rect 48038 297508 48044 297560
rect 48096 297548 48102 297560
rect 77754 297548 77760 297560
rect 48096 297520 77760 297548
rect 48096 297508 48102 297520
rect 77754 297508 77760 297520
rect 77812 297508 77818 297560
rect 60458 297440 60464 297492
rect 60516 297480 60522 297492
rect 124398 297480 124404 297492
rect 60516 297452 124404 297480
rect 60516 297440 60522 297452
rect 124398 297440 124404 297452
rect 124456 297440 124462 297492
rect 41230 297372 41236 297424
rect 41288 297412 41294 297424
rect 117222 297412 117228 297424
rect 41288 297384 117228 297412
rect 41288 297372 41294 297384
rect 117222 297372 117228 297384
rect 117280 297372 117286 297424
rect 117958 296964 117964 297016
rect 118016 297004 118022 297016
rect 123018 297004 123024 297016
rect 118016 296976 123024 297004
rect 118016 296964 118022 296976
rect 123018 296964 123024 296976
rect 123076 296964 123082 297016
rect 88702 296896 88708 296948
rect 88760 296936 88766 296948
rect 151078 296936 151084 296948
rect 88760 296908 151084 296936
rect 88760 296896 88766 296908
rect 151078 296896 151084 296908
rect 151136 296896 151142 296948
rect 100938 296828 100944 296880
rect 100996 296868 101002 296880
rect 182818 296868 182824 296880
rect 100996 296840 182824 296868
rect 100996 296828 101002 296840
rect 182818 296828 182824 296840
rect 182876 296828 182882 296880
rect 93210 296760 93216 296812
rect 93268 296800 93274 296812
rect 202230 296800 202236 296812
rect 93268 296772 202236 296800
rect 93268 296760 93274 296772
rect 202230 296760 202236 296772
rect 202288 296760 202294 296812
rect 110598 296692 110604 296744
rect 110656 296732 110662 296744
rect 225598 296732 225604 296744
rect 110656 296704 225604 296732
rect 110656 296692 110662 296704
rect 225598 296692 225604 296704
rect 225656 296692 225662 296744
rect 29638 295740 29644 295792
rect 29696 295780 29702 295792
rect 118050 295780 118056 295792
rect 29696 295752 118056 295780
rect 29696 295740 29702 295752
rect 118050 295740 118056 295752
rect 118108 295740 118114 295792
rect 91922 295672 91928 295724
rect 91980 295712 91986 295724
rect 141418 295712 141424 295724
rect 91980 295684 141424 295712
rect 91980 295672 91986 295684
rect 141418 295672 141424 295684
rect 141476 295672 141482 295724
rect 117682 295604 117688 295656
rect 117740 295644 117746 295656
rect 199378 295644 199384 295656
rect 117740 295616 199384 295644
rect 117740 295604 117746 295616
rect 199378 295604 199384 295616
rect 199436 295604 199442 295656
rect 83550 295536 83556 295588
rect 83608 295576 83614 295588
rect 181438 295576 181444 295588
rect 83608 295548 181444 295576
rect 83608 295536 83614 295548
rect 181438 295536 181444 295548
rect 181496 295536 181502 295588
rect 99650 295468 99656 295520
rect 99708 295508 99714 295520
rect 256694 295508 256700 295520
rect 99708 295480 256700 295508
rect 99708 295468 99714 295480
rect 256694 295468 256700 295480
rect 256752 295468 256758 295520
rect 68830 295400 68836 295452
rect 68888 295440 68894 295452
rect 234614 295440 234620 295452
rect 68888 295412 234620 295440
rect 68888 295400 68894 295412
rect 234614 295400 234620 295412
rect 234672 295400 234678 295452
rect 17218 295332 17224 295384
rect 17276 295372 17282 295384
rect 92566 295372 92572 295384
rect 17276 295344 92572 295372
rect 17276 295332 17282 295344
rect 92566 295332 92572 295344
rect 92624 295372 92630 295384
rect 92934 295372 92940 295384
rect 92624 295344 92940 295372
rect 92624 295332 92630 295344
rect 92934 295332 92940 295344
rect 92992 295332 92998 295384
rect 111886 295332 111892 295384
rect 111944 295372 111950 295384
rect 307846 295372 307852 295384
rect 111944 295344 307852 295372
rect 111944 295332 111950 295344
rect 307846 295332 307852 295344
rect 307904 295332 307910 295384
rect 87414 294788 87420 294840
rect 87472 294828 87478 294840
rect 106918 294828 106924 294840
rect 87472 294800 106924 294828
rect 87472 294788 87478 294800
rect 106918 294788 106924 294800
rect 106976 294788 106982 294840
rect 79042 294760 79048 294772
rect 55186 294732 79048 294760
rect 25498 294584 25504 294636
rect 25556 294624 25562 294636
rect 53650 294624 53656 294636
rect 25556 294596 53656 294624
rect 25556 294584 25562 294596
rect 53650 294584 53656 294596
rect 53708 294624 53714 294636
rect 55186 294624 55214 294732
rect 79042 294720 79048 294732
rect 79100 294720 79106 294772
rect 84838 294720 84844 294772
rect 84896 294760 84902 294772
rect 104158 294760 104164 294772
rect 84896 294732 104164 294760
rect 84896 294720 84902 294732
rect 104158 294720 104164 294732
rect 104216 294720 104222 294772
rect 57790 294652 57796 294704
rect 57848 294692 57854 294704
rect 91278 294692 91284 294704
rect 57848 294664 91284 294692
rect 57848 294652 57854 294664
rect 91278 294652 91284 294664
rect 91336 294652 91342 294704
rect 53708 294596 55214 294624
rect 53708 294584 53714 294596
rect 70670 294584 70676 294636
rect 70728 294624 70734 294636
rect 115842 294624 115848 294636
rect 70728 294596 115848 294624
rect 70728 294584 70734 294596
rect 115842 294584 115848 294596
rect 115900 294584 115906 294636
rect 106734 294380 106740 294432
rect 106792 294420 106798 294432
rect 112438 294420 112444 294432
rect 106792 294392 112444 294420
rect 106792 294380 106798 294392
rect 112438 294380 112444 294392
rect 112496 294380 112502 294432
rect 71774 294312 71780 294364
rect 71832 294352 71838 294364
rect 72326 294352 72332 294364
rect 71832 294324 72332 294352
rect 71832 294312 71838 294324
rect 72326 294312 72332 294324
rect 72384 294312 72390 294364
rect 85482 294312 85488 294364
rect 85540 294352 85546 294364
rect 86310 294352 86316 294364
rect 85540 294324 86316 294352
rect 85540 294312 85546 294324
rect 86310 294312 86316 294324
rect 86368 294312 86374 294364
rect 93946 294312 93952 294364
rect 94004 294352 94010 294364
rect 94774 294352 94780 294364
rect 94004 294324 94780 294352
rect 94004 294312 94010 294324
rect 94774 294312 94780 294324
rect 94832 294312 94838 294364
rect 108022 294312 108028 294364
rect 108080 294352 108086 294364
rect 117130 294352 117136 294364
rect 108080 294324 117136 294352
rect 108080 294312 108086 294324
rect 117130 294312 117136 294324
rect 117188 294312 117194 294364
rect 71314 294244 71320 294296
rect 71372 294284 71378 294296
rect 72418 294284 72424 294296
rect 71372 294256 72424 294284
rect 71372 294244 71378 294256
rect 72418 294244 72424 294256
rect 72476 294244 72482 294296
rect 85574 294244 85580 294296
rect 85632 294284 85638 294296
rect 86494 294284 86500 294296
rect 85632 294256 86500 294284
rect 85632 294244 85638 294256
rect 86494 294244 86500 294256
rect 86552 294244 86558 294296
rect 105446 294244 105452 294296
rect 105504 294284 105510 294296
rect 125502 294284 125508 294296
rect 105504 294256 125508 294284
rect 105504 294244 105510 294256
rect 125502 294244 125508 294256
rect 125560 294244 125566 294296
rect 113818 294176 113824 294228
rect 113876 294216 113882 294228
rect 152458 294216 152464 294228
rect 113876 294188 152464 294216
rect 113876 294176 113882 294188
rect 152458 294176 152464 294188
rect 152516 294176 152522 294228
rect 112530 294108 112536 294160
rect 112588 294148 112594 294160
rect 255314 294148 255320 294160
rect 112588 294120 255320 294148
rect 112588 294108 112594 294120
rect 255314 294108 255320 294120
rect 255372 294108 255378 294160
rect 80974 294040 80980 294092
rect 81032 294080 81038 294092
rect 239030 294080 239036 294092
rect 81032 294052 239036 294080
rect 81032 294040 81038 294052
rect 239030 294040 239036 294052
rect 239088 294040 239094 294092
rect 47578 293972 47584 294024
rect 47636 294012 47642 294024
rect 101398 294012 101404 294024
rect 47636 293984 101404 294012
rect 47636 293972 47642 293984
rect 101398 293972 101404 293984
rect 101456 294012 101462 294024
rect 101582 294012 101588 294024
rect 101456 293984 101588 294012
rect 101456 293972 101462 293984
rect 101582 293972 101588 293984
rect 101640 293972 101646 294024
rect 104158 293972 104164 294024
rect 104216 294012 104222 294024
rect 110414 294012 110420 294024
rect 104216 293984 110420 294012
rect 104216 293972 104222 293984
rect 110414 293972 110420 293984
rect 110472 293972 110478 294024
rect 117222 293972 117228 294024
rect 117280 294012 117286 294024
rect 119614 294012 119620 294024
rect 117280 293984 119620 294012
rect 117280 293972 117286 293984
rect 119614 293972 119620 293984
rect 119672 293972 119678 294024
rect 303706 294012 303712 294024
rect 119724 293984 303712 294012
rect 119338 293904 119344 293956
rect 119396 293944 119402 293956
rect 119724 293944 119752 293984
rect 303706 293972 303712 293984
rect 303764 293972 303770 294024
rect 119396 293916 119752 293944
rect 119396 293904 119402 293916
rect 125502 293904 125508 293956
rect 125560 293944 125566 293956
rect 130010 293944 130016 293956
rect 125560 293916 130016 293944
rect 125560 293904 125566 293916
rect 130010 293904 130016 293916
rect 130068 293904 130074 293956
rect 115198 293292 115204 293344
rect 115256 293332 115262 293344
rect 125686 293332 125692 293344
rect 115256 293304 125692 293332
rect 115256 293292 115262 293304
rect 125686 293292 125692 293304
rect 125744 293292 125750 293344
rect 53098 293224 53104 293276
rect 53156 293264 53162 293276
rect 54478 293264 54484 293276
rect 53156 293236 54484 293264
rect 53156 293224 53162 293236
rect 54478 293224 54484 293236
rect 54536 293264 54542 293276
rect 97074 293264 97080 293276
rect 54536 293236 97080 293264
rect 54536 293224 54542 293236
rect 97074 293224 97080 293236
rect 97132 293224 97138 293276
rect 110414 293224 110420 293276
rect 110472 293264 110478 293276
rect 278130 293264 278136 293276
rect 110472 293236 278136 293264
rect 110472 293224 110478 293236
rect 278130 293224 278136 293236
rect 278188 293224 278194 293276
rect 93854 292748 93860 292800
rect 93912 292788 93918 292800
rect 133138 292788 133144 292800
rect 93912 292760 133144 292788
rect 93912 292748 93918 292760
rect 133138 292748 133144 292760
rect 133196 292748 133202 292800
rect 77110 292680 77116 292732
rect 77168 292720 77174 292732
rect 125226 292720 125232 292732
rect 77168 292692 125232 292720
rect 77168 292680 77174 292692
rect 125226 292680 125232 292692
rect 125284 292720 125290 292732
rect 125502 292720 125508 292732
rect 125284 292692 125508 292720
rect 125284 292680 125290 292692
rect 125502 292680 125508 292692
rect 125560 292680 125566 292732
rect 103514 292612 103520 292664
rect 103572 292652 103578 292664
rect 271138 292652 271144 292664
rect 103572 292624 271144 292652
rect 103572 292612 103578 292624
rect 271138 292612 271144 292624
rect 271196 292612 271202 292664
rect 55122 292544 55128 292596
rect 55180 292584 55186 292596
rect 96430 292584 96436 292596
rect 55180 292556 96436 292584
rect 55180 292544 55186 292556
rect 96430 292544 96436 292556
rect 96488 292544 96494 292596
rect 97718 292544 97724 292596
rect 97776 292584 97782 292596
rect 273898 292584 273904 292596
rect 97776 292556 273904 292584
rect 97776 292544 97782 292556
rect 273898 292544 273904 292556
rect 273956 292544 273962 292596
rect 121638 292476 121644 292528
rect 121696 292516 121702 292528
rect 147858 292516 147864 292528
rect 121696 292488 147864 292516
rect 121696 292476 121702 292488
rect 147858 292476 147864 292488
rect 147916 292476 147922 292528
rect 125502 292408 125508 292460
rect 125560 292448 125566 292460
rect 142430 292448 142436 292460
rect 125560 292420 142436 292448
rect 125560 292408 125566 292420
rect 142430 292408 142436 292420
rect 142488 292408 142494 292460
rect 117130 291932 117136 291984
rect 117188 291972 117194 291984
rect 117188 291944 132494 291972
rect 117188 291932 117194 291944
rect 109586 291864 109592 291916
rect 109644 291904 109650 291916
rect 109644 291876 113174 291904
rect 109644 291864 109650 291876
rect 113146 291224 113174 291876
rect 117314 291864 117320 291916
rect 117372 291904 117378 291916
rect 132466 291904 132494 291944
rect 166350 291904 166356 291916
rect 117372 291876 122834 291904
rect 132466 291876 166356 291904
rect 117372 291864 117378 291876
rect 122806 291836 122834 291876
rect 166350 291864 166356 291876
rect 166408 291864 166414 291916
rect 307938 291836 307944 291848
rect 122806 291808 307944 291836
rect 307938 291796 307944 291808
rect 307996 291796 308002 291848
rect 290458 291224 290464 291236
rect 113146 291196 290464 291224
rect 290458 291184 290464 291196
rect 290516 291184 290522 291236
rect 32398 290436 32404 290488
rect 32456 290476 32462 290488
rect 67634 290476 67640 290488
rect 32456 290448 67640 290476
rect 32456 290436 32462 290448
rect 67634 290436 67640 290448
rect 67692 290436 67698 290488
rect 121638 289824 121644 289876
rect 121696 289864 121702 289876
rect 234706 289864 234712 289876
rect 121696 289836 234712 289864
rect 121696 289824 121702 289836
rect 234706 289824 234712 289836
rect 234764 289824 234770 289876
rect 66162 289756 66168 289808
rect 66220 289796 66226 289808
rect 68186 289796 68192 289808
rect 66220 289768 68192 289796
rect 66220 289756 66226 289768
rect 68186 289756 68192 289768
rect 68244 289756 68250 289808
rect 121730 288396 121736 288448
rect 121788 288436 121794 288448
rect 287330 288436 287336 288448
rect 121788 288408 287336 288436
rect 121788 288396 121794 288408
rect 287330 288396 287336 288408
rect 287388 288396 287394 288448
rect 49510 288328 49516 288380
rect 49568 288368 49574 288380
rect 67634 288368 67640 288380
rect 49568 288340 67640 288368
rect 49568 288328 49574 288340
rect 67634 288328 67640 288340
rect 67692 288328 67698 288380
rect 121638 288328 121644 288380
rect 121696 288368 121702 288380
rect 140958 288368 140964 288380
rect 121696 288340 140964 288368
rect 121696 288328 121702 288340
rect 140958 288328 140964 288340
rect 141016 288368 141022 288380
rect 141602 288368 141608 288380
rect 141016 288340 141608 288368
rect 141016 288328 141022 288340
rect 141602 288328 141608 288340
rect 141660 288328 141666 288380
rect 141602 287648 141608 287700
rect 141660 287688 141666 287700
rect 467098 287688 467104 287700
rect 141660 287660 467104 287688
rect 141660 287648 141666 287660
rect 467098 287648 467104 287660
rect 467156 287648 467162 287700
rect 121822 287036 121828 287088
rect 121880 287076 121886 287088
rect 224310 287076 224316 287088
rect 121880 287048 224316 287076
rect 121880 287036 121886 287048
rect 224310 287036 224316 287048
rect 224368 287036 224374 287088
rect 121730 286900 121736 286952
rect 121788 286940 121794 286952
rect 125870 286940 125876 286952
rect 121788 286912 125876 286940
rect 121788 286900 121794 286912
rect 125870 286900 125876 286912
rect 125928 286900 125934 286952
rect 121638 286832 121644 286884
rect 121696 286872 121702 286884
rect 132678 286872 132684 286884
rect 121696 286844 132684 286872
rect 121696 286832 121702 286844
rect 132678 286832 132684 286844
rect 132736 286832 132742 286884
rect 121546 286628 121552 286680
rect 121604 286668 121610 286680
rect 123110 286668 123116 286680
rect 121604 286640 123116 286668
rect 121604 286628 121610 286640
rect 123110 286628 123116 286640
rect 123168 286628 123174 286680
rect 125870 286288 125876 286340
rect 125928 286328 125934 286340
rect 468478 286328 468484 286340
rect 125928 286300 468484 286328
rect 125928 286288 125934 286300
rect 468478 286288 468484 286300
rect 468536 286288 468542 286340
rect 46750 284316 46756 284368
rect 46808 284356 46814 284368
rect 67634 284356 67640 284368
rect 46808 284328 67640 284356
rect 46808 284316 46814 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 121638 284316 121644 284368
rect 121696 284356 121702 284368
rect 214650 284356 214656 284368
rect 121696 284328 214656 284356
rect 121696 284316 121702 284328
rect 214650 284316 214656 284328
rect 214708 284316 214714 284368
rect 56502 284248 56508 284300
rect 56560 284288 56566 284300
rect 67726 284288 67732 284300
rect 56560 284260 67732 284288
rect 56560 284248 56566 284260
rect 67726 284248 67732 284260
rect 67784 284248 67790 284300
rect 121546 284248 121552 284300
rect 121604 284288 121610 284300
rect 143718 284288 143724 284300
rect 121604 284260 143724 284288
rect 121604 284248 121610 284260
rect 143718 284248 143724 284260
rect 143776 284248 143782 284300
rect 121546 282888 121552 282940
rect 121604 282928 121610 282940
rect 282914 282928 282920 282940
rect 121604 282900 282920 282928
rect 121604 282888 121610 282900
rect 282914 282888 282920 282900
rect 282972 282888 282978 282940
rect 43990 282820 43996 282872
rect 44048 282860 44054 282872
rect 67634 282860 67640 282872
rect 44048 282832 67640 282860
rect 44048 282820 44054 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 222930 282140 222936 282192
rect 222988 282180 222994 282192
rect 336734 282180 336740 282192
rect 222988 282152 336740 282180
rect 222988 282140 222994 282152
rect 336734 282140 336740 282152
rect 336792 282140 336798 282192
rect 121638 281596 121644 281648
rect 121696 281636 121702 281648
rect 221458 281636 221464 281648
rect 121696 281608 221464 281636
rect 121696 281596 121702 281608
rect 221458 281596 221464 281608
rect 221516 281596 221522 281648
rect 121546 281528 121552 281580
rect 121604 281568 121610 281580
rect 227162 281568 227168 281580
rect 121604 281540 227168 281568
rect 121604 281528 121610 281540
rect 227162 281528 227168 281540
rect 227220 281528 227226 281580
rect 50798 280168 50804 280220
rect 50856 280208 50862 280220
rect 67634 280208 67640 280220
rect 50856 280180 67640 280208
rect 50856 280168 50862 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121546 280168 121552 280220
rect 121604 280208 121610 280220
rect 284570 280208 284576 280220
rect 121604 280180 284576 280208
rect 121604 280168 121610 280180
rect 284570 280168 284576 280180
rect 284628 280168 284634 280220
rect 33134 280100 33140 280152
rect 33192 280140 33198 280152
rect 34146 280140 34152 280152
rect 33192 280112 34152 280140
rect 33192 280100 33198 280112
rect 34146 280100 34152 280112
rect 34204 280140 34210 280152
rect 67726 280140 67732 280152
rect 34204 280112 67732 280140
rect 34204 280100 34210 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 55030 280032 55036 280084
rect 55088 280072 55094 280084
rect 67634 280072 67640 280084
rect 55088 280044 67640 280072
rect 55088 280032 55094 280044
rect 67634 280032 67640 280044
rect 67692 280032 67698 280084
rect 4798 279420 4804 279472
rect 4856 279460 4862 279472
rect 33134 279460 33140 279472
rect 4856 279432 33140 279460
rect 4856 279420 4862 279432
rect 33134 279420 33140 279432
rect 33192 279420 33198 279472
rect 271230 279420 271236 279472
rect 271288 279460 271294 279472
rect 346394 279460 346400 279472
rect 271288 279432 346400 279460
rect 271288 279420 271294 279432
rect 346394 279420 346400 279432
rect 346452 279420 346458 279472
rect 121546 278808 121552 278860
rect 121604 278848 121610 278860
rect 204990 278848 204996 278860
rect 121604 278820 204996 278848
rect 121604 278808 121610 278820
rect 204990 278808 204996 278820
rect 205048 278808 205054 278860
rect 121638 278740 121644 278792
rect 121696 278780 121702 278792
rect 269850 278780 269856 278792
rect 121696 278752 269856 278780
rect 121696 278740 121702 278752
rect 269850 278740 269856 278752
rect 269908 278740 269914 278792
rect 273990 277992 273996 278044
rect 274048 278032 274054 278044
rect 347774 278032 347780 278044
rect 274048 278004 347780 278032
rect 274048 277992 274054 278004
rect 347774 277992 347780 278004
rect 347832 277992 347838 278044
rect 55030 277448 55036 277500
rect 55088 277488 55094 277500
rect 67634 277488 67640 277500
rect 55088 277460 67640 277488
rect 55088 277448 55094 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 121546 277448 121552 277500
rect 121604 277488 121610 277500
rect 192478 277488 192484 277500
rect 121604 277460 192484 277488
rect 121604 277448 121610 277460
rect 192478 277448 192484 277460
rect 192536 277448 192542 277500
rect 52086 277380 52092 277432
rect 52144 277420 52150 277432
rect 67726 277420 67732 277432
rect 52144 277392 67732 277420
rect 52144 277380 52150 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121638 277380 121644 277432
rect 121696 277420 121702 277432
rect 302234 277420 302240 277432
rect 121696 277392 302240 277420
rect 121696 277380 121702 277392
rect 302234 277380 302240 277392
rect 302292 277380 302298 277432
rect 121546 276632 121552 276684
rect 121604 276672 121610 276684
rect 129918 276672 129924 276684
rect 121604 276644 129924 276672
rect 121604 276632 121610 276644
rect 129918 276632 129924 276644
rect 129976 276632 129982 276684
rect 53558 276020 53564 276072
rect 53616 276060 53622 276072
rect 67634 276060 67640 276072
rect 53616 276032 67640 276060
rect 53616 276020 53622 276032
rect 67634 276020 67640 276032
rect 67692 276020 67698 276072
rect 129918 276020 129924 276072
rect 129976 276060 129982 276072
rect 130378 276060 130384 276072
rect 129976 276032 130384 276060
rect 129976 276020 129982 276032
rect 130378 276020 130384 276032
rect 130436 276020 130442 276072
rect 61838 274728 61844 274780
rect 61896 274768 61902 274780
rect 67634 274768 67640 274780
rect 61896 274740 67640 274768
rect 61896 274728 61902 274740
rect 67634 274728 67640 274740
rect 67692 274728 67698 274780
rect 52178 274660 52184 274712
rect 52236 274700 52242 274712
rect 67818 274700 67824 274712
rect 52236 274672 67824 274700
rect 52236 274660 52242 274672
rect 67818 274660 67824 274672
rect 67876 274660 67882 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 211798 274700 211804 274712
rect 121604 274672 211804 274700
rect 121604 274660 121610 274672
rect 211798 274660 211804 274672
rect 211856 274660 211862 274712
rect 39758 274592 39764 274644
rect 39816 274632 39822 274644
rect 67726 274632 67732 274644
rect 39816 274604 67732 274632
rect 39816 274592 39822 274604
rect 67726 274592 67732 274604
rect 67784 274592 67790 274644
rect 121638 274592 121644 274644
rect 121696 274632 121702 274644
rect 125778 274632 125784 274644
rect 121696 274604 125784 274632
rect 121696 274592 121702 274604
rect 125778 274592 125784 274604
rect 125836 274592 125842 274644
rect 121730 273912 121736 273964
rect 121788 273952 121794 273964
rect 287146 273952 287152 273964
rect 121788 273924 287152 273952
rect 121788 273912 121794 273924
rect 287146 273912 287152 273924
rect 287204 273912 287210 273964
rect 56502 273232 56508 273284
rect 56560 273272 56566 273284
rect 67634 273272 67640 273284
rect 56560 273244 67640 273272
rect 56560 273232 56566 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 121546 273232 121552 273284
rect 121604 273272 121610 273284
rect 210418 273272 210424 273284
rect 121604 273244 210424 273272
rect 121604 273232 121610 273244
rect 210418 273232 210424 273244
rect 210476 273232 210482 273284
rect 121638 273164 121644 273216
rect 121696 273204 121702 273216
rect 126974 273204 126980 273216
rect 121696 273176 126980 273204
rect 121696 273164 121702 273176
rect 126974 273164 126980 273176
rect 127032 273164 127038 273216
rect 66070 271872 66076 271924
rect 66128 271912 66134 271924
rect 67634 271912 67640 271924
rect 66128 271884 67640 271912
rect 66128 271872 66134 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 121546 271872 121552 271924
rect 121604 271912 121610 271924
rect 173894 271912 173900 271924
rect 121604 271884 173900 271912
rect 121604 271872 121610 271884
rect 173894 271872 173900 271884
rect 173952 271872 173958 271924
rect 54846 271804 54852 271856
rect 54904 271844 54910 271856
rect 67726 271844 67732 271856
rect 54904 271816 67732 271844
rect 54904 271804 54910 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 49510 270512 49516 270564
rect 49568 270552 49574 270564
rect 67634 270552 67640 270564
rect 49568 270524 67640 270552
rect 49568 270512 49574 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121546 270512 121552 270564
rect 121604 270552 121610 270564
rect 213270 270552 213276 270564
rect 121604 270524 213276 270552
rect 121604 270512 121610 270524
rect 213270 270512 213276 270524
rect 213328 270512 213334 270564
rect 121822 269764 121828 269816
rect 121880 269804 121886 269816
rect 471238 269804 471244 269816
rect 121880 269776 471244 269804
rect 121880 269764 121886 269776
rect 471238 269764 471244 269776
rect 471296 269764 471302 269816
rect 57514 269152 57520 269204
rect 57572 269192 57578 269204
rect 67726 269192 67732 269204
rect 57572 269164 67732 269192
rect 57572 269152 57578 269164
rect 67726 269152 67732 269164
rect 67784 269152 67790 269204
rect 121546 269152 121552 269204
rect 121604 269192 121610 269204
rect 237374 269192 237380 269204
rect 121604 269164 237380 269192
rect 121604 269152 121610 269164
rect 237374 269152 237380 269164
rect 237432 269152 237438 269204
rect 50890 269084 50896 269136
rect 50948 269124 50954 269136
rect 67634 269124 67640 269136
rect 50948 269096 67640 269124
rect 50948 269084 50954 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121638 269084 121644 269136
rect 121696 269124 121702 269136
rect 248414 269124 248420 269136
rect 121696 269096 248420 269124
rect 121696 269084 121702 269096
rect 248414 269084 248420 269096
rect 248472 269084 248478 269136
rect 121546 269016 121552 269068
rect 121604 269056 121610 269068
rect 146294 269056 146300 269068
rect 121604 269028 146300 269056
rect 121604 269016 121610 269028
rect 146294 269016 146300 269028
rect 146352 269016 146358 269068
rect 52270 268336 52276 268388
rect 52328 268376 52334 268388
rect 67634 268376 67640 268388
rect 52328 268348 67640 268376
rect 52328 268336 52334 268348
rect 67634 268336 67640 268348
rect 67692 268336 67698 268388
rect 51718 268200 51724 268252
rect 51776 268240 51782 268252
rect 52270 268240 52276 268252
rect 51776 268212 52276 268240
rect 51776 268200 51782 268212
rect 52270 268200 52276 268212
rect 52328 268200 52334 268252
rect 121546 267724 121552 267776
rect 121604 267764 121610 267776
rect 295334 267764 295340 267776
rect 121604 267736 295340 267764
rect 121604 267724 121610 267736
rect 295334 267724 295340 267736
rect 295392 267724 295398 267776
rect 41138 267656 41144 267708
rect 41196 267696 41202 267708
rect 67634 267696 67640 267708
rect 41196 267668 67640 267696
rect 41196 267656 41202 267668
rect 67634 267656 67640 267668
rect 67692 267656 67698 267708
rect 46842 267588 46848 267640
rect 46900 267628 46906 267640
rect 67726 267628 67732 267640
rect 46900 267600 67732 267628
rect 46900 267588 46906 267600
rect 67726 267588 67732 267600
rect 67784 267588 67790 267640
rect 121454 266432 121460 266484
rect 121512 266472 121518 266484
rect 280154 266472 280160 266484
rect 121512 266444 280160 266472
rect 121512 266432 121518 266444
rect 280154 266432 280160 266444
rect 280212 266432 280218 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 14458 266404 14464 266416
rect 3108 266376 14464 266404
rect 3108 266364 3114 266376
rect 14458 266364 14464 266376
rect 14516 266364 14522 266416
rect 121730 266364 121736 266416
rect 121788 266404 121794 266416
rect 309318 266404 309324 266416
rect 121788 266376 309324 266404
rect 121788 266364 121794 266376
rect 309318 266364 309324 266376
rect 309376 266364 309382 266416
rect 57606 266296 57612 266348
rect 57664 266336 57670 266348
rect 67634 266336 67640 266348
rect 57664 266308 67640 266336
rect 57664 266296 57670 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 216122 265044 216128 265056
rect 121512 265016 216128 265044
rect 121512 265004 121518 265016
rect 216122 265004 216128 265016
rect 216180 265004 216186 265056
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 310698 264976 310704 264988
rect 121604 264948 310704 264976
rect 121604 264936 121610 264948
rect 310698 264936 310704 264948
rect 310756 264936 310762 264988
rect 50706 264868 50712 264920
rect 50764 264908 50770 264920
rect 67634 264908 67640 264920
rect 50764 264880 67640 264908
rect 50764 264868 50770 264880
rect 67634 264868 67640 264880
rect 67692 264868 67698 264920
rect 121454 264868 121460 264920
rect 121512 264908 121518 264920
rect 133966 264908 133972 264920
rect 121512 264880 133972 264908
rect 121512 264868 121518 264880
rect 133966 264868 133972 264880
rect 134024 264868 134030 264920
rect 22738 264188 22744 264240
rect 22796 264228 22802 264240
rect 50706 264228 50712 264240
rect 22796 264200 50712 264228
rect 22796 264188 22802 264200
rect 50706 264188 50712 264200
rect 50764 264188 50770 264240
rect 48130 263576 48136 263628
rect 48188 263616 48194 263628
rect 67726 263616 67732 263628
rect 48188 263588 67732 263616
rect 48188 263576 48194 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 233234 263616 233240 263628
rect 121604 263588 233240 263616
rect 121604 263576 121610 263588
rect 233234 263576 233240 263588
rect 233292 263576 233298 263628
rect 61930 263508 61936 263560
rect 61988 263548 61994 263560
rect 67634 263548 67640 263560
rect 61988 263520 67640 263548
rect 61988 263508 61994 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 125594 263548 125600 263560
rect 121512 263520 125600 263548
rect 121512 263508 121518 263520
rect 125594 263508 125600 263520
rect 125652 263508 125658 263560
rect 56318 262216 56324 262268
rect 56376 262256 56382 262268
rect 67634 262256 67640 262268
rect 56376 262228 67640 262256
rect 56376 262216 56382 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 285674 262256 285680 262268
rect 121512 262228 285680 262256
rect 121512 262216 121518 262228
rect 285674 262216 285680 262228
rect 285732 262216 285738 262268
rect 121546 262148 121552 262200
rect 121604 262188 121610 262200
rect 132586 262188 132592 262200
rect 121604 262160 132592 262188
rect 121604 262148 121610 262160
rect 132586 262148 132592 262160
rect 132644 262148 132650 262200
rect 276658 261468 276664 261520
rect 276716 261508 276722 261520
rect 350534 261508 350540 261520
rect 276716 261480 350540 261508
rect 276716 261468 276722 261480
rect 350534 261468 350540 261480
rect 350592 261468 350598 261520
rect 61930 260924 61936 260976
rect 61988 260964 61994 260976
rect 67634 260964 67640 260976
rect 61988 260936 67640 260964
rect 61988 260924 61994 260936
rect 67634 260924 67640 260936
rect 67692 260924 67698 260976
rect 60274 260856 60280 260908
rect 60332 260896 60338 260908
rect 67726 260896 67732 260908
rect 60332 260868 67732 260896
rect 60332 260856 60338 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121730 260856 121736 260908
rect 121788 260896 121794 260908
rect 291838 260896 291844 260908
rect 121788 260868 291844 260896
rect 121788 260856 121794 260868
rect 291838 260856 291844 260868
rect 291896 260856 291902 260908
rect 60458 260788 60464 260840
rect 60516 260828 60522 260840
rect 67634 260828 67640 260840
rect 60516 260800 67640 260828
rect 60516 260788 60522 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 131666 260828 131672 260840
rect 121512 260800 131672 260828
rect 121512 260788 121518 260800
rect 131666 260788 131672 260800
rect 131724 260788 131730 260840
rect 131666 260108 131672 260160
rect 131724 260148 131730 260160
rect 353938 260148 353944 260160
rect 131724 260120 353944 260148
rect 131724 260108 131730 260120
rect 353938 260108 353944 260120
rect 353996 260108 354002 260160
rect 53650 259428 53656 259480
rect 53708 259468 53714 259480
rect 67634 259468 67640 259480
rect 53708 259440 67640 259468
rect 53708 259428 53714 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 207658 259468 207664 259480
rect 121512 259440 207664 259468
rect 121512 259428 121518 259440
rect 207658 259428 207664 259440
rect 207716 259428 207722 259480
rect 125410 259360 125416 259412
rect 125468 259400 125474 259412
rect 579798 259400 579804 259412
rect 125468 259372 579804 259400
rect 125468 259360 125474 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 121454 259292 121460 259344
rect 121512 259332 121518 259344
rect 127158 259332 127164 259344
rect 121512 259304 127164 259332
rect 121512 259292 121518 259304
rect 127158 259292 127164 259304
rect 127216 259292 127222 259344
rect 65978 258136 65984 258188
rect 66036 258176 66042 258188
rect 67634 258176 67640 258188
rect 66036 258148 67640 258176
rect 66036 258136 66042 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 58986 258068 58992 258120
rect 59044 258108 59050 258120
rect 67726 258108 67732 258120
rect 59044 258080 67732 258108
rect 59044 258068 59050 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121546 258068 121552 258120
rect 121604 258108 121610 258120
rect 288710 258108 288716 258120
rect 121604 258080 288716 258108
rect 121604 258068 121610 258080
rect 288710 258068 288716 258080
rect 288768 258068 288774 258120
rect 34514 258000 34520 258052
rect 34572 258040 34578 258052
rect 35802 258040 35808 258052
rect 34572 258012 35808 258040
rect 34572 258000 34578 258012
rect 35802 258000 35808 258012
rect 35860 258040 35866 258052
rect 67634 258040 67640 258052
rect 35860 258012 67640 258040
rect 35860 258000 35866 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 15838 257320 15844 257372
rect 15896 257360 15902 257372
rect 34514 257360 34520 257372
rect 15896 257332 34520 257360
rect 15896 257320 15902 257332
rect 34514 257320 34520 257332
rect 34572 257320 34578 257372
rect 233878 257320 233884 257372
rect 233936 257360 233942 257372
rect 296714 257360 296720 257372
rect 233936 257332 296720 257360
rect 233936 257320 233942 257332
rect 296714 257320 296720 257332
rect 296772 257320 296778 257372
rect 63218 256708 63224 256760
rect 63276 256748 63282 256760
rect 67634 256748 67640 256760
rect 63276 256720 67640 256748
rect 63276 256708 63282 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 242894 256748 242900 256760
rect 121604 256720 242900 256748
rect 121604 256708 121610 256720
rect 242894 256708 242900 256720
rect 242952 256708 242958 256760
rect 121454 256640 121460 256692
rect 121512 256680 121518 256692
rect 128538 256680 128544 256692
rect 121512 256652 128544 256680
rect 121512 256640 121518 256652
rect 128538 256640 128544 256652
rect 128596 256640 128602 256692
rect 54846 255280 54852 255332
rect 54904 255320 54910 255332
rect 67726 255320 67732 255332
rect 54904 255292 67732 255320
rect 54904 255280 54910 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 59262 255212 59268 255264
rect 59320 255252 59326 255264
rect 67634 255252 67640 255264
rect 59320 255224 67640 255252
rect 59320 255212 59326 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 125502 254532 125508 254584
rect 125560 254572 125566 254584
rect 580442 254572 580448 254584
rect 125560 254544 580448 254572
rect 125560 254532 125566 254544
rect 580442 254532 580448 254544
rect 580500 254532 580506 254584
rect 121546 254192 121552 254244
rect 121604 254232 121610 254244
rect 123478 254232 123484 254244
rect 121604 254204 123484 254232
rect 121604 254192 121610 254204
rect 123478 254192 123484 254204
rect 123536 254192 123542 254244
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 17310 253960 17316 253972
rect 3476 253932 17316 253960
rect 3476 253920 3482 253932
rect 17310 253920 17316 253932
rect 17368 253920 17374 253972
rect 60918 253920 60924 253972
rect 60976 253960 60982 253972
rect 67726 253960 67732 253972
rect 60976 253932 67732 253960
rect 60976 253920 60982 253932
rect 67726 253920 67732 253932
rect 67784 253920 67790 253972
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 235994 253960 236000 253972
rect 121512 253932 236000 253960
rect 121512 253920 121518 253932
rect 235994 253920 236000 253932
rect 236052 253920 236058 253972
rect 42794 253852 42800 253904
rect 42852 253892 42858 253904
rect 43806 253892 43812 253904
rect 42852 253864 43812 253892
rect 42852 253852 42858 253864
rect 43806 253852 43812 253864
rect 43864 253892 43870 253904
rect 67634 253892 67640 253904
rect 43864 253864 67640 253892
rect 43864 253852 43870 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 35158 253172 35164 253224
rect 35216 253212 35222 253224
rect 42794 253212 42800 253224
rect 35216 253184 42800 253212
rect 35216 253172 35222 253184
rect 42794 253172 42800 253184
rect 42852 253172 42858 253224
rect 63310 252560 63316 252612
rect 63368 252600 63374 252612
rect 67634 252600 67640 252612
rect 63368 252572 67640 252600
rect 63368 252560 63374 252572
rect 67634 252560 67640 252572
rect 67692 252560 67698 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 282270 252600 282276 252612
rect 121512 252572 282276 252600
rect 121512 252560 121518 252572
rect 282270 252560 282276 252572
rect 282328 252560 282334 252612
rect 121546 251812 121552 251864
rect 121604 251852 121610 251864
rect 231854 251852 231860 251864
rect 121604 251824 231860 251852
rect 121604 251812 121610 251824
rect 231854 251812 231860 251824
rect 231912 251812 231918 251864
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 276658 251240 276664 251252
rect 121512 251212 276664 251240
rect 121512 251200 121518 251212
rect 276658 251200 276664 251212
rect 276716 251200 276722 251252
rect 57790 249772 57796 249824
rect 57848 249812 57854 249824
rect 67726 249812 67732 249824
rect 57848 249784 67732 249812
rect 57848 249772 57854 249784
rect 67726 249772 67732 249784
rect 67784 249772 67790 249824
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 206462 249812 206468 249824
rect 121604 249784 206468 249812
rect 121604 249772 121610 249784
rect 206462 249772 206468 249784
rect 206520 249772 206526 249824
rect 39850 249704 39856 249756
rect 39908 249744 39914 249756
rect 67634 249744 67640 249756
rect 39908 249716 67640 249744
rect 39908 249704 39914 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121454 249704 121460 249756
rect 121512 249744 121518 249756
rect 131114 249744 131120 249756
rect 121512 249716 131120 249744
rect 121512 249704 121518 249716
rect 131114 249704 131120 249716
rect 131172 249704 131178 249756
rect 67450 248888 67456 248940
rect 67508 248928 67514 248940
rect 68830 248928 68836 248940
rect 67508 248900 68836 248928
rect 67508 248888 67514 248900
rect 68830 248888 68836 248900
rect 68888 248888 68894 248940
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 310606 248452 310612 248464
rect 121512 248424 310612 248452
rect 121512 248412 121518 248424
rect 310606 248412 310612 248424
rect 310664 248412 310670 248464
rect 130378 247664 130384 247716
rect 130436 247704 130442 247716
rect 580534 247704 580540 247716
rect 130436 247676 580540 247704
rect 130436 247664 130442 247676
rect 580534 247664 580540 247676
rect 580592 247664 580598 247716
rect 65886 247120 65892 247172
rect 65944 247160 65950 247172
rect 67634 247160 67640 247172
rect 65944 247132 67640 247160
rect 65944 247120 65950 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 59078 247052 59084 247104
rect 59136 247092 59142 247104
rect 67726 247092 67732 247104
rect 59136 247064 67732 247092
rect 59136 247052 59142 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 218698 247092 218704 247104
rect 121512 247064 218704 247092
rect 121512 247052 121518 247064
rect 218698 247052 218704 247064
rect 218756 247052 218762 247104
rect 54938 246984 54944 247036
rect 54996 247024 55002 247036
rect 67634 247024 67640 247036
rect 54996 246996 67640 247024
rect 54996 246984 55002 246996
rect 67634 246984 67640 246996
rect 67692 246984 67698 247036
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 237466 245664 237472 245676
rect 121512 245636 237472 245664
rect 121512 245624 121518 245636
rect 237466 245624 237472 245636
rect 237524 245624 237530 245676
rect 57698 245556 57704 245608
rect 57756 245596 57762 245608
rect 67634 245596 67640 245608
rect 57756 245568 67640 245596
rect 57756 245556 57762 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 64782 244944 64788 244996
rect 64840 244984 64846 244996
rect 68370 244984 68376 244996
rect 64840 244956 68376 244984
rect 64840 244944 64846 244956
rect 68370 244944 68376 244956
rect 68428 244944 68434 244996
rect 61654 244604 61660 244656
rect 61712 244644 61718 244656
rect 66898 244644 66904 244656
rect 61712 244616 66904 244644
rect 61712 244604 61718 244616
rect 66898 244604 66904 244616
rect 66956 244604 66962 244656
rect 67358 244332 67364 244384
rect 67416 244372 67422 244384
rect 68278 244372 68284 244384
rect 67416 244344 68284 244372
rect 67416 244332 67422 244344
rect 68278 244332 68284 244344
rect 68336 244332 68342 244384
rect 63126 244264 63132 244316
rect 63184 244304 63190 244316
rect 67634 244304 67640 244316
rect 63184 244276 67640 244304
rect 63184 244264 63190 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 306466 244304 306472 244316
rect 121604 244276 306472 244304
rect 121604 244264 121610 244276
rect 306466 244264 306472 244276
rect 306524 244264 306530 244316
rect 321646 244264 321652 244316
rect 321704 244304 321710 244316
rect 580166 244304 580172 244316
rect 321704 244276 580172 244304
rect 321704 244264 321710 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 49602 244196 49608 244248
rect 49660 244236 49666 244248
rect 67726 244236 67732 244248
rect 49660 244208 67732 244236
rect 49660 244196 49666 244208
rect 67726 244196 67732 244208
rect 67784 244196 67790 244248
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 125686 244236 125692 244248
rect 121512 244208 125692 244236
rect 121512 244196 121518 244208
rect 125686 244196 125692 244208
rect 125744 244196 125750 244248
rect 66162 242904 66168 242956
rect 66220 242944 66226 242956
rect 67818 242944 67824 242956
rect 66220 242916 67824 242944
rect 66220 242904 66226 242916
rect 67818 242904 67824 242916
rect 67876 242904 67882 242956
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 275278 242944 275284 242956
rect 121604 242916 275284 242944
rect 121604 242904 121610 242916
rect 275278 242904 275284 242916
rect 275336 242904 275342 242956
rect 62022 242836 62028 242888
rect 62080 242876 62086 242888
rect 67634 242876 67640 242888
rect 62080 242848 67640 242876
rect 62080 242836 62086 242848
rect 67634 242836 67640 242848
rect 67692 242836 67698 242888
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 142154 242876 142160 242888
rect 121512 242848 142160 242876
rect 121512 242836 121518 242848
rect 142154 242836 142160 242848
rect 142212 242876 142218 242888
rect 321646 242876 321652 242888
rect 142212 242848 321652 242876
rect 142212 242836 142218 242848
rect 321646 242836 321652 242848
rect 321704 242836 321710 242888
rect 121546 242768 121552 242820
rect 121604 242808 121610 242820
rect 129734 242808 129740 242820
rect 121604 242780 129740 242808
rect 121604 242768 121610 242780
rect 129734 242768 129740 242780
rect 129792 242768 129798 242820
rect 122098 241544 122104 241596
rect 122156 241584 122162 241596
rect 209130 241584 209136 241596
rect 122156 241556 209136 241584
rect 122156 241544 122162 241556
rect 209130 241544 209136 241556
rect 209188 241544 209194 241596
rect 60366 241476 60372 241528
rect 60424 241516 60430 241528
rect 67634 241516 67640 241528
rect 60424 241488 67640 241516
rect 60424 241476 60430 241488
rect 67634 241476 67640 241488
rect 67692 241476 67698 241528
rect 121454 241476 121460 241528
rect 121512 241516 121518 241528
rect 232038 241516 232044 241528
rect 121512 241488 232044 241516
rect 121512 241476 121518 241488
rect 232038 241476 232044 241488
rect 232096 241476 232102 241528
rect 3418 240116 3424 240168
rect 3476 240156 3482 240168
rect 3476 240128 11744 240156
rect 3476 240116 3482 240128
rect 11716 240088 11744 240128
rect 61746 240116 61752 240168
rect 61804 240156 61810 240168
rect 67634 240156 67640 240168
rect 61804 240128 67640 240156
rect 61804 240116 61810 240128
rect 67634 240116 67640 240128
rect 67692 240116 67698 240168
rect 119890 240116 119896 240168
rect 119948 240156 119954 240168
rect 288526 240156 288532 240168
rect 119948 240128 288532 240156
rect 119948 240116 119954 240128
rect 288526 240116 288532 240128
rect 288584 240116 288590 240168
rect 37090 240088 37096 240100
rect 11716 240060 37096 240088
rect 37090 240048 37096 240060
rect 37148 240048 37154 240100
rect 118970 239912 118976 239964
rect 119028 239952 119034 239964
rect 119982 239952 119988 239964
rect 119028 239924 119988 239952
rect 119028 239912 119034 239924
rect 119982 239912 119988 239924
rect 120040 239912 120046 239964
rect 70394 239776 70400 239828
rect 70452 239816 70458 239828
rect 71302 239816 71308 239828
rect 70452 239788 71308 239816
rect 70452 239776 70458 239788
rect 71302 239776 71308 239788
rect 71360 239776 71366 239828
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 78674 239776 78680 239828
rect 78732 239816 78738 239828
rect 79674 239816 79680 239828
rect 78732 239788 79680 239816
rect 78732 239776 78738 239788
rect 79674 239776 79680 239788
rect 79732 239776 79738 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 89714 239776 89720 239828
rect 89772 239816 89778 239828
rect 90622 239816 90628 239828
rect 89772 239788 90628 239816
rect 89772 239776 89778 239788
rect 90622 239776 90628 239788
rect 90680 239776 90686 239828
rect 93946 239776 93952 239828
rect 94004 239816 94010 239828
rect 95130 239816 95136 239828
rect 94004 239788 95136 239816
rect 94004 239776 94010 239788
rect 95130 239776 95136 239788
rect 95188 239776 95194 239828
rect 99374 239776 99380 239828
rect 99432 239816 99438 239828
rect 100282 239816 100288 239828
rect 99432 239788 100288 239816
rect 99432 239776 99438 239788
rect 100282 239776 100288 239788
rect 100340 239776 100346 239828
rect 100754 239776 100760 239828
rect 100812 239816 100818 239828
rect 101570 239816 101576 239828
rect 100812 239788 101576 239816
rect 100812 239776 100818 239788
rect 101570 239776 101576 239788
rect 101628 239776 101634 239828
rect 104894 239776 104900 239828
rect 104952 239816 104958 239828
rect 106078 239816 106084 239828
rect 104952 239788 106084 239816
rect 104952 239776 104958 239788
rect 106078 239776 106084 239788
rect 106136 239776 106142 239828
rect 107654 239776 107660 239828
rect 107712 239816 107718 239828
rect 108654 239816 108660 239828
rect 107712 239788 108660 239816
rect 107712 239776 107718 239788
rect 108654 239776 108660 239788
rect 108712 239776 108718 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 65978 239504 65984 239556
rect 66036 239544 66042 239556
rect 254026 239544 254032 239556
rect 66036 239516 254032 239544
rect 66036 239504 66042 239516
rect 254026 239504 254032 239516
rect 254084 239504 254090 239556
rect 63310 239436 63316 239488
rect 63368 239476 63374 239488
rect 272610 239476 272616 239488
rect 63368 239448 272616 239476
rect 63368 239436 63374 239448
rect 272610 239436 272616 239448
rect 272668 239436 272674 239488
rect 63218 239368 63224 239420
rect 63276 239408 63282 239420
rect 299474 239408 299480 239420
rect 63276 239380 299480 239408
rect 63276 239368 63282 239380
rect 299474 239368 299480 239380
rect 299532 239368 299538 239420
rect 84286 239300 84292 239352
rect 84344 239340 84350 239352
rect 85482 239340 85488 239352
rect 84344 239312 85488 239340
rect 84344 239300 84350 239312
rect 85482 239300 85488 239312
rect 85540 239300 85546 239352
rect 50982 238824 50988 238876
rect 51040 238864 51046 238876
rect 82262 238864 82268 238876
rect 51040 238836 82268 238864
rect 51040 238824 51046 238836
rect 82262 238824 82268 238836
rect 82320 238824 82326 238876
rect 103514 238824 103520 238876
rect 103572 238824 103578 238876
rect 115106 238824 115112 238876
rect 115164 238864 115170 238876
rect 132494 238864 132500 238876
rect 115164 238836 132500 238864
rect 115164 238824 115170 238836
rect 132494 238824 132500 238836
rect 132552 238824 132558 238876
rect 37090 238756 37096 238808
rect 37148 238796 37154 238808
rect 103532 238796 103560 238824
rect 37148 238768 103560 238796
rect 37148 238756 37154 238768
rect 106734 238756 106740 238808
rect 106792 238796 106798 238808
rect 139394 238796 139400 238808
rect 106792 238768 139400 238796
rect 106792 238756 106798 238768
rect 139394 238756 139400 238768
rect 139452 238756 139458 238808
rect 52362 238688 52368 238740
rect 52420 238728 52426 238740
rect 98362 238728 98368 238740
rect 52420 238700 98368 238728
rect 52420 238688 52426 238700
rect 98362 238688 98368 238700
rect 98420 238688 98426 238740
rect 118326 238688 118332 238740
rect 118384 238728 118390 238740
rect 123018 238728 123024 238740
rect 118384 238700 123024 238728
rect 118384 238688 118390 238700
rect 123018 238688 123024 238700
rect 123076 238688 123082 238740
rect 59170 238620 59176 238672
rect 59228 238660 59234 238672
rect 91922 238660 91928 238672
rect 59228 238632 91928 238660
rect 59228 238620 59234 238632
rect 91922 238620 91928 238632
rect 91980 238620 91986 238672
rect 53742 238552 53748 238604
rect 53800 238592 53806 238604
rect 95786 238592 95792 238604
rect 53800 238564 95792 238592
rect 53800 238552 53806 238564
rect 95786 238552 95792 238564
rect 95844 238552 95850 238604
rect 113818 238552 113824 238604
rect 113876 238592 113882 238604
rect 128722 238592 128728 238604
rect 113876 238564 128728 238592
rect 113876 238552 113882 238564
rect 128722 238552 128728 238564
rect 128780 238552 128786 238604
rect 60550 238484 60556 238536
rect 60608 238524 60614 238536
rect 72602 238524 72608 238536
rect 60608 238496 72608 238524
rect 60608 238484 60614 238496
rect 72602 238484 72608 238496
rect 72660 238484 72666 238536
rect 99006 238484 99012 238536
rect 99064 238524 99070 238536
rect 124214 238524 124220 238536
rect 99064 238496 124220 238524
rect 99064 238484 99070 238496
rect 124214 238484 124220 238496
rect 124272 238484 124278 238536
rect 89346 238416 89352 238468
rect 89404 238456 89410 238468
rect 133874 238456 133880 238468
rect 89404 238428 133880 238456
rect 89404 238416 89410 238428
rect 133874 238416 133880 238428
rect 133932 238416 133938 238468
rect 105446 238076 105452 238128
rect 105504 238116 105510 238128
rect 184198 238116 184204 238128
rect 105504 238088 184204 238116
rect 105504 238076 105510 238088
rect 184198 238076 184204 238088
rect 184256 238076 184262 238128
rect 96430 238008 96436 238060
rect 96488 238048 96494 238060
rect 276750 238048 276756 238060
rect 96488 238020 276756 238048
rect 96488 238008 96494 238020
rect 276750 238008 276756 238020
rect 276808 238008 276814 238060
rect 102870 237396 102876 237448
rect 102928 237436 102934 237448
rect 105538 237436 105544 237448
rect 102928 237408 105544 237436
rect 102928 237396 102934 237408
rect 105538 237396 105544 237408
rect 105596 237396 105602 237448
rect 48222 237328 48228 237380
rect 48280 237368 48286 237380
rect 107378 237368 107384 237380
rect 48280 237340 107384 237368
rect 48280 237328 48286 237340
rect 107378 237328 107384 237340
rect 107436 237328 107442 237380
rect 110598 237328 110604 237380
rect 110656 237368 110662 237380
rect 136634 237368 136640 237380
rect 110656 237340 136640 237368
rect 110656 237328 110662 237340
rect 136634 237328 136640 237340
rect 136692 237328 136698 237380
rect 14458 237260 14464 237312
rect 14516 237300 14522 237312
rect 14516 237272 45554 237300
rect 14516 237260 14522 237272
rect 45526 237232 45554 237272
rect 117038 237260 117044 237312
rect 117096 237300 117102 237312
rect 127066 237300 127072 237312
rect 117096 237272 127072 237300
rect 117096 237260 117102 237272
rect 127066 237260 127072 237272
rect 127124 237260 127130 237312
rect 57882 237232 57888 237244
rect 45526 237204 57888 237232
rect 57882 237192 57888 237204
rect 57940 237232 57946 237244
rect 86770 237232 86776 237244
rect 57940 237204 86776 237232
rect 57940 237192 57946 237204
rect 86770 237192 86776 237204
rect 86828 237192 86834 237244
rect 60642 237124 60648 237176
rect 60700 237164 60706 237176
rect 117682 237164 117688 237176
rect 60700 237136 117688 237164
rect 60700 237124 60706 237136
rect 117682 237124 117688 237136
rect 117740 237124 117746 237176
rect 110598 236784 110604 236836
rect 110656 236824 110662 236836
rect 111058 236824 111064 236836
rect 110656 236796 111064 236824
rect 110656 236784 110662 236796
rect 111058 236784 111064 236796
rect 111116 236784 111122 236836
rect 69290 236716 69296 236768
rect 69348 236756 69354 236768
rect 230474 236756 230480 236768
rect 69348 236728 230480 236756
rect 69348 236716 69354 236728
rect 230474 236716 230480 236728
rect 230532 236716 230538 236768
rect 282178 236716 282184 236768
rect 282236 236756 282242 236768
rect 331214 236756 331220 236768
rect 282236 236728 331220 236756
rect 282236 236716 282242 236728
rect 331214 236716 331220 236728
rect 331272 236716 331278 236768
rect 64782 236648 64788 236700
rect 64840 236688 64846 236700
rect 306558 236688 306564 236700
rect 64840 236660 306564 236688
rect 64840 236648 64846 236660
rect 306558 236648 306564 236660
rect 306616 236648 306622 236700
rect 17310 235900 17316 235952
rect 17368 235940 17374 235952
rect 34330 235940 34336 235952
rect 17368 235912 34336 235940
rect 17368 235900 17374 235912
rect 34330 235900 34336 235912
rect 34388 235940 34394 235952
rect 112530 235940 112536 235952
rect 34388 235912 112536 235940
rect 34388 235900 34394 235912
rect 112530 235900 112536 235912
rect 112588 235900 112594 235952
rect 114462 235900 114468 235952
rect 114520 235940 114526 235952
rect 124306 235940 124312 235952
rect 114520 235912 124312 235940
rect 114520 235900 114526 235912
rect 124306 235900 124312 235912
rect 124364 235900 124370 235952
rect 91278 235832 91284 235884
rect 91336 235872 91342 235884
rect 140866 235872 140872 235884
rect 91336 235844 140872 235872
rect 91336 235832 91342 235844
rect 140866 235832 140872 235844
rect 140924 235832 140930 235884
rect 117682 235220 117688 235272
rect 117740 235260 117746 235272
rect 177390 235260 177396 235272
rect 117740 235232 177396 235260
rect 117740 235220 117746 235232
rect 177390 235220 177396 235232
rect 177448 235220 177454 235272
rect 45462 234540 45468 234592
rect 45520 234580 45526 234592
rect 109034 234580 109040 234592
rect 45520 234552 109040 234580
rect 45520 234540 45526 234552
rect 109034 234540 109040 234552
rect 109092 234540 109098 234592
rect 81618 234472 81624 234524
rect 81676 234512 81682 234524
rect 135254 234512 135260 234524
rect 81676 234484 135260 234512
rect 81676 234472 81682 234484
rect 135254 234472 135260 234484
rect 135312 234472 135318 234524
rect 109034 234132 109040 234184
rect 109092 234172 109098 234184
rect 109954 234172 109960 234184
rect 109092 234144 109960 234172
rect 109092 234132 109098 234144
rect 109954 234132 109960 234144
rect 110012 234132 110018 234184
rect 74534 233928 74540 233980
rect 74592 233968 74598 233980
rect 75178 233968 75184 233980
rect 74592 233940 75184 233968
rect 74592 233928 74598 233940
rect 75178 233928 75184 233940
rect 75236 233928 75242 233980
rect 122374 233928 122380 233980
rect 122432 233968 122438 233980
rect 313366 233968 313372 233980
rect 122432 233940 313372 233968
rect 122432 233928 122438 233940
rect 313366 233928 313372 233940
rect 313424 233928 313430 233980
rect 66162 233860 66168 233912
rect 66220 233900 66226 233912
rect 276842 233900 276848 233912
rect 66220 233872 276848 233900
rect 66220 233860 66226 233872
rect 276842 233860 276848 233872
rect 276900 233860 276906 233912
rect 83458 233180 83464 233232
rect 83516 233220 83522 233232
rect 143534 233220 143540 233232
rect 83516 233192 143540 233220
rect 83516 233180 83522 233192
rect 143534 233180 143540 233192
rect 143592 233180 143598 233232
rect 92566 232500 92572 232552
rect 92624 232540 92630 232552
rect 238846 232540 238852 232552
rect 92624 232512 238852 232540
rect 92624 232500 92630 232512
rect 238846 232500 238852 232512
rect 238904 232500 238910 232552
rect 84102 231820 84108 231872
rect 84160 231860 84166 231872
rect 84838 231860 84844 231872
rect 84160 231832 84844 231860
rect 84160 231820 84166 231832
rect 84838 231820 84844 231832
rect 84896 231820 84902 231872
rect 94038 231072 94044 231124
rect 94096 231112 94102 231124
rect 271230 231112 271236 231124
rect 94096 231084 271236 231112
rect 94096 231072 94102 231084
rect 271230 231072 271236 231084
rect 271288 231072 271294 231124
rect 76006 230392 76012 230444
rect 76064 230432 76070 230444
rect 128354 230432 128360 230444
rect 76064 230404 128360 230432
rect 76064 230392 76070 230404
rect 128354 230392 128360 230404
rect 128412 230392 128418 230444
rect 128354 229780 128360 229832
rect 128412 229820 128418 229832
rect 187050 229820 187056 229832
rect 128412 229792 187056 229820
rect 128412 229780 128418 229792
rect 187050 229780 187056 229792
rect 187108 229780 187114 229832
rect 97626 229712 97632 229764
rect 97684 229752 97690 229764
rect 303798 229752 303804 229764
rect 97684 229724 303804 229752
rect 97684 229712 97690 229724
rect 303798 229712 303804 229724
rect 303856 229712 303862 229764
rect 78766 226992 78772 227044
rect 78824 227032 78830 227044
rect 231946 227032 231952 227044
rect 78824 227004 231952 227032
rect 78824 226992 78830 227004
rect 231946 226992 231952 227004
rect 232004 226992 232010 227044
rect 82814 226244 82820 226296
rect 82872 226284 82878 226296
rect 133874 226284 133880 226296
rect 82872 226256 133880 226284
rect 82872 226244 82878 226256
rect 133874 226244 133880 226256
rect 133932 226284 133938 226296
rect 135162 226284 135168 226296
rect 133932 226256 135168 226284
rect 133932 226244 133938 226256
rect 135162 226244 135168 226256
rect 135220 226244 135226 226296
rect 135162 224952 135168 225004
rect 135220 224992 135226 225004
rect 358078 224992 358084 225004
rect 135220 224964 358084 224992
rect 135220 224952 135226 224964
rect 358078 224952 358084 224964
rect 358136 224952 358142 225004
rect 71866 224204 71872 224256
rect 71924 224244 71930 224256
rect 268378 224244 268384 224256
rect 71924 224216 268384 224244
rect 71924 224204 71930 224216
rect 268378 224204 268384 224216
rect 268436 224204 268442 224256
rect 61838 222844 61844 222896
rect 61896 222884 61902 222896
rect 244274 222884 244280 222896
rect 61896 222856 244280 222884
rect 61896 222844 61902 222856
rect 244274 222844 244280 222856
rect 244332 222844 244338 222896
rect 53558 220124 53564 220176
rect 53616 220164 53622 220176
rect 142798 220164 142804 220176
rect 53616 220136 142804 220164
rect 53616 220124 53622 220136
rect 142798 220124 142804 220136
rect 142856 220124 142862 220176
rect 103606 220056 103612 220108
rect 103664 220096 103670 220108
rect 287238 220096 287244 220108
rect 103664 220068 287244 220096
rect 103664 220056 103670 220068
rect 287238 220056 287244 220068
rect 287296 220056 287302 220108
rect 60366 218696 60372 218748
rect 60424 218736 60430 218748
rect 247034 218736 247040 218748
rect 60424 218708 247040 218736
rect 60424 218696 60430 218708
rect 247034 218696 247040 218708
rect 247092 218696 247098 218748
rect 74626 217336 74632 217388
rect 74684 217376 74690 217388
rect 265618 217376 265624 217388
rect 74684 217348 265624 217376
rect 74684 217336 74690 217348
rect 265618 217336 265624 217348
rect 265676 217336 265682 217388
rect 57514 217268 57520 217320
rect 57572 217308 57578 217320
rect 252554 217308 252560 217320
rect 57572 217280 252560 217308
rect 57572 217268 57578 217280
rect 252554 217268 252560 217280
rect 252612 217268 252618 217320
rect 231118 216044 231124 216096
rect 231176 216084 231182 216096
rect 245654 216084 245660 216096
rect 231176 216056 245660 216084
rect 231176 216044 231182 216056
rect 245654 216044 245660 216056
rect 245712 216044 245718 216096
rect 88334 215976 88340 216028
rect 88392 216016 88398 216028
rect 285950 216016 285956 216028
rect 88392 215988 285956 216016
rect 88392 215976 88398 215988
rect 285950 215976 285956 215988
rect 286008 215976 286014 216028
rect 73246 215908 73252 215960
rect 73304 215948 73310 215960
rect 273990 215948 273996 215960
rect 73304 215920 273996 215948
rect 73304 215908 73310 215920
rect 273990 215908 273996 215920
rect 274048 215908 274054 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 22738 215268 22744 215280
rect 3384 215240 22744 215268
rect 3384 215228 3390 215240
rect 22738 215228 22744 215240
rect 22796 215228 22802 215280
rect 50890 214548 50896 214600
rect 50948 214588 50954 214600
rect 295426 214588 295432 214600
rect 50948 214560 295432 214588
rect 50948 214548 50954 214560
rect 295426 214548 295432 214560
rect 295484 214548 295490 214600
rect 61746 213256 61752 213308
rect 61804 213296 61810 213308
rect 261478 213296 261484 213308
rect 61804 213268 261484 213296
rect 61804 213256 61810 213268
rect 261478 213256 261484 213268
rect 261536 213256 261542 213308
rect 48130 213188 48136 213240
rect 48188 213228 48194 213240
rect 305086 213228 305092 213240
rect 48188 213200 305092 213228
rect 48188 213188 48194 213200
rect 305086 213188 305092 213200
rect 305144 213188 305150 213240
rect 123478 211828 123484 211880
rect 123536 211868 123542 211880
rect 255958 211868 255964 211880
rect 123536 211840 255964 211868
rect 123536 211828 123542 211840
rect 255958 211828 255964 211840
rect 256016 211828 256022 211880
rect 77386 211760 77392 211812
rect 77444 211800 77450 211812
rect 233326 211800 233332 211812
rect 77444 211772 233332 211800
rect 77444 211760 77450 211772
rect 233326 211760 233332 211772
rect 233384 211760 233390 211812
rect 46750 210400 46756 210452
rect 46808 210440 46814 210452
rect 302418 210440 302424 210452
rect 46808 210412 302424 210440
rect 46808 210400 46814 210412
rect 302418 210400 302424 210412
rect 302476 210400 302482 210452
rect 89806 209040 89812 209092
rect 89864 209080 89870 209092
rect 233418 209080 233424 209092
rect 89864 209052 233424 209080
rect 89864 209040 89870 209052
rect 233418 209040 233424 209052
rect 233476 209040 233482 209092
rect 55030 207748 55036 207800
rect 55088 207788 55094 207800
rect 213362 207788 213368 207800
rect 55088 207760 213368 207788
rect 55088 207748 55094 207760
rect 213362 207748 213368 207760
rect 213420 207748 213426 207800
rect 104894 207680 104900 207732
rect 104952 207720 104958 207732
rect 284386 207720 284392 207732
rect 104952 207692 284392 207720
rect 104952 207680 104958 207692
rect 284386 207680 284392 207692
rect 284444 207680 284450 207732
rect 56318 207612 56324 207664
rect 56376 207652 56382 207664
rect 241514 207652 241520 207664
rect 56376 207624 241520 207652
rect 56376 207612 56382 207624
rect 241514 207612 241520 207624
rect 241572 207612 241578 207664
rect 100846 206388 100852 206440
rect 100904 206428 100910 206440
rect 232130 206428 232136 206440
rect 100904 206400 232136 206428
rect 100904 206388 100910 206400
rect 232130 206388 232136 206400
rect 232188 206388 232194 206440
rect 69106 206320 69112 206372
rect 69164 206360 69170 206372
rect 230566 206360 230572 206372
rect 69164 206332 230572 206360
rect 69164 206320 69170 206332
rect 230566 206320 230572 206332
rect 230624 206320 230630 206372
rect 102134 206252 102140 206304
rect 102192 206292 102198 206304
rect 289906 206292 289912 206304
rect 102192 206264 289912 206292
rect 102192 206252 102198 206264
rect 289906 206252 289912 206264
rect 289964 206252 289970 206304
rect 163498 205028 163504 205080
rect 163556 205068 163562 205080
rect 264330 205068 264336 205080
rect 163556 205040 264336 205068
rect 163556 205028 163562 205040
rect 264330 205028 264336 205040
rect 264388 205028 264394 205080
rect 105538 204960 105544 205012
rect 105596 205000 105602 205012
rect 220170 205000 220176 205012
rect 105596 204972 220176 205000
rect 105596 204960 105602 204972
rect 220170 204960 220176 204972
rect 220228 204960 220234 205012
rect 52086 204892 52092 204944
rect 52144 204932 52150 204944
rect 269942 204932 269948 204944
rect 52144 204904 269948 204932
rect 52144 204892 52150 204904
rect 269942 204892 269948 204904
rect 270000 204892 270006 204944
rect 93946 203600 93952 203652
rect 94004 203640 94010 203652
rect 258810 203640 258816 203652
rect 94004 203612 258816 203640
rect 94004 203600 94010 203612
rect 258810 203600 258816 203612
rect 258868 203600 258874 203652
rect 14458 203532 14464 203584
rect 14516 203572 14522 203584
rect 83458 203572 83464 203584
rect 14516 203544 83464 203572
rect 14516 203532 14522 203544
rect 83458 203532 83464 203544
rect 83516 203532 83522 203584
rect 113174 203532 113180 203584
rect 113232 203572 113238 203584
rect 306650 203572 306656 203584
rect 113232 203544 306656 203572
rect 113232 203532 113238 203544
rect 306650 203532 306656 203544
rect 306708 203532 306714 203584
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 120074 202824 120080 202836
rect 3476 202796 120080 202824
rect 3476 202784 3482 202796
rect 120074 202784 120080 202796
rect 120132 202784 120138 202836
rect 100754 202172 100760 202224
rect 100812 202212 100818 202224
rect 234798 202212 234804 202224
rect 100812 202184 234804 202212
rect 100812 202172 100818 202184
rect 234798 202172 234804 202184
rect 234856 202172 234862 202224
rect 151078 202104 151084 202156
rect 151136 202144 151142 202156
rect 305178 202144 305184 202156
rect 151136 202116 305184 202144
rect 151136 202104 151142 202116
rect 305178 202104 305184 202116
rect 305236 202104 305242 202156
rect 133138 200812 133144 200864
rect 133196 200852 133202 200864
rect 240226 200852 240232 200864
rect 133196 200824 240232 200852
rect 133196 200812 133202 200824
rect 240226 200812 240232 200824
rect 240284 200812 240290 200864
rect 152458 200744 152464 200796
rect 152516 200784 152522 200796
rect 303890 200784 303896 200796
rect 152516 200756 303896 200784
rect 152516 200744 152522 200756
rect 303890 200744 303896 200756
rect 303948 200744 303954 200796
rect 96614 199656 96620 199708
rect 96672 199696 96678 199708
rect 218790 199696 218796 199708
rect 96672 199668 218796 199696
rect 96672 199656 96678 199668
rect 218790 199656 218796 199668
rect 218848 199656 218854 199708
rect 166350 199588 166356 199640
rect 166408 199628 166414 199640
rect 291194 199628 291200 199640
rect 166408 199600 291200 199628
rect 166408 199588 166414 199600
rect 291194 199588 291200 199600
rect 291252 199588 291258 199640
rect 93854 199520 93860 199572
rect 93912 199560 93918 199572
rect 234890 199560 234896 199572
rect 93912 199532 234896 199560
rect 93912 199520 93918 199532
rect 234890 199520 234896 199532
rect 234948 199520 234954 199572
rect 280798 199520 280804 199572
rect 280856 199560 280862 199572
rect 300946 199560 300952 199572
rect 280856 199532 300952 199560
rect 280856 199520 280862 199532
rect 300946 199520 300952 199532
rect 301004 199520 301010 199572
rect 107746 199452 107752 199504
rect 107804 199492 107810 199504
rect 299658 199492 299664 199504
rect 107804 199464 299664 199492
rect 107804 199452 107810 199464
rect 299658 199452 299664 199464
rect 299716 199452 299722 199504
rect 52178 199384 52184 199436
rect 52236 199424 52242 199436
rect 296898 199424 296904 199436
rect 52236 199396 296904 199424
rect 52236 199384 52242 199396
rect 296898 199384 296904 199396
rect 296956 199384 296962 199436
rect 157978 198024 157984 198076
rect 158036 198064 158042 198076
rect 294046 198064 294052 198076
rect 158036 198036 294052 198064
rect 158036 198024 158042 198036
rect 294046 198024 294052 198036
rect 294104 198024 294110 198076
rect 73154 197956 73160 198008
rect 73212 197996 73218 198008
rect 275370 197996 275376 198008
rect 73212 197968 275376 197996
rect 73212 197956 73218 197968
rect 275370 197956 275376 197968
rect 275428 197956 275434 198008
rect 67542 196732 67548 196784
rect 67600 196772 67606 196784
rect 230658 196772 230664 196784
rect 67600 196744 230664 196772
rect 67600 196732 67606 196744
rect 230658 196732 230664 196744
rect 230716 196732 230722 196784
rect 92474 196664 92480 196716
rect 92532 196704 92538 196716
rect 285858 196704 285864 196716
rect 92532 196676 285864 196704
rect 92532 196664 92538 196676
rect 285858 196664 285864 196676
rect 285916 196664 285922 196716
rect 86218 196596 86224 196648
rect 86276 196636 86282 196648
rect 582558 196636 582564 196648
rect 86276 196608 582564 196636
rect 86276 196596 86282 196608
rect 582558 196596 582564 196608
rect 582616 196596 582622 196648
rect 84286 195372 84292 195424
rect 84344 195412 84350 195424
rect 233510 195412 233516 195424
rect 84344 195384 233516 195412
rect 84344 195372 84350 195384
rect 233510 195372 233516 195384
rect 233568 195372 233574 195424
rect 107654 195304 107660 195356
rect 107712 195344 107718 195356
rect 285766 195344 285772 195356
rect 107712 195316 285772 195344
rect 107712 195304 107718 195316
rect 285766 195304 285772 195316
rect 285824 195304 285830 195356
rect 70486 195236 70492 195288
rect 70544 195276 70550 195288
rect 276934 195276 276940 195288
rect 70544 195248 276940 195276
rect 70544 195236 70550 195248
rect 276934 195236 276940 195248
rect 276992 195236 276998 195288
rect 145558 194080 145564 194132
rect 145616 194120 145622 194132
rect 196710 194120 196716 194132
rect 145616 194092 196716 194120
rect 145616 194080 145622 194092
rect 196710 194080 196716 194092
rect 196768 194080 196774 194132
rect 110414 194012 110420 194064
rect 110472 194052 110478 194064
rect 236086 194052 236092 194064
rect 110472 194024 236092 194052
rect 110472 194012 110478 194024
rect 236086 194012 236092 194024
rect 236144 194012 236150 194064
rect 50798 193944 50804 193996
rect 50856 193984 50862 193996
rect 244366 193984 244372 193996
rect 50856 193956 244372 193984
rect 50856 193944 50862 193956
rect 244366 193944 244372 193956
rect 244424 193944 244430 193996
rect 56502 193876 56508 193928
rect 56560 193916 56566 193928
rect 260834 193916 260840 193928
rect 56560 193888 260840 193916
rect 56560 193876 56566 193888
rect 260834 193876 260840 193888
rect 260892 193876 260898 193928
rect 54846 193808 54852 193860
rect 54904 193848 54910 193860
rect 296990 193848 296996 193860
rect 54904 193820 296996 193848
rect 54904 193808 54910 193820
rect 296990 193808 296996 193820
rect 297048 193808 297054 193860
rect 352558 193128 352564 193180
rect 352616 193168 352622 193180
rect 580166 193168 580172 193180
rect 352616 193140 580172 193168
rect 352616 193128 352622 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 142798 192516 142804 192568
rect 142856 192556 142862 192568
rect 242986 192556 242992 192568
rect 142856 192528 242992 192556
rect 142856 192516 142862 192528
rect 242986 192516 242992 192528
rect 243044 192516 243050 192568
rect 61930 192448 61936 192500
rect 61988 192488 61994 192500
rect 294138 192488 294144 192500
rect 61988 192460 294144 192488
rect 61988 192448 61994 192460
rect 294138 192448 294144 192460
rect 294196 192448 294202 192500
rect 103514 191292 103520 191344
rect 103572 191332 103578 191344
rect 180242 191332 180248 191344
rect 103572 191304 180248 191332
rect 103572 191292 103578 191304
rect 180242 191292 180248 191304
rect 180300 191292 180306 191344
rect 111794 191224 111800 191276
rect 111852 191264 111858 191276
rect 251358 191264 251364 191276
rect 111852 191236 251364 191264
rect 111852 191224 111858 191236
rect 251358 191224 251364 191236
rect 251416 191224 251422 191276
rect 114554 191156 114560 191208
rect 114612 191196 114618 191208
rect 280246 191196 280252 191208
rect 114612 191168 280252 191196
rect 114612 191156 114618 191168
rect 280246 191156 280252 191168
rect 280304 191156 280310 191208
rect 70394 191088 70400 191140
rect 70452 191128 70458 191140
rect 247126 191128 247132 191140
rect 70452 191100 247132 191128
rect 70452 191088 70458 191100
rect 247126 191088 247132 191100
rect 247184 191088 247190 191140
rect 214650 189728 214656 189780
rect 214708 189768 214714 189780
rect 292758 189768 292764 189780
rect 214708 189740 292764 189768
rect 214708 189728 214714 189740
rect 292758 189728 292764 189740
rect 292816 189728 292822 189780
rect 105538 189048 105544 189100
rect 105596 189088 105602 189100
rect 214742 189088 214748 189100
rect 105596 189060 214748 189088
rect 105596 189048 105602 189060
rect 214742 189048 214748 189060
rect 214800 189048 214806 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 17218 189020 17224 189032
rect 3476 188992 17224 189020
rect 3476 188980 3482 188992
rect 17218 188980 17224 188992
rect 17276 188980 17282 189032
rect 192478 188436 192484 188488
rect 192536 188476 192542 188488
rect 302510 188476 302516 188488
rect 192536 188448 302516 188476
rect 192536 188436 192542 188448
rect 302510 188436 302516 188448
rect 302568 188436 302574 188488
rect 89714 188368 89720 188420
rect 89772 188408 89778 188420
rect 241606 188408 241612 188420
rect 89772 188380 241612 188408
rect 89772 188368 89778 188380
rect 241606 188368 241612 188380
rect 241664 188368 241670 188420
rect 99374 188300 99380 188352
rect 99432 188340 99438 188352
rect 252646 188340 252652 188352
rect 99432 188312 252652 188340
rect 99432 188300 99438 188312
rect 252646 188300 252652 188312
rect 252704 188300 252710 188352
rect 101950 187756 101956 187808
rect 102008 187796 102014 187808
rect 171870 187796 171876 187808
rect 102008 187768 171876 187796
rect 102008 187756 102014 187768
rect 171870 187756 171876 187768
rect 171928 187756 171934 187808
rect 104802 187688 104808 187740
rect 104860 187728 104866 187740
rect 184290 187728 184296 187740
rect 104860 187700 184296 187728
rect 104860 187688 104866 187700
rect 184290 187688 184296 187700
rect 184348 187688 184354 187740
rect 224310 187008 224316 187060
rect 224368 187048 224374 187060
rect 298278 187048 298284 187060
rect 224368 187020 298284 187048
rect 224368 187008 224374 187020
rect 298278 187008 298284 187020
rect 298336 187008 298342 187060
rect 155218 186940 155224 186992
rect 155276 186980 155282 186992
rect 295518 186980 295524 186992
rect 155276 186952 295524 186980
rect 155276 186940 155282 186952
rect 295518 186940 295524 186952
rect 295576 186940 295582 186992
rect 128262 186396 128268 186448
rect 128320 186436 128326 186448
rect 171962 186436 171968 186448
rect 128320 186408 171968 186436
rect 128320 186396 128326 186408
rect 171962 186396 171968 186408
rect 172020 186396 172026 186448
rect 99282 186328 99288 186380
rect 99340 186368 99346 186380
rect 214650 186368 214656 186380
rect 99340 186340 214656 186368
rect 99340 186328 99346 186340
rect 214650 186328 214656 186340
rect 214708 186328 214714 186380
rect 40678 185784 40684 185836
rect 40736 185824 40742 185836
rect 109034 185824 109040 185836
rect 40736 185796 109040 185824
rect 40736 185784 40742 185796
rect 109034 185784 109040 185796
rect 109092 185784 109098 185836
rect 61654 185716 61660 185768
rect 61712 185756 61718 185768
rect 244550 185756 244556 185768
rect 61712 185728 244556 185756
rect 61712 185716 61718 185728
rect 244550 185716 244556 185728
rect 244608 185716 244614 185768
rect 58986 185648 58992 185700
rect 59044 185688 59050 185700
rect 249794 185688 249800 185700
rect 59044 185660 249800 185688
rect 59044 185648 59050 185660
rect 249794 185648 249800 185660
rect 249852 185648 249858 185700
rect 282270 185648 282276 185700
rect 282328 185688 282334 185700
rect 308030 185688 308036 185700
rect 282328 185660 308036 185688
rect 282328 185648 282334 185660
rect 308030 185648 308036 185660
rect 308088 185648 308094 185700
rect 84194 185580 84200 185632
rect 84252 185620 84258 185632
rect 283006 185620 283012 185632
rect 84252 185592 283012 185620
rect 84252 185580 84258 185592
rect 283006 185580 283012 185592
rect 283064 185580 283070 185632
rect 119982 184968 119988 185020
rect 120040 185008 120046 185020
rect 170490 185008 170496 185020
rect 120040 184980 170496 185008
rect 120040 184968 120046 184980
rect 170490 184968 170496 184980
rect 170548 184968 170554 185020
rect 114462 184900 114468 184952
rect 114520 184940 114526 184952
rect 213454 184940 213460 184952
rect 114520 184912 213460 184940
rect 114520 184900 114526 184912
rect 213454 184900 213460 184912
rect 213512 184900 213518 184952
rect 115934 184288 115940 184340
rect 115992 184328 115998 184340
rect 248598 184328 248604 184340
rect 115992 184300 248604 184328
rect 115992 184288 115998 184300
rect 248598 184288 248604 184300
rect 248656 184288 248662 184340
rect 271230 184288 271236 184340
rect 271288 184328 271294 184340
rect 299566 184328 299572 184340
rect 271288 184300 299572 184328
rect 271288 184288 271294 184300
rect 299566 184288 299572 184300
rect 299624 184288 299630 184340
rect 80146 184220 80152 184272
rect 80204 184260 80210 184272
rect 284478 184260 284484 184272
rect 80204 184232 284484 184260
rect 80204 184220 80210 184232
rect 284478 184220 284484 184232
rect 284536 184220 284542 184272
rect 69014 184152 69020 184204
rect 69072 184192 69078 184204
rect 281534 184192 281540 184204
rect 69072 184164 281540 184192
rect 69072 184152 69078 184164
rect 281534 184152 281540 184164
rect 281592 184152 281598 184204
rect 100662 183540 100668 183592
rect 100720 183580 100726 183592
rect 167638 183580 167644 183592
rect 100720 183552 167644 183580
rect 100720 183540 100726 183552
rect 167638 183540 167644 183552
rect 167696 183540 167702 183592
rect 159358 183064 159364 183116
rect 159416 183104 159422 183116
rect 198090 183104 198096 183116
rect 159416 183076 198096 183104
rect 159416 183064 159422 183076
rect 198090 183064 198096 183076
rect 198148 183064 198154 183116
rect 180150 182996 180156 183048
rect 180208 183036 180214 183048
rect 227714 183036 227720 183048
rect 180208 183008 227720 183036
rect 180208 182996 180214 183008
rect 227714 182996 227720 183008
rect 227772 182996 227778 183048
rect 65886 182928 65892 182980
rect 65944 182968 65950 182980
rect 251266 182968 251272 182980
rect 65944 182940 251272 182968
rect 65944 182928 65950 182940
rect 251266 182928 251272 182940
rect 251324 182928 251330 182980
rect 59078 182860 59084 182912
rect 59136 182900 59142 182912
rect 245838 182900 245844 182912
rect 59136 182872 245844 182900
rect 59136 182860 59142 182872
rect 245838 182860 245844 182872
rect 245896 182860 245902 182912
rect 80054 182792 80060 182844
rect 80112 182832 80118 182844
rect 280430 182832 280436 182844
rect 80112 182804 280436 182832
rect 80112 182792 80118 182804
rect 280430 182792 280436 182804
rect 280488 182792 280494 182844
rect 264330 182724 264336 182776
rect 264388 182764 264394 182776
rect 269114 182764 269120 182776
rect 264388 182736 269120 182764
rect 264388 182724 264394 182736
rect 269114 182724 269120 182736
rect 269172 182724 269178 182776
rect 118418 182248 118424 182300
rect 118476 182288 118482 182300
rect 166350 182288 166356 182300
rect 118476 182260 166356 182288
rect 118476 182248 118482 182260
rect 166350 182248 166356 182260
rect 166408 182248 166414 182300
rect 97718 182180 97724 182232
rect 97776 182220 97782 182232
rect 169110 182220 169116 182232
rect 97776 182192 169116 182220
rect 97776 182180 97782 182192
rect 169110 182180 169116 182192
rect 169168 182180 169174 182232
rect 278130 181772 278136 181824
rect 278188 181812 278194 181824
rect 301038 181812 301044 181824
rect 278188 181784 301044 181812
rect 278188 181772 278194 181784
rect 301038 181772 301044 181784
rect 301096 181772 301102 181824
rect 213270 181704 213276 181756
rect 213328 181744 213334 181756
rect 240134 181744 240140 181756
rect 213328 181716 240140 181744
rect 213328 181704 213334 181716
rect 240134 181704 240140 181716
rect 240192 181704 240198 181756
rect 261478 181704 261484 181756
rect 261536 181744 261542 181756
rect 292574 181744 292580 181756
rect 261536 181716 292580 181744
rect 261536 181704 261542 181716
rect 292574 181704 292580 181716
rect 292632 181704 292638 181756
rect 198182 181636 198188 181688
rect 198240 181676 198246 181688
rect 256786 181676 256792 181688
rect 198240 181648 256792 181676
rect 198240 181636 198246 181648
rect 256786 181636 256792 181648
rect 256844 181636 256850 181688
rect 269758 181636 269764 181688
rect 269816 181676 269822 181688
rect 307754 181676 307760 181688
rect 269816 181648 307760 181676
rect 269816 181636 269822 181648
rect 307754 181636 307760 181648
rect 307812 181636 307818 181688
rect 86954 181568 86960 181620
rect 87012 181608 87018 181620
rect 236178 181608 236184 181620
rect 87012 181580 236184 181608
rect 87012 181568 87018 181580
rect 236178 181568 236184 181580
rect 236236 181568 236242 181620
rect 264238 181568 264244 181620
rect 264296 181608 264302 181620
rect 335354 181608 335360 181620
rect 264296 181580 335360 181608
rect 264296 181568 264302 181580
rect 335354 181568 335360 181580
rect 335412 181568 335418 181620
rect 53650 181500 53656 181552
rect 53708 181540 53714 181552
rect 291470 181540 291476 181552
rect 53708 181512 291476 181540
rect 53708 181500 53714 181512
rect 291470 181500 291476 181512
rect 291528 181500 291534 181552
rect 60274 181432 60280 181484
rect 60332 181472 60338 181484
rect 301130 181472 301136 181484
rect 60332 181444 301136 181472
rect 60332 181432 60338 181444
rect 301130 181432 301136 181444
rect 301188 181432 301194 181484
rect 129458 180956 129464 181008
rect 129516 180996 129522 181008
rect 166442 180996 166448 181008
rect 129516 180968 166448 180996
rect 129516 180956 129522 180968
rect 166442 180956 166448 180968
rect 166500 180956 166506 181008
rect 122650 180888 122656 180940
rect 122708 180928 122714 180940
rect 167914 180928 167920 180940
rect 122708 180900 167920 180928
rect 122708 180888 122714 180900
rect 167914 180888 167920 180900
rect 167972 180888 167978 180940
rect 114094 180820 114100 180872
rect 114152 180860 114158 180872
rect 169202 180860 169208 180872
rect 114152 180832 169208 180860
rect 114152 180820 114158 180832
rect 169202 180820 169208 180832
rect 169260 180820 169266 180872
rect 226978 180412 226984 180464
rect 227036 180452 227042 180464
rect 248506 180452 248512 180464
rect 227036 180424 248512 180452
rect 227036 180412 227042 180424
rect 248506 180412 248512 180424
rect 248564 180412 248570 180464
rect 213362 180344 213368 180396
rect 213420 180384 213426 180396
rect 241698 180384 241704 180396
rect 213420 180356 241704 180384
rect 213420 180344 213426 180356
rect 241698 180344 241704 180356
rect 241756 180344 241762 180396
rect 166258 180276 166264 180328
rect 166316 180316 166322 180328
rect 199470 180316 199476 180328
rect 166316 180288 199476 180316
rect 166316 180276 166322 180288
rect 199470 180276 199476 180288
rect 199528 180276 199534 180328
rect 204990 180276 204996 180328
rect 205048 180316 205054 180328
rect 238754 180316 238760 180328
rect 205048 180288 238760 180316
rect 205048 180276 205054 180288
rect 238754 180276 238760 180288
rect 238812 180276 238818 180328
rect 273898 180276 273904 180328
rect 273956 180316 273962 180328
rect 288434 180316 288440 180328
rect 273956 180288 288440 180316
rect 273956 180276 273962 180288
rect 288434 180276 288440 180288
rect 288492 180276 288498 180328
rect 162118 180208 162124 180260
rect 162176 180248 162182 180260
rect 206370 180248 206376 180260
rect 162176 180220 206376 180248
rect 162176 180208 162182 180220
rect 206370 180208 206376 180220
rect 206428 180208 206434 180260
rect 207658 180208 207664 180260
rect 207716 180248 207722 180260
rect 258074 180248 258080 180260
rect 207716 180220 258080 180248
rect 207716 180208 207722 180220
rect 258074 180208 258080 180220
rect 258132 180208 258138 180260
rect 271138 180208 271144 180260
rect 271196 180248 271202 180260
rect 299750 180248 299756 180260
rect 271196 180220 299756 180248
rect 271196 180208 271202 180220
rect 299750 180208 299756 180220
rect 299808 180208 299814 180260
rect 182818 180140 182824 180192
rect 182876 180180 182882 180192
rect 244458 180180 244464 180192
rect 182876 180152 244464 180180
rect 182876 180140 182882 180152
rect 244458 180140 244464 180152
rect 244516 180140 244522 180192
rect 258810 180140 258816 180192
rect 258868 180180 258874 180192
rect 296806 180180 296812 180192
rect 258868 180152 296812 180180
rect 258868 180140 258874 180152
rect 296806 180140 296812 180152
rect 296864 180140 296870 180192
rect 69198 180072 69204 180124
rect 69256 180112 69262 180124
rect 280338 180112 280344 180124
rect 69256 180084 280344 180112
rect 69256 180072 69262 180084
rect 280338 180072 280344 180084
rect 280396 180072 280402 180124
rect 133138 179460 133144 179512
rect 133196 179500 133202 179512
rect 165062 179500 165068 179512
rect 133196 179472 165068 179500
rect 133196 179460 133202 179472
rect 165062 179460 165068 179472
rect 165120 179460 165126 179512
rect 126790 179392 126796 179444
rect 126848 179432 126854 179444
rect 166534 179432 166540 179444
rect 126848 179404 166540 179432
rect 126848 179392 126854 179404
rect 166534 179392 166540 179404
rect 166592 179392 166598 179444
rect 272518 179324 272524 179376
rect 272576 179364 272582 179376
rect 279326 179364 279332 179376
rect 272576 179336 279332 179364
rect 272576 179324 272582 179336
rect 279326 179324 279332 179336
rect 279384 179324 279390 179376
rect 211798 178984 211804 179036
rect 211856 179024 211862 179036
rect 245746 179024 245752 179036
rect 211856 178996 245752 179024
rect 211856 178984 211862 178996
rect 245746 178984 245752 178996
rect 245804 178984 245810 179036
rect 203518 178916 203524 178968
rect 203576 178956 203582 178968
rect 243078 178956 243084 178968
rect 203576 178928 243084 178956
rect 203576 178916 203582 178928
rect 243078 178916 243084 178928
rect 243136 178916 243142 178968
rect 178770 178848 178776 178900
rect 178828 178888 178834 178900
rect 238938 178888 238944 178900
rect 178828 178860 238944 178888
rect 178828 178848 178834 178860
rect 238938 178848 238944 178860
rect 238996 178848 239002 178900
rect 169018 178780 169024 178832
rect 169076 178820 169082 178832
rect 240318 178820 240324 178832
rect 169076 178792 240324 178820
rect 169076 178780 169082 178792
rect 240318 178780 240324 178792
rect 240376 178780 240382 178832
rect 269850 178780 269856 178832
rect 269908 178820 269914 178832
rect 278774 178820 278780 178832
rect 269908 178792 278780 178820
rect 269908 178780 269914 178792
rect 278774 178780 278780 178792
rect 278832 178780 278838 178832
rect 220078 178712 220084 178764
rect 220136 178752 220142 178764
rect 299382 178752 299388 178764
rect 220136 178724 299388 178752
rect 220136 178712 220142 178724
rect 299382 178712 299388 178724
rect 299440 178712 299446 178764
rect 214558 178644 214564 178696
rect 214616 178684 214622 178696
rect 340966 178684 340972 178696
rect 214616 178656 340972 178684
rect 214616 178644 214622 178656
rect 340966 178644 340972 178656
rect 341024 178644 341030 178696
rect 134794 178372 134800 178424
rect 134852 178412 134858 178424
rect 165522 178412 165528 178424
rect 134852 178384 165528 178412
rect 134852 178372 134858 178384
rect 165522 178372 165528 178384
rect 165580 178372 165586 178424
rect 132402 178304 132408 178356
rect 132460 178344 132466 178356
rect 165430 178344 165436 178356
rect 132460 178316 165436 178344
rect 132460 178304 132466 178316
rect 165430 178304 165436 178316
rect 165488 178304 165494 178356
rect 123754 178236 123760 178288
rect 123812 178276 123818 178288
rect 169294 178276 169300 178288
rect 123812 178248 169300 178276
rect 123812 178236 123818 178248
rect 169294 178236 169300 178248
rect 169352 178236 169358 178288
rect 115842 178168 115848 178220
rect 115900 178208 115906 178220
rect 167822 178208 167828 178220
rect 115900 178180 167828 178208
rect 115900 178168 115906 178180
rect 167822 178168 167828 178180
rect 167880 178168 167886 178220
rect 148226 178100 148232 178152
rect 148284 178140 148290 178152
rect 210510 178140 210516 178152
rect 148284 178112 210516 178140
rect 148284 178100 148290 178112
rect 210510 178100 210516 178112
rect 210568 178100 210574 178152
rect 130746 178032 130752 178084
rect 130804 178072 130810 178084
rect 214098 178072 214104 178084
rect 130804 178044 214104 178072
rect 130804 178032 130810 178044
rect 214098 178032 214104 178044
rect 214156 178032 214162 178084
rect 298738 178032 298744 178084
rect 298796 178072 298802 178084
rect 299474 178072 299480 178084
rect 298796 178044 299480 178072
rect 298796 178032 298802 178044
rect 299474 178032 299480 178044
rect 299532 178032 299538 178084
rect 222838 177964 222844 178016
rect 222896 178004 222902 178016
rect 229370 178004 229376 178016
rect 222896 177976 229376 178004
rect 222896 177964 222902 177976
rect 229370 177964 229376 177976
rect 229428 177964 229434 178016
rect 102042 177828 102048 177880
rect 102100 177868 102106 177880
rect 105538 177868 105544 177880
rect 102100 177840 105544 177868
rect 102100 177828 102106 177840
rect 105538 177828 105544 177840
rect 105596 177828 105602 177880
rect 276750 177624 276756 177676
rect 276808 177664 276814 177676
rect 287054 177664 287060 177676
rect 276808 177636 287060 177664
rect 276808 177624 276814 177636
rect 287054 177624 287060 177636
rect 287112 177624 287118 177676
rect 276934 177556 276940 177608
rect 276992 177596 276998 177608
rect 288618 177596 288624 177608
rect 276992 177568 288624 177596
rect 276992 177556 276998 177568
rect 288618 177556 288624 177568
rect 288676 177556 288682 177608
rect 221458 177488 221464 177540
rect 221516 177528 221522 177540
rect 229094 177528 229100 177540
rect 221516 177500 229100 177528
rect 221516 177488 221522 177500
rect 229094 177488 229100 177500
rect 229152 177488 229158 177540
rect 272610 177488 272616 177540
rect 272668 177528 272674 177540
rect 284294 177528 284300 177540
rect 272668 177500 284300 177528
rect 272668 177488 272674 177500
rect 284294 177488 284300 177500
rect 284352 177488 284358 177540
rect 220170 177420 220176 177472
rect 220228 177460 220234 177472
rect 237650 177460 237656 177472
rect 220228 177432 237656 177460
rect 220228 177420 220234 177432
rect 237650 177420 237656 177432
rect 237708 177420 237714 177472
rect 276658 177420 276664 177472
rect 276716 177460 276722 177472
rect 291378 177460 291384 177472
rect 276716 177432 291384 177460
rect 276716 177420 276722 177432
rect 291378 177420 291384 177432
rect 291436 177420 291442 177472
rect 218790 177352 218796 177404
rect 218848 177392 218854 177404
rect 237558 177392 237564 177404
rect 218848 177364 237564 177392
rect 218848 177352 218854 177364
rect 237558 177352 237564 177364
rect 237616 177352 237622 177404
rect 268378 177352 268384 177404
rect 268436 177392 268442 177404
rect 292666 177392 292672 177404
rect 268436 177364 292672 177392
rect 268436 177352 268442 177364
rect 292666 177352 292672 177364
rect 292724 177352 292730 177404
rect 227162 177284 227168 177336
rect 227220 177324 227226 177336
rect 247218 177324 247224 177336
rect 227220 177296 247224 177324
rect 227220 177284 227226 177296
rect 247218 177284 247224 177296
rect 247276 177284 247282 177336
rect 255958 177284 255964 177336
rect 256016 177324 256022 177336
rect 290090 177324 290096 177336
rect 256016 177296 290096 177324
rect 256016 177284 256022 177296
rect 290090 177284 290096 177296
rect 290148 177284 290154 177336
rect 291838 177148 291844 177200
rect 291896 177188 291902 177200
rect 295610 177188 295616 177200
rect 291896 177160 295616 177188
rect 291896 177148 291902 177160
rect 295610 177148 295616 177160
rect 295668 177148 295674 177200
rect 128170 177012 128176 177064
rect 128228 177052 128234 177064
rect 169754 177052 169760 177064
rect 128228 177024 169760 177052
rect 128228 177012 128234 177024
rect 169754 177012 169760 177024
rect 169812 177012 169818 177064
rect 107010 176944 107016 176996
rect 107068 176984 107074 176996
rect 164418 176984 164424 176996
rect 107068 176956 164424 176984
rect 107068 176944 107074 176956
rect 164418 176944 164424 176956
rect 164476 176944 164482 176996
rect 105722 176876 105728 176928
rect 105780 176916 105786 176928
rect 169018 176916 169024 176928
rect 105780 176888 169024 176916
rect 105780 176876 105786 176888
rect 169018 176876 169024 176888
rect 169076 176876 169082 176928
rect 103330 176808 103336 176860
rect 103388 176848 103394 176860
rect 167730 176848 167736 176860
rect 103388 176820 167736 176848
rect 103388 176808 103394 176820
rect 167730 176808 167736 176820
rect 167788 176808 167794 176860
rect 136082 176740 136088 176792
rect 136140 176780 136146 176792
rect 213822 176780 213828 176792
rect 136140 176752 213828 176780
rect 136140 176740 136146 176752
rect 213822 176740 213828 176752
rect 213880 176740 213886 176792
rect 108114 176672 108120 176724
rect 108172 176712 108178 176724
rect 188430 176712 188436 176724
rect 108172 176684 188436 176712
rect 108172 176672 108178 176684
rect 188430 176672 188436 176684
rect 188488 176672 188494 176724
rect 158898 176264 158904 176316
rect 158956 176304 158962 176316
rect 166258 176304 166264 176316
rect 158956 176276 166264 176304
rect 158956 176264 158962 176276
rect 166258 176264 166264 176276
rect 166316 176264 166322 176316
rect 164418 176196 164424 176248
rect 164476 176236 164482 176248
rect 214558 176236 214564 176248
rect 164476 176208 214564 176236
rect 164476 176196 164482 176208
rect 214558 176196 214564 176208
rect 214616 176196 214622 176248
rect 110690 176128 110696 176180
rect 110748 176168 110754 176180
rect 170582 176168 170588 176180
rect 110748 176140 170588 176168
rect 110748 176128 110754 176140
rect 170582 176128 170588 176140
rect 170640 176128 170646 176180
rect 210418 176128 210424 176180
rect 210476 176168 210482 176180
rect 229186 176168 229192 176180
rect 210476 176140 229192 176168
rect 210476 176128 210482 176140
rect 229186 176128 229192 176140
rect 229244 176128 229250 176180
rect 275370 176128 275376 176180
rect 275428 176168 275434 176180
rect 281626 176168 281632 176180
rect 275428 176140 281632 176168
rect 275428 176128 275434 176140
rect 281626 176128 281632 176140
rect 281684 176128 281690 176180
rect 124490 176060 124496 176112
rect 124548 176100 124554 176112
rect 211798 176100 211804 176112
rect 124548 176072 211804 176100
rect 124548 176060 124554 176072
rect 211798 176060 211804 176072
rect 211856 176060 211862 176112
rect 218698 176060 218704 176112
rect 218756 176100 218762 176112
rect 229278 176100 229284 176112
rect 218756 176072 229284 176100
rect 218756 176060 218762 176072
rect 229278 176060 229284 176072
rect 229336 176060 229342 176112
rect 276842 176060 276848 176112
rect 276900 176100 276906 176112
rect 289814 176100 289820 176112
rect 276900 176072 289820 176100
rect 276900 176060 276906 176072
rect 289814 176060 289820 176072
rect 289872 176060 289878 176112
rect 120810 175992 120816 176044
rect 120868 176032 120874 176044
rect 210602 176032 210608 176044
rect 120868 176004 210608 176032
rect 120868 175992 120874 176004
rect 210602 175992 210608 176004
rect 210660 175992 210666 176044
rect 225598 175992 225604 176044
rect 225656 176032 225662 176044
rect 243170 176032 243176 176044
rect 225656 176004 243176 176032
rect 225656 175992 225662 176004
rect 243170 175992 243176 176004
rect 243228 175992 243234 176044
rect 273990 175992 273996 176044
rect 274048 176032 274054 176044
rect 289998 176032 290004 176044
rect 274048 176004 290004 176032
rect 274048 175992 274054 176004
rect 289998 175992 290004 176004
rect 290056 175992 290062 176044
rect 290458 175992 290464 176044
rect 290516 176032 290522 176044
rect 292850 176032 292856 176044
rect 290516 176004 292856 176032
rect 290516 175992 290522 176004
rect 292850 175992 292856 176004
rect 292908 175992 292914 176044
rect 11698 175924 11704 175976
rect 11756 175964 11762 175976
rect 111058 175964 111064 175976
rect 11756 175936 111064 175964
rect 11756 175924 11762 175936
rect 111058 175924 111064 175936
rect 111116 175924 111122 175976
rect 116946 175924 116952 175976
rect 117004 175964 117010 175976
rect 213270 175964 213276 175976
rect 117004 175936 213276 175964
rect 117004 175924 117010 175936
rect 213270 175924 213276 175936
rect 213328 175924 213334 175976
rect 224218 175924 224224 175976
rect 224276 175964 224282 175976
rect 251450 175964 251456 175976
rect 224276 175936 251456 175964
rect 224276 175924 224282 175936
rect 251450 175924 251456 175936
rect 251508 175924 251514 175976
rect 275278 175924 275284 175976
rect 275336 175964 275342 175976
rect 294230 175964 294236 175976
rect 275336 175936 294236 175964
rect 275336 175924 275342 175936
rect 294230 175924 294236 175936
rect 294288 175924 294294 175976
rect 165062 175176 165068 175228
rect 165120 175216 165126 175228
rect 214006 175216 214012 175228
rect 165120 175188 214012 175216
rect 165120 175176 165126 175188
rect 214006 175176 214012 175188
rect 214064 175176 214070 175228
rect 236638 175176 236644 175228
rect 236696 175216 236702 175228
rect 237374 175216 237380 175228
rect 236696 175188 237380 175216
rect 236696 175176 236702 175188
rect 237374 175176 237380 175188
rect 237432 175176 237438 175228
rect 165522 175108 165528 175160
rect 165580 175148 165586 175160
rect 213914 175148 213920 175160
rect 165580 175120 213920 175148
rect 165580 175108 165586 175120
rect 213914 175108 213920 175120
rect 213972 175108 213978 175160
rect 254578 173952 254584 174004
rect 254636 173992 254642 174004
rect 265802 173992 265808 174004
rect 254636 173964 265808 173992
rect 254636 173952 254642 173964
rect 265802 173952 265808 173964
rect 265860 173952 265866 174004
rect 242526 173884 242532 173936
rect 242584 173924 242590 173936
rect 264422 173924 264428 173936
rect 242584 173896 264428 173924
rect 242584 173884 242590 173896
rect 264422 173884 264428 173896
rect 264480 173884 264486 173936
rect 165430 173816 165436 173868
rect 165488 173856 165494 173868
rect 213914 173856 213920 173868
rect 165488 173828 213920 173856
rect 165488 173816 165494 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231762 173816 231768 173868
rect 231820 173856 231826 173868
rect 242986 173856 242992 173868
rect 231820 173828 242992 173856
rect 231820 173816 231826 173828
rect 242986 173816 242992 173828
rect 243044 173816 243050 173868
rect 231118 173748 231124 173800
rect 231176 173788 231182 173800
rect 240226 173788 240232 173800
rect 231176 173760 240232 173788
rect 231176 173748 231182 173760
rect 240226 173748 240232 173760
rect 240284 173748 240290 173800
rect 231486 173680 231492 173732
rect 231544 173720 231550 173732
rect 238754 173720 238760 173732
rect 231544 173692 238760 173720
rect 231544 173680 231550 173692
rect 238754 173680 238760 173692
rect 238812 173680 238818 173732
rect 243722 173136 243728 173188
rect 243780 173176 243786 173188
rect 265710 173176 265716 173188
rect 243780 173148 265716 173176
rect 243780 173136 243786 173148
rect 265710 173136 265716 173148
rect 265768 173136 265774 173188
rect 262858 172592 262864 172644
rect 262916 172632 262922 172644
rect 265526 172632 265532 172644
rect 262916 172604 265532 172632
rect 262916 172592 262922 172604
rect 265526 172592 265532 172604
rect 265584 172592 265590 172644
rect 238110 172524 238116 172576
rect 238168 172564 238174 172576
rect 265894 172564 265900 172576
rect 238168 172536 265900 172564
rect 238168 172524 238174 172536
rect 265894 172524 265900 172536
rect 265952 172524 265958 172576
rect 166442 172456 166448 172508
rect 166500 172496 166506 172508
rect 213914 172496 213920 172508
rect 166500 172468 213920 172496
rect 166500 172456 166506 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 231762 172456 231768 172508
rect 231820 172496 231826 172508
rect 240134 172496 240140 172508
rect 231820 172468 240140 172496
rect 231820 172456 231826 172468
rect 240134 172456 240140 172468
rect 240192 172456 240198 172508
rect 169754 172388 169760 172440
rect 169812 172428 169818 172440
rect 214006 172428 214012 172440
rect 169812 172400 214012 172428
rect 169812 172388 169818 172400
rect 214006 172388 214012 172400
rect 214064 172388 214070 172440
rect 282086 171776 282092 171828
rect 282144 171816 282150 171828
rect 287054 171816 287060 171828
rect 282144 171788 287060 171816
rect 282144 171776 282150 171788
rect 287054 171776 287060 171788
rect 287112 171776 287118 171828
rect 167546 171300 167552 171352
rect 167604 171340 167610 171352
rect 170674 171340 170680 171352
rect 167604 171312 170680 171340
rect 167604 171300 167610 171312
rect 170674 171300 170680 171312
rect 170732 171300 170738 171352
rect 257338 171232 257344 171284
rect 257396 171272 257402 171284
rect 265618 171272 265624 171284
rect 257396 171244 265624 171272
rect 257396 171232 257402 171244
rect 265618 171232 265624 171244
rect 265676 171232 265682 171284
rect 246390 171164 246396 171216
rect 246448 171204 246454 171216
rect 265802 171204 265808 171216
rect 246448 171176 265808 171204
rect 246448 171164 246454 171176
rect 265802 171164 265808 171176
rect 265860 171164 265866 171216
rect 241146 171096 241152 171148
rect 241204 171136 241210 171148
rect 265894 171136 265900 171148
rect 241204 171108 265900 171136
rect 241204 171096 241210 171108
rect 265894 171096 265900 171108
rect 265952 171096 265958 171148
rect 166534 171028 166540 171080
rect 166592 171068 166598 171080
rect 214006 171068 214012 171080
rect 166592 171040 214012 171068
rect 166592 171028 166598 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 245654 171068 245660 171080
rect 231820 171040 245660 171068
rect 231820 171028 231826 171040
rect 245654 171028 245660 171040
rect 245712 171028 245718 171080
rect 171962 170960 171968 171012
rect 172020 171000 172026 171012
rect 215110 171000 215116 171012
rect 172020 170972 215116 171000
rect 172020 170960 172026 170972
rect 215110 170960 215116 170972
rect 215168 170960 215174 171012
rect 231118 170960 231124 171012
rect 231176 171000 231182 171012
rect 245838 171000 245844 171012
rect 231176 170972 245844 171000
rect 231176 170960 231182 170972
rect 245838 170960 245844 170972
rect 245896 170960 245902 171012
rect 231486 170892 231492 170944
rect 231544 170932 231550 170944
rect 244274 170932 244280 170944
rect 231544 170904 244280 170932
rect 231544 170892 231550 170904
rect 244274 170892 244280 170904
rect 244332 170892 244338 170944
rect 229738 170416 229744 170468
rect 229796 170456 229802 170468
rect 239030 170456 239036 170468
rect 229796 170428 239036 170456
rect 229796 170416 229802 170428
rect 239030 170416 239036 170428
rect 239088 170416 239094 170468
rect 229830 170348 229836 170400
rect 229888 170388 229894 170400
rect 241606 170388 241612 170400
rect 229888 170360 241612 170388
rect 229888 170348 229894 170360
rect 241606 170348 241612 170360
rect 241664 170348 241670 170400
rect 258902 169872 258908 169924
rect 258960 169912 258966 169924
rect 265250 169912 265256 169924
rect 258960 169884 265256 169912
rect 258960 169872 258966 169884
rect 265250 169872 265256 169884
rect 265308 169872 265314 169924
rect 282270 169872 282276 169924
rect 282328 169912 282334 169924
rect 288434 169912 288440 169924
rect 282328 169884 288440 169912
rect 282328 169872 282334 169884
rect 288434 169872 288440 169884
rect 288492 169872 288498 169924
rect 244918 169804 244924 169856
rect 244976 169844 244982 169856
rect 265434 169844 265440 169856
rect 244976 169816 265440 169844
rect 244976 169804 244982 169816
rect 265434 169804 265440 169816
rect 265492 169804 265498 169856
rect 239674 169736 239680 169788
rect 239732 169776 239738 169788
rect 265618 169776 265624 169788
rect 239732 169748 265624 169776
rect 239732 169736 239738 169748
rect 265618 169736 265624 169748
rect 265676 169736 265682 169788
rect 281718 169736 281724 169788
rect 281776 169776 281782 169788
rect 284294 169776 284300 169788
rect 281776 169748 284300 169776
rect 281776 169736 281782 169748
rect 284294 169736 284300 169748
rect 284352 169736 284358 169788
rect 169294 169668 169300 169720
rect 169352 169708 169358 169720
rect 213914 169708 213920 169720
rect 169352 169680 213920 169708
rect 169352 169668 169358 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 231486 169668 231492 169720
rect 231544 169708 231550 169720
rect 237558 169708 237564 169720
rect 231544 169680 237564 169708
rect 231544 169668 231550 169680
rect 237558 169668 237564 169680
rect 237616 169668 237622 169720
rect 282822 169668 282828 169720
rect 282880 169708 282886 169720
rect 301130 169708 301136 169720
rect 282880 169680 301136 169708
rect 282880 169668 282886 169680
rect 301130 169668 301136 169680
rect 301188 169668 301194 169720
rect 211798 169600 211804 169652
rect 211856 169640 211862 169652
rect 214006 169640 214012 169652
rect 211856 169612 214012 169640
rect 211856 169600 211862 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 230750 169532 230756 169584
rect 230808 169572 230814 169584
rect 237650 169572 237656 169584
rect 230808 169544 237656 169572
rect 230808 169532 230814 169544
rect 237650 169532 237656 169544
rect 237708 169532 237714 169584
rect 256234 168512 256240 168564
rect 256292 168552 256298 168564
rect 265342 168552 265348 168564
rect 256292 168524 265348 168552
rect 256292 168512 256298 168524
rect 265342 168512 265348 168524
rect 265400 168512 265406 168564
rect 242434 168444 242440 168496
rect 242492 168484 242498 168496
rect 265802 168484 265808 168496
rect 242492 168456 265808 168484
rect 242492 168444 242498 168456
rect 265802 168444 265808 168456
rect 265860 168444 265866 168496
rect 239766 168376 239772 168428
rect 239824 168416 239830 168428
rect 265618 168416 265624 168428
rect 239824 168388 265624 168416
rect 239824 168376 239830 168388
rect 265618 168376 265624 168388
rect 265676 168376 265682 168428
rect 167914 168308 167920 168360
rect 167972 168348 167978 168360
rect 213914 168348 213920 168360
rect 167972 168320 213920 168348
rect 167972 168308 167978 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 238938 168348 238944 168360
rect 231820 168320 238944 168348
rect 231820 168308 231826 168320
rect 238938 168308 238944 168320
rect 238996 168308 239002 168360
rect 282454 168308 282460 168360
rect 282512 168348 282518 168360
rect 289814 168348 289820 168360
rect 282512 168320 289820 168348
rect 282512 168308 282518 168320
rect 289814 168308 289820 168320
rect 289872 168308 289878 168360
rect 210602 168240 210608 168292
rect 210660 168280 210666 168292
rect 214006 168280 214012 168292
rect 210660 168252 214012 168280
rect 210660 168240 210666 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 232498 167628 232504 167680
rect 232556 167668 232562 167680
rect 243078 167668 243084 167680
rect 232556 167640 243084 167668
rect 232556 167628 232562 167640
rect 243078 167628 243084 167640
rect 243136 167628 243142 167680
rect 250530 167084 250536 167136
rect 250588 167124 250594 167136
rect 265342 167124 265348 167136
rect 250588 167096 265348 167124
rect 250588 167084 250594 167096
rect 265342 167084 265348 167096
rect 265400 167084 265406 167136
rect 243630 167016 243636 167068
rect 243688 167056 243694 167068
rect 264422 167056 264428 167068
rect 243688 167028 264428 167056
rect 243688 167016 243694 167028
rect 264422 167016 264428 167028
rect 264480 167016 264486 167068
rect 231670 166948 231676 167000
rect 231728 166988 231734 167000
rect 241514 166988 241520 167000
rect 231728 166960 241520 166988
rect 231728 166948 231734 166960
rect 241514 166948 241520 166960
rect 241572 166948 241578 167000
rect 282086 166948 282092 167000
rect 282144 166988 282150 167000
rect 295426 166988 295432 167000
rect 282144 166960 295432 166988
rect 282144 166948 282150 166960
rect 295426 166948 295432 166960
rect 295484 166948 295490 167000
rect 353938 166948 353944 167000
rect 353996 166988 354002 167000
rect 580166 166988 580172 167000
rect 353996 166960 580172 166988
rect 353996 166948 354002 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 170490 166880 170496 166932
rect 170548 166920 170554 166932
rect 213914 166920 213920 166932
rect 170548 166892 213920 166920
rect 170548 166880 170554 166892
rect 213914 166880 213920 166892
rect 213972 166880 213978 166932
rect 231762 166880 231768 166932
rect 231820 166920 231826 166932
rect 238846 166920 238852 166932
rect 231820 166892 238852 166920
rect 231820 166880 231826 166892
rect 238846 166880 238852 166892
rect 238904 166880 238910 166932
rect 166350 166812 166356 166864
rect 166408 166852 166414 166864
rect 214006 166852 214012 166864
rect 166408 166824 214012 166852
rect 166408 166812 166414 166824
rect 214006 166812 214012 166824
rect 214064 166812 214070 166864
rect 282638 166268 282644 166320
rect 282696 166308 282702 166320
rect 294138 166308 294144 166320
rect 282696 166280 294144 166308
rect 282696 166268 282702 166280
rect 294138 166268 294144 166280
rect 294196 166268 294202 166320
rect 253474 165724 253480 165776
rect 253532 165764 253538 165776
rect 265802 165764 265808 165776
rect 253532 165736 265808 165764
rect 253532 165724 253538 165736
rect 265802 165724 265808 165736
rect 265860 165724 265866 165776
rect 246298 165656 246304 165708
rect 246356 165696 246362 165708
rect 265710 165696 265716 165708
rect 246356 165668 265716 165696
rect 246356 165656 246362 165668
rect 265710 165656 265716 165668
rect 265768 165656 265774 165708
rect 238294 165588 238300 165640
rect 238352 165628 238358 165640
rect 265342 165628 265348 165640
rect 238352 165600 265348 165628
rect 238352 165588 238358 165600
rect 265342 165588 265348 165600
rect 265400 165588 265406 165640
rect 167822 165520 167828 165572
rect 167880 165560 167886 165572
rect 213914 165560 213920 165572
rect 167880 165532 213920 165560
rect 167880 165520 167886 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 231118 165520 231124 165572
rect 231176 165560 231182 165572
rect 233418 165560 233424 165572
rect 231176 165532 233424 165560
rect 231176 165520 231182 165532
rect 233418 165520 233424 165532
rect 233476 165520 233482 165572
rect 282086 165520 282092 165572
rect 282144 165560 282150 165572
rect 289906 165560 289912 165572
rect 282144 165532 289912 165560
rect 282144 165520 282150 165532
rect 289906 165520 289912 165532
rect 289964 165520 289970 165572
rect 231670 165452 231676 165504
rect 231728 165492 231734 165504
rect 241698 165492 241704 165504
rect 231728 165464 241704 165492
rect 231728 165452 231734 165464
rect 241698 165452 241704 165464
rect 241756 165452 241762 165504
rect 231762 165384 231768 165436
rect 231820 165424 231826 165436
rect 243170 165424 243176 165436
rect 231820 165396 243176 165424
rect 231820 165384 231826 165396
rect 243170 165384 243176 165396
rect 243228 165384 243234 165436
rect 249058 164840 249064 164892
rect 249116 164880 249122 164892
rect 265250 164880 265256 164892
rect 249116 164852 265256 164880
rect 249116 164840 249122 164852
rect 265250 164840 265256 164852
rect 265308 164840 265314 164892
rect 255958 164296 255964 164348
rect 256016 164336 256022 164348
rect 265158 164336 265164 164348
rect 256016 164308 265164 164336
rect 256016 164296 256022 164308
rect 265158 164296 265164 164308
rect 265216 164296 265222 164348
rect 240778 164228 240784 164280
rect 240836 164268 240842 164280
rect 265342 164268 265348 164280
rect 240836 164240 265348 164268
rect 240836 164228 240842 164240
rect 265342 164228 265348 164240
rect 265400 164228 265406 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 25498 164200 25504 164212
rect 3292 164172 25504 164200
rect 3292 164160 3298 164172
rect 25498 164160 25504 164172
rect 25556 164160 25562 164212
rect 169202 164160 169208 164212
rect 169260 164200 169266 164212
rect 213914 164200 213920 164212
rect 169260 164172 213920 164200
rect 169260 164160 169266 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 231118 164160 231124 164212
rect 231176 164200 231182 164212
rect 233234 164200 233240 164212
rect 231176 164172 233240 164200
rect 231176 164160 231182 164172
rect 233234 164160 233240 164172
rect 233292 164160 233298 164212
rect 282822 164160 282828 164212
rect 282880 164200 282886 164212
rect 291470 164200 291476 164212
rect 282880 164172 291476 164200
rect 282880 164160 282886 164172
rect 291470 164160 291476 164172
rect 291528 164160 291534 164212
rect 231762 164092 231768 164144
rect 231820 164132 231826 164144
rect 240410 164132 240416 164144
rect 231820 164104 240416 164132
rect 231820 164092 231826 164104
rect 240410 164092 240416 164104
rect 240468 164092 240474 164144
rect 231670 164024 231676 164076
rect 231728 164064 231734 164076
rect 244550 164064 244556 164076
rect 231728 164036 244556 164064
rect 231728 164024 231734 164036
rect 244550 164024 244556 164036
rect 244608 164024 244614 164076
rect 242158 163480 242164 163532
rect 242216 163520 242222 163532
rect 265158 163520 265164 163532
rect 242216 163492 265164 163520
rect 242216 163480 242222 163492
rect 265158 163480 265164 163492
rect 265216 163480 265222 163532
rect 234062 163004 234068 163056
rect 234120 163044 234126 163056
rect 265802 163044 265808 163056
rect 234120 163016 265808 163044
rect 234120 163004 234126 163016
rect 265802 163004 265808 163016
rect 265860 163004 265866 163056
rect 258718 162868 258724 162920
rect 258776 162908 258782 162920
rect 265526 162908 265532 162920
rect 258776 162880 265532 162908
rect 258776 162868 258782 162880
rect 265526 162868 265532 162880
rect 265584 162868 265590 162920
rect 282730 162868 282736 162920
rect 282788 162908 282794 162920
rect 288618 162908 288624 162920
rect 282788 162880 288624 162908
rect 282788 162868 282794 162880
rect 288618 162868 288624 162880
rect 288676 162868 288682 162920
rect 170582 162800 170588 162852
rect 170640 162840 170646 162852
rect 213914 162840 213920 162852
rect 170640 162812 213920 162840
rect 170640 162800 170646 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 231026 162800 231032 162852
rect 231084 162840 231090 162852
rect 233326 162840 233332 162852
rect 231084 162812 233332 162840
rect 231084 162800 231090 162812
rect 233326 162800 233332 162812
rect 233384 162800 233390 162852
rect 282546 162800 282552 162852
rect 282604 162840 282610 162852
rect 294230 162840 294236 162852
rect 282604 162812 294236 162840
rect 282604 162800 282610 162812
rect 294230 162800 294236 162812
rect 294288 162800 294294 162852
rect 282822 162732 282828 162784
rect 282880 162772 282886 162784
rect 292850 162772 292856 162784
rect 282880 162744 292856 162772
rect 282880 162732 282886 162744
rect 292850 162732 292856 162744
rect 292908 162732 292914 162784
rect 231670 162664 231676 162716
rect 231728 162704 231734 162716
rect 244366 162704 244372 162716
rect 231728 162676 244372 162704
rect 231728 162664 231734 162676
rect 244366 162664 244372 162676
rect 244424 162664 244430 162716
rect 231762 162460 231768 162512
rect 231820 162500 231826 162512
rect 236638 162500 236644 162512
rect 231820 162472 236644 162500
rect 231820 162460 231826 162472
rect 236638 162460 236644 162472
rect 236696 162460 236702 162512
rect 233878 162120 233884 162172
rect 233936 162160 233942 162172
rect 247126 162160 247132 162172
rect 233936 162132 247132 162160
rect 233936 162120 233942 162132
rect 247126 162120 247132 162132
rect 247184 162120 247190 162172
rect 253382 161576 253388 161628
rect 253440 161616 253446 161628
rect 264422 161616 264428 161628
rect 253440 161588 264428 161616
rect 253440 161576 253446 161588
rect 264422 161576 264428 161588
rect 264480 161576 264486 161628
rect 247678 161508 247684 161560
rect 247736 161548 247742 161560
rect 265526 161548 265532 161560
rect 247736 161520 265532 161548
rect 247736 161508 247742 161520
rect 265526 161508 265532 161520
rect 265584 161508 265590 161560
rect 241054 161440 241060 161492
rect 241112 161480 241118 161492
rect 264514 161480 264520 161492
rect 241112 161452 264520 161480
rect 241112 161440 241118 161452
rect 264514 161440 264520 161452
rect 264572 161440 264578 161492
rect 188430 161372 188436 161424
rect 188488 161412 188494 161424
rect 213914 161412 213920 161424
rect 188488 161384 213920 161412
rect 188488 161372 188494 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 231670 161372 231676 161424
rect 231728 161412 231734 161424
rect 248598 161412 248604 161424
rect 231728 161384 248604 161412
rect 231728 161372 231734 161384
rect 248598 161372 248604 161384
rect 248656 161372 248662 161424
rect 282822 161372 282828 161424
rect 282880 161412 282886 161424
rect 302326 161412 302332 161424
rect 282880 161384 302332 161412
rect 282880 161372 282886 161384
rect 302326 161372 302332 161384
rect 302384 161372 302390 161424
rect 231762 161304 231768 161356
rect 231820 161344 231826 161356
rect 238754 161344 238760 161356
rect 231820 161316 238760 161344
rect 231820 161304 231826 161316
rect 238754 161304 238760 161316
rect 238812 161304 238818 161356
rect 282362 161304 282368 161356
rect 282420 161344 282426 161356
rect 292758 161344 292764 161356
rect 282420 161316 292764 161344
rect 282420 161304 282426 161316
rect 292758 161304 292764 161316
rect 292816 161304 292822 161356
rect 167730 160692 167736 160744
rect 167788 160732 167794 160744
rect 214098 160732 214104 160744
rect 167788 160704 214104 160732
rect 167788 160692 167794 160704
rect 214098 160692 214104 160704
rect 214156 160692 214162 160744
rect 247862 160216 247868 160268
rect 247920 160256 247926 160268
rect 265894 160256 265900 160268
rect 247920 160228 265900 160256
rect 247920 160216 247926 160228
rect 265894 160216 265900 160228
rect 265952 160216 265958 160268
rect 245010 160148 245016 160200
rect 245068 160188 245074 160200
rect 265802 160188 265808 160200
rect 245068 160160 265808 160188
rect 245068 160148 245074 160160
rect 265802 160148 265808 160160
rect 265860 160148 265866 160200
rect 242342 160080 242348 160132
rect 242400 160120 242406 160132
rect 265986 160120 265992 160132
rect 242400 160092 265992 160120
rect 242400 160080 242406 160092
rect 265986 160080 265992 160092
rect 266044 160080 266050 160132
rect 169018 160012 169024 160064
rect 169076 160052 169082 160064
rect 213914 160052 213920 160064
rect 169076 160024 213920 160052
rect 169076 160012 169082 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231762 160012 231768 160064
rect 231820 160052 231826 160064
rect 247218 160052 247224 160064
rect 231820 160024 247224 160052
rect 231820 160012 231826 160024
rect 247218 160012 247224 160024
rect 247276 160012 247282 160064
rect 184290 159944 184296 159996
rect 184348 159984 184354 159996
rect 214006 159984 214012 159996
rect 184348 159956 214012 159984
rect 184348 159944 184354 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 231670 159944 231676 159996
rect 231728 159984 231734 159996
rect 240318 159984 240324 159996
rect 231728 159956 240324 159984
rect 231728 159944 231734 159956
rect 240318 159944 240324 159956
rect 240376 159944 240382 159996
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 234706 159508 234712 159520
rect 231728 159480 234712 159508
rect 231728 159468 231734 159480
rect 234706 159468 234712 159480
rect 234764 159468 234770 159520
rect 261754 158788 261760 158840
rect 261812 158828 261818 158840
rect 265434 158828 265440 158840
rect 261812 158800 265440 158828
rect 261812 158788 261818 158800
rect 265434 158788 265440 158800
rect 265492 158788 265498 158840
rect 246574 158720 246580 158772
rect 246632 158760 246638 158772
rect 265526 158760 265532 158772
rect 246632 158732 265532 158760
rect 246632 158720 246638 158732
rect 265526 158720 265532 158732
rect 265584 158720 265590 158772
rect 282270 158652 282276 158704
rect 282328 158692 282334 158704
rect 299750 158692 299756 158704
rect 282328 158664 299756 158692
rect 282328 158652 282334 158664
rect 299750 158652 299756 158664
rect 299808 158652 299814 158704
rect 170674 157972 170680 158024
rect 170732 158012 170738 158024
rect 214926 158012 214932 158024
rect 170732 157984 214932 158012
rect 170732 157972 170738 157984
rect 214926 157972 214932 157984
rect 214984 157972 214990 158024
rect 256142 157972 256148 158024
rect 256200 158012 256206 158024
rect 265802 158012 265808 158024
rect 256200 157984 265808 158012
rect 256200 157972 256206 157984
rect 265802 157972 265808 157984
rect 265860 157972 265866 158024
rect 245102 157428 245108 157480
rect 245160 157468 245166 157480
rect 265802 157468 265808 157480
rect 245160 157440 265808 157468
rect 245160 157428 245166 157440
rect 265802 157428 265808 157440
rect 265860 157428 265866 157480
rect 237374 157360 237380 157412
rect 237432 157400 237438 157412
rect 265986 157400 265992 157412
rect 237432 157372 265992 157400
rect 237432 157360 237438 157372
rect 265986 157360 265992 157372
rect 266044 157360 266050 157412
rect 167638 157292 167644 157344
rect 167696 157332 167702 157344
rect 214006 157332 214012 157344
rect 167696 157304 214012 157332
rect 167696 157292 167702 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 231670 157292 231676 157344
rect 231728 157332 231734 157344
rect 258074 157332 258080 157344
rect 231728 157304 258080 157332
rect 231728 157292 231734 157304
rect 258074 157292 258080 157304
rect 258132 157292 258138 157344
rect 282822 157292 282828 157344
rect 282880 157332 282886 157344
rect 301038 157332 301044 157344
rect 282880 157304 301044 157332
rect 282880 157292 282886 157304
rect 301038 157292 301044 157304
rect 301096 157292 301102 157344
rect 171870 157224 171876 157276
rect 171928 157264 171934 157276
rect 213914 157264 213920 157276
rect 171928 157236 213920 157264
rect 171928 157224 171934 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 231762 157224 231768 157276
rect 231820 157264 231826 157276
rect 244458 157264 244464 157276
rect 231820 157236 244464 157264
rect 231820 157224 231826 157236
rect 244458 157224 244464 157236
rect 244516 157224 244522 157276
rect 239582 156612 239588 156664
rect 239640 156652 239646 156664
rect 265066 156652 265072 156664
rect 239640 156624 265072 156652
rect 239640 156612 239646 156624
rect 265066 156612 265072 156624
rect 265124 156612 265130 156664
rect 232774 156136 232780 156188
rect 232832 156176 232838 156188
rect 237466 156176 237472 156188
rect 232832 156148 237472 156176
rect 232832 156136 232838 156148
rect 237466 156136 237472 156148
rect 237524 156136 237530 156188
rect 250438 156000 250444 156052
rect 250496 156040 250502 156052
rect 265894 156040 265900 156052
rect 250496 156012 265900 156040
rect 250496 156000 250502 156012
rect 265894 156000 265900 156012
rect 265952 156000 265958 156052
rect 238018 155932 238024 155984
rect 238076 155972 238082 155984
rect 265802 155972 265808 155984
rect 238076 155944 265808 155972
rect 238076 155932 238082 155944
rect 265802 155932 265808 155944
rect 265860 155932 265866 155984
rect 169110 155864 169116 155916
rect 169168 155904 169174 155916
rect 213914 155904 213920 155916
rect 169168 155876 213920 155904
rect 169168 155864 169174 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 230934 155864 230940 155916
rect 230992 155904 230998 155916
rect 233510 155904 233516 155916
rect 230992 155876 233516 155904
rect 230992 155864 230998 155876
rect 233510 155864 233516 155876
rect 233568 155864 233574 155916
rect 282822 155864 282828 155916
rect 282880 155904 282886 155916
rect 302510 155904 302516 155916
rect 282880 155876 302516 155904
rect 282880 155864 282886 155876
rect 302510 155864 302516 155876
rect 302568 155864 302574 155916
rect 230566 155796 230572 155848
rect 230624 155836 230630 155848
rect 232130 155836 232136 155848
rect 230624 155808 232136 155836
rect 230624 155796 230630 155808
rect 232130 155796 232136 155808
rect 232188 155796 232194 155848
rect 263134 154708 263140 154760
rect 263192 154748 263198 154760
rect 265802 154748 265808 154760
rect 263192 154720 265808 154748
rect 263192 154708 263198 154720
rect 265802 154708 265808 154720
rect 265860 154708 265866 154760
rect 240962 154640 240968 154692
rect 241020 154680 241026 154692
rect 265986 154680 265992 154692
rect 241020 154652 265992 154680
rect 241020 154640 241026 154652
rect 265986 154640 265992 154652
rect 266044 154640 266050 154692
rect 233970 154572 233976 154624
rect 234028 154612 234034 154624
rect 265710 154612 265716 154624
rect 234028 154584 265716 154612
rect 234028 154572 234034 154584
rect 265710 154572 265716 154584
rect 265768 154572 265774 154624
rect 231394 154504 231400 154556
rect 231452 154544 231458 154556
rect 252554 154544 252560 154556
rect 231452 154516 252560 154544
rect 231452 154504 231458 154516
rect 252554 154504 252560 154516
rect 252612 154504 252618 154556
rect 231762 154300 231768 154352
rect 231820 154340 231826 154352
rect 236178 154340 236184 154352
rect 231820 154312 236184 154340
rect 231820 154300 231826 154312
rect 236178 154300 236184 154312
rect 236236 154300 236242 154352
rect 281902 154164 281908 154216
rect 281960 154204 281966 154216
rect 285950 154204 285956 154216
rect 281960 154176 285956 154204
rect 281960 154164 281966 154176
rect 285950 154164 285956 154176
rect 286008 154164 286014 154216
rect 231118 154096 231124 154148
rect 231176 154136 231182 154148
rect 237374 154136 237380 154148
rect 231176 154108 237380 154136
rect 231176 154096 231182 154108
rect 237374 154096 237380 154108
rect 237432 154096 237438 154148
rect 239398 153824 239404 153876
rect 239456 153864 239462 153876
rect 265894 153864 265900 153876
rect 239456 153836 265900 153864
rect 239456 153824 239462 153836
rect 265894 153824 265900 153836
rect 265952 153824 265958 153876
rect 231302 153348 231308 153400
rect 231360 153388 231366 153400
rect 233878 153388 233884 153400
rect 231360 153360 233884 153388
rect 231360 153348 231366 153360
rect 233878 153348 233884 153360
rect 233936 153348 233942 153400
rect 196802 153280 196808 153332
rect 196860 153320 196866 153332
rect 213914 153320 213920 153332
rect 196860 153292 213920 153320
rect 196860 153280 196866 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 258810 153280 258816 153332
rect 258868 153320 258874 153332
rect 265802 153320 265808 153332
rect 258868 153292 265808 153320
rect 258868 153280 258874 153292
rect 265802 153280 265808 153292
rect 265860 153280 265866 153332
rect 281718 153280 281724 153332
rect 281776 153320 281782 153332
rect 284478 153320 284484 153332
rect 281776 153292 284484 153320
rect 281776 153280 281782 153292
rect 284478 153280 284484 153292
rect 284536 153280 284542 153332
rect 167638 153212 167644 153264
rect 167696 153252 167702 153264
rect 214006 153252 214012 153264
rect 167696 153224 214012 153252
rect 167696 153212 167702 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 238202 153212 238208 153264
rect 238260 153252 238266 153264
rect 265342 153252 265348 153264
rect 238260 153224 265348 153252
rect 238260 153212 238266 153224
rect 265342 153212 265348 153224
rect 265400 153212 265406 153264
rect 230750 153144 230756 153196
rect 230808 153184 230814 153196
rect 255314 153184 255320 153196
rect 230808 153156 255320 153184
rect 230808 153144 230814 153156
rect 255314 153144 255320 153156
rect 255372 153144 255378 153196
rect 282178 153144 282184 153196
rect 282236 153184 282242 153196
rect 308030 153184 308036 153196
rect 282236 153156 308036 153184
rect 282236 153144 282242 153156
rect 308030 153144 308036 153156
rect 308088 153144 308094 153196
rect 468478 153144 468484 153196
rect 468536 153184 468542 153196
rect 579798 153184 579804 153196
rect 468536 153156 579804 153184
rect 468536 153144 468542 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 231762 153076 231768 153128
rect 231820 153116 231826 153128
rect 245746 153116 245752 153128
rect 231820 153088 245752 153116
rect 231820 153076 231826 153088
rect 245746 153076 245752 153088
rect 245804 153076 245810 153128
rect 231670 152668 231676 152720
rect 231728 152708 231734 152720
rect 234614 152708 234620 152720
rect 231728 152680 234620 152708
rect 231728 152668 231734 152680
rect 234614 152668 234620 152680
rect 234672 152668 234678 152720
rect 211798 152396 211804 152448
rect 211856 152436 211862 152448
rect 213914 152436 213920 152448
rect 211856 152408 213920 152436
rect 211856 152396 211862 152408
rect 213914 152396 213920 152408
rect 213972 152396 213978 152448
rect 235442 151920 235448 151972
rect 235500 151960 235506 151972
rect 265250 151960 265256 151972
rect 235500 151932 265256 151960
rect 235500 151920 235506 151932
rect 265250 151920 265256 151932
rect 265308 151920 265314 151972
rect 253198 151852 253204 151904
rect 253256 151892 253262 151904
rect 265802 151892 265808 151904
rect 253256 151864 265808 151892
rect 253256 151852 253262 151864
rect 265802 151852 265808 151864
rect 265860 151852 265866 151904
rect 171778 151784 171784 151836
rect 171836 151824 171842 151836
rect 213914 151824 213920 151836
rect 171836 151796 213920 151824
rect 171836 151784 171842 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 231670 151716 231676 151768
rect 231728 151756 231734 151768
rect 252646 151756 252652 151768
rect 231728 151728 252652 151756
rect 231728 151716 231734 151728
rect 252646 151716 252652 151728
rect 252704 151716 252710 151768
rect 282822 151716 282828 151768
rect 282880 151756 282886 151768
rect 299658 151756 299664 151768
rect 282880 151728 299664 151756
rect 282880 151716 282886 151728
rect 299658 151716 299664 151728
rect 299716 151716 299722 151768
rect 231762 151648 231768 151700
rect 231820 151688 231826 151700
rect 251358 151688 251364 151700
rect 231820 151660 251364 151688
rect 231820 151648 231826 151660
rect 251358 151648 251364 151660
rect 251416 151648 251422 151700
rect 281994 151648 282000 151700
rect 282052 151688 282058 151700
rect 289998 151688 290004 151700
rect 282052 151660 290004 151688
rect 282052 151648 282058 151660
rect 289998 151648 290004 151660
rect 290056 151648 290062 151700
rect 260466 150560 260472 150612
rect 260524 150600 260530 150612
rect 265710 150600 265716 150612
rect 260524 150572 265716 150600
rect 260524 150560 260530 150572
rect 265710 150560 265716 150572
rect 265768 150560 265774 150612
rect 245194 150492 245200 150544
rect 245252 150532 245258 150544
rect 265802 150532 265808 150544
rect 245252 150504 265808 150532
rect 245252 150492 245258 150504
rect 265802 150492 265808 150504
rect 265860 150492 265866 150544
rect 173342 150424 173348 150476
rect 173400 150464 173406 150476
rect 213914 150464 213920 150476
rect 173400 150436 213920 150464
rect 173400 150424 173406 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 236822 150424 236828 150476
rect 236880 150464 236886 150476
rect 265434 150464 265440 150476
rect 236880 150436 265440 150464
rect 236880 150424 236886 150436
rect 265434 150424 265440 150436
rect 265492 150424 265498 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 32398 150396 32404 150408
rect 3476 150368 32404 150396
rect 3476 150356 3482 150368
rect 32398 150356 32404 150368
rect 32456 150356 32462 150408
rect 210510 150356 210516 150408
rect 210568 150396 210574 150408
rect 214006 150396 214012 150408
rect 210568 150368 214012 150396
rect 210568 150356 210574 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 230934 150356 230940 150408
rect 230992 150396 230998 150408
rect 256786 150396 256792 150408
rect 230992 150368 256792 150396
rect 230992 150356 230998 150368
rect 256786 150356 256792 150368
rect 256844 150356 256850 150408
rect 282822 150356 282828 150408
rect 282880 150396 282886 150408
rect 296898 150396 296904 150408
rect 282880 150368 296904 150396
rect 282880 150356 282886 150368
rect 296898 150356 296904 150368
rect 296956 150356 296962 150408
rect 231026 150288 231032 150340
rect 231084 150328 231090 150340
rect 234890 150328 234896 150340
rect 231084 150300 234896 150328
rect 231084 150288 231090 150300
rect 234890 150288 234896 150300
rect 234948 150288 234954 150340
rect 282178 150288 282184 150340
rect 282236 150328 282242 150340
rect 291378 150328 291384 150340
rect 282236 150300 291384 150328
rect 282236 150288 282242 150300
rect 291378 150288 291384 150300
rect 291436 150288 291442 150340
rect 231210 149744 231216 149796
rect 231268 149784 231274 149796
rect 250438 149784 250444 149796
rect 231268 149756 250444 149784
rect 231268 149744 231274 149756
rect 250438 149744 250444 149756
rect 250496 149744 250502 149796
rect 236914 149676 236920 149728
rect 236972 149716 236978 149728
rect 265894 149716 265900 149728
rect 236972 149688 265900 149716
rect 236972 149676 236978 149688
rect 265894 149676 265900 149688
rect 265952 149676 265958 149728
rect 231302 149472 231308 149524
rect 231360 149512 231366 149524
rect 235994 149512 236000 149524
rect 231360 149484 236000 149512
rect 231360 149472 231366 149484
rect 235994 149472 236000 149484
rect 236052 149472 236058 149524
rect 259086 149132 259092 149184
rect 259144 149172 259150 149184
rect 265342 149172 265348 149184
rect 259144 149144 265348 149172
rect 259144 149132 259150 149144
rect 265342 149132 265348 149144
rect 265400 149132 265406 149184
rect 250714 149064 250720 149116
rect 250772 149104 250778 149116
rect 265802 149104 265808 149116
rect 250772 149076 265808 149104
rect 250772 149064 250778 149076
rect 265802 149064 265808 149076
rect 265860 149064 265866 149116
rect 166258 148996 166264 149048
rect 166316 149036 166322 149048
rect 213914 149036 213920 149048
rect 166316 149008 213920 149036
rect 166316 148996 166322 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 251450 149036 251456 149048
rect 231820 149008 251456 149036
rect 231820 148996 231826 149008
rect 251450 148996 251456 149008
rect 251508 148996 251514 149048
rect 282086 148928 282092 148980
rect 282144 148968 282150 148980
rect 309318 148968 309324 148980
rect 282144 148940 309324 148968
rect 282144 148928 282150 148940
rect 309318 148928 309324 148940
rect 309376 148928 309382 148980
rect 257522 148316 257528 148368
rect 257580 148356 257586 148368
rect 265434 148356 265440 148368
rect 257580 148328 265440 148356
rect 257580 148316 257586 148328
rect 265434 148316 265440 148328
rect 265492 148316 265498 148368
rect 235534 147704 235540 147756
rect 235592 147744 235598 147756
rect 265710 147744 265716 147756
rect 235592 147716 265716 147744
rect 235592 147704 235598 147716
rect 265710 147704 265716 147716
rect 265768 147704 265774 147756
rect 187142 147636 187148 147688
rect 187200 147676 187206 147688
rect 213914 147676 213920 147688
rect 187200 147648 213920 147676
rect 187200 147636 187206 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 233878 147636 233884 147688
rect 233936 147676 233942 147688
rect 265526 147676 265532 147688
rect 233936 147648 265532 147676
rect 233936 147636 233942 147648
rect 265526 147636 265532 147648
rect 265584 147636 265590 147688
rect 230934 147568 230940 147620
rect 230992 147608 230998 147620
rect 234798 147608 234804 147620
rect 230992 147580 234804 147608
rect 230992 147568 230998 147580
rect 234798 147568 234804 147580
rect 234856 147568 234862 147620
rect 281718 147568 281724 147620
rect 281776 147608 281782 147620
rect 305178 147608 305184 147620
rect 281776 147580 305184 147608
rect 281776 147568 281782 147580
rect 305178 147568 305184 147580
rect 305236 147568 305242 147620
rect 230750 147500 230756 147552
rect 230808 147540 230814 147552
rect 232498 147540 232504 147552
rect 230808 147512 232504 147540
rect 230808 147500 230814 147512
rect 232498 147500 232504 147512
rect 232556 147500 232562 147552
rect 231394 146956 231400 147008
rect 231452 146996 231458 147008
rect 242526 146996 242532 147008
rect 231452 146968 242532 146996
rect 231452 146956 231458 146968
rect 242526 146956 242532 146968
rect 242584 146956 242590 147008
rect 242250 146888 242256 146940
rect 242308 146928 242314 146940
rect 265066 146928 265072 146940
rect 242308 146900 265072 146928
rect 242308 146888 242314 146900
rect 265066 146888 265072 146900
rect 265124 146888 265130 146940
rect 261570 146344 261576 146396
rect 261628 146384 261634 146396
rect 265894 146384 265900 146396
rect 261628 146356 265900 146384
rect 261628 146344 261634 146356
rect 265894 146344 265900 146356
rect 265952 146344 265958 146396
rect 171870 146276 171876 146328
rect 171928 146316 171934 146328
rect 213914 146316 213920 146328
rect 171928 146288 213920 146316
rect 171928 146276 171934 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 235626 146276 235632 146328
rect 235684 146316 235690 146328
rect 265526 146316 265532 146328
rect 235684 146288 265532 146316
rect 235684 146276 235690 146288
rect 265526 146276 265532 146288
rect 265584 146276 265590 146328
rect 231762 146208 231768 146260
rect 231820 146248 231826 146260
rect 249794 146248 249800 146260
rect 231820 146220 249800 146248
rect 231820 146208 231826 146220
rect 249794 146208 249800 146220
rect 249852 146208 249858 146260
rect 282822 146208 282828 146260
rect 282880 146248 282886 146260
rect 307938 146248 307944 146260
rect 282880 146220 307944 146248
rect 282880 146208 282886 146220
rect 307938 146208 307944 146220
rect 307996 146208 308002 146260
rect 231670 146140 231676 146192
rect 231728 146180 231734 146192
rect 247034 146180 247040 146192
rect 231728 146152 247040 146180
rect 231728 146140 231734 146152
rect 247034 146140 247040 146152
rect 247092 146140 247098 146192
rect 282730 146140 282736 146192
rect 282788 146180 282794 146192
rect 296990 146180 296996 146192
rect 282788 146152 296996 146180
rect 282788 146140 282794 146152
rect 296990 146140 296996 146152
rect 297048 146140 297054 146192
rect 254762 145052 254768 145104
rect 254820 145092 254826 145104
rect 265894 145092 265900 145104
rect 254820 145064 265900 145092
rect 254820 145052 254826 145064
rect 265894 145052 265900 145064
rect 265952 145052 265958 145104
rect 243814 144984 243820 145036
rect 243872 145024 243878 145036
rect 265710 145024 265716 145036
rect 243872 144996 265716 145024
rect 243872 144984 243878 144996
rect 265710 144984 265716 144996
rect 265768 144984 265774 145036
rect 189810 144916 189816 144968
rect 189868 144956 189874 144968
rect 213914 144956 213920 144968
rect 189868 144928 213920 144956
rect 189868 144916 189874 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 234154 144916 234160 144968
rect 234212 144956 234218 144968
rect 265802 144956 265808 144968
rect 234212 144928 265808 144956
rect 234212 144916 234218 144928
rect 265802 144916 265808 144928
rect 265860 144916 265866 144968
rect 231762 144848 231768 144900
rect 231820 144888 231826 144900
rect 248414 144888 248420 144900
rect 231820 144860 248420 144888
rect 231820 144848 231826 144860
rect 248414 144848 248420 144860
rect 248472 144848 248478 144900
rect 282822 144848 282828 144900
rect 282880 144888 282886 144900
rect 298186 144888 298192 144900
rect 282880 144860 298192 144888
rect 282880 144848 282886 144860
rect 298186 144848 298192 144860
rect 298244 144848 298250 144900
rect 174630 144168 174636 144220
rect 174688 144208 174694 144220
rect 214650 144208 214656 144220
rect 174688 144180 214656 144208
rect 174688 144168 174694 144180
rect 214650 144168 214656 144180
rect 214708 144168 214714 144220
rect 230750 144168 230756 144220
rect 230808 144208 230814 144220
rect 232682 144208 232688 144220
rect 230808 144180 232688 144208
rect 230808 144168 230814 144180
rect 232682 144168 232688 144180
rect 232740 144168 232746 144220
rect 265986 144208 265992 144220
rect 238726 144180 265992 144208
rect 232590 144100 232596 144152
rect 232648 144140 232654 144152
rect 238726 144140 238754 144180
rect 265986 144168 265992 144180
rect 266044 144168 266050 144220
rect 232648 144112 238754 144140
rect 232648 144100 232654 144112
rect 282822 143692 282828 143744
rect 282880 143732 282886 143744
rect 287146 143732 287152 143744
rect 282880 143704 287152 143732
rect 282880 143692 282886 143704
rect 287146 143692 287152 143704
rect 287204 143692 287210 143744
rect 182818 143556 182824 143608
rect 182876 143596 182882 143608
rect 213914 143596 213920 143608
rect 182876 143568 213920 143596
rect 182876 143556 182882 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 262950 143556 262956 143608
rect 263008 143596 263014 143608
rect 265526 143596 265532 143608
rect 263008 143568 265532 143596
rect 263008 143556 263014 143568
rect 265526 143556 265532 143568
rect 265584 143556 265590 143608
rect 231762 143488 231768 143540
rect 231820 143528 231826 143540
rect 242894 143528 242900 143540
rect 231820 143500 242900 143528
rect 231820 143488 231826 143500
rect 242894 143488 242900 143500
rect 242952 143488 242958 143540
rect 282086 143488 282092 143540
rect 282144 143528 282150 143540
rect 306558 143528 306564 143540
rect 282144 143500 306564 143528
rect 282144 143488 282150 143500
rect 306558 143488 306564 143500
rect 306616 143488 306622 143540
rect 230474 143420 230480 143472
rect 230532 143460 230538 143472
rect 232774 143460 232780 143472
rect 230532 143432 232780 143460
rect 230532 143420 230538 143432
rect 232774 143420 232780 143432
rect 232832 143420 232838 143472
rect 282270 143420 282276 143472
rect 282328 143460 282334 143472
rect 298278 143460 298284 143472
rect 282328 143432 298284 143460
rect 282328 143420 282334 143432
rect 298278 143420 298284 143432
rect 298336 143420 298342 143472
rect 282178 142944 282184 142996
rect 282236 142984 282242 142996
rect 285674 142984 285680 142996
rect 282236 142956 285680 142984
rect 282236 142944 282242 142956
rect 285674 142944 285680 142956
rect 285732 142944 285738 142996
rect 167730 142808 167736 142860
rect 167788 142848 167794 142860
rect 214006 142848 214012 142860
rect 167788 142820 214012 142848
rect 167788 142808 167794 142820
rect 214006 142808 214012 142820
rect 214064 142808 214070 142860
rect 232682 142808 232688 142860
rect 232740 142848 232746 142860
rect 265802 142848 265808 142860
rect 232740 142820 265808 142848
rect 232740 142808 232746 142820
rect 265802 142808 265808 142820
rect 265860 142808 265866 142860
rect 195422 142196 195428 142248
rect 195480 142236 195486 142248
rect 213914 142236 213920 142248
rect 195480 142208 213920 142236
rect 195480 142196 195486 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 184290 142128 184296 142180
rect 184348 142168 184354 142180
rect 214006 142168 214012 142180
rect 184348 142140 214012 142168
rect 184348 142128 184354 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 252094 142128 252100 142180
rect 252152 142168 252158 142180
rect 265342 142168 265348 142180
rect 252152 142140 265348 142168
rect 252152 142128 252158 142140
rect 265342 142128 265348 142140
rect 265400 142128 265406 142180
rect 282822 142060 282828 142112
rect 282880 142100 282886 142112
rect 310698 142100 310704 142112
rect 282880 142072 310704 142100
rect 282880 142060 282886 142072
rect 310698 142060 310704 142072
rect 310756 142060 310762 142112
rect 282730 141992 282736 142044
rect 282788 142032 282794 142044
rect 295518 142032 295524 142044
rect 282788 142004 295524 142032
rect 282788 141992 282794 142004
rect 295518 141992 295524 142004
rect 295576 141992 295582 142044
rect 176010 140836 176016 140888
rect 176068 140876 176074 140888
rect 213914 140876 213920 140888
rect 176068 140848 213920 140876
rect 176068 140836 176074 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 250806 140836 250812 140888
rect 250864 140876 250870 140888
rect 265526 140876 265532 140888
rect 250864 140848 265532 140876
rect 250864 140836 250870 140848
rect 265526 140836 265532 140848
rect 265584 140836 265590 140888
rect 169018 140768 169024 140820
rect 169076 140808 169082 140820
rect 214006 140808 214012 140820
rect 169076 140780 214012 140808
rect 169076 140768 169082 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 232774 140768 232780 140820
rect 232832 140808 232838 140820
rect 264422 140808 264428 140820
rect 232832 140780 264428 140808
rect 232832 140768 232838 140780
rect 264422 140768 264428 140780
rect 264480 140768 264486 140820
rect 231486 140700 231492 140752
rect 231544 140740 231550 140752
rect 262214 140740 262220 140752
rect 231544 140712 262220 140740
rect 231544 140700 231550 140712
rect 262214 140700 262220 140712
rect 262272 140700 262278 140752
rect 282822 140700 282828 140752
rect 282880 140740 282886 140752
rect 287330 140740 287336 140752
rect 282880 140712 287336 140740
rect 282880 140700 282886 140712
rect 287330 140700 287336 140712
rect 287388 140700 287394 140752
rect 231762 140632 231768 140684
rect 231820 140672 231826 140684
rect 260834 140672 260840 140684
rect 231820 140644 260840 140672
rect 231820 140632 231826 140644
rect 260834 140632 260840 140644
rect 260892 140632 260898 140684
rect 230934 140564 230940 140616
rect 230992 140604 230998 140616
rect 248506 140604 248512 140616
rect 230992 140576 248512 140604
rect 230992 140564 230998 140576
rect 248506 140564 248512 140576
rect 248564 140564 248570 140616
rect 169110 140020 169116 140072
rect 169168 140060 169174 140072
rect 214466 140060 214472 140072
rect 169168 140032 214472 140060
rect 169168 140020 169174 140032
rect 214466 140020 214472 140032
rect 214524 140020 214530 140072
rect 253566 140020 253572 140072
rect 253624 140060 253630 140072
rect 265802 140060 265808 140072
rect 253624 140032 265808 140060
rect 253624 140020 253630 140032
rect 265802 140020 265808 140032
rect 265860 140020 265866 140072
rect 236730 139476 236736 139528
rect 236788 139516 236794 139528
rect 265802 139516 265808 139528
rect 236788 139488 265808 139516
rect 236788 139476 236794 139488
rect 265802 139476 265808 139488
rect 265860 139476 265866 139528
rect 170582 139408 170588 139460
rect 170640 139448 170646 139460
rect 213914 139448 213920 139460
rect 170640 139420 213920 139448
rect 170640 139408 170646 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 230014 139408 230020 139460
rect 230072 139448 230078 139460
rect 265710 139448 265716 139460
rect 230072 139420 265716 139448
rect 230072 139408 230078 139420
rect 265710 139408 265716 139420
rect 265768 139408 265774 139460
rect 231762 139340 231768 139392
rect 231820 139380 231826 139392
rect 251266 139380 251272 139392
rect 231820 139352 251272 139380
rect 231820 139340 231826 139352
rect 251266 139340 251272 139352
rect 251324 139340 251330 139392
rect 282822 139340 282828 139392
rect 282880 139380 282886 139392
rect 307846 139380 307852 139392
rect 282880 139352 307852 139380
rect 282880 139340 282886 139352
rect 307846 139340 307852 139352
rect 307904 139340 307910 139392
rect 282730 139272 282736 139324
rect 282788 139312 282794 139324
rect 305270 139312 305276 139324
rect 282788 139284 305276 139312
rect 282788 139272 282794 139284
rect 305270 139272 305276 139284
rect 305328 139272 305334 139324
rect 231670 139204 231676 139256
rect 231728 139244 231734 139256
rect 236086 139244 236092 139256
rect 231728 139216 236092 139244
rect 231728 139204 231734 139216
rect 236086 139204 236092 139216
rect 236144 139204 236150 139256
rect 181438 138660 181444 138712
rect 181496 138700 181502 138712
rect 214006 138700 214012 138712
rect 181496 138672 214012 138700
rect 181496 138660 181502 138672
rect 214006 138660 214012 138672
rect 214064 138660 214070 138712
rect 231026 138660 231032 138712
rect 231084 138700 231090 138712
rect 241146 138700 241152 138712
rect 231084 138672 241152 138700
rect 231084 138660 231090 138672
rect 241146 138660 241152 138672
rect 241204 138660 241210 138712
rect 251910 138048 251916 138100
rect 251968 138088 251974 138100
rect 265158 138088 265164 138100
rect 251968 138060 265164 138088
rect 251968 138048 251974 138060
rect 265158 138048 265164 138060
rect 265216 138048 265222 138100
rect 170490 137980 170496 138032
rect 170548 138020 170554 138032
rect 213914 138020 213920 138032
rect 170548 137992 213920 138020
rect 170548 137980 170554 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 240870 137980 240876 138032
rect 240928 138020 240934 138032
rect 265802 138020 265808 138032
rect 240928 137992 265808 138020
rect 240928 137980 240934 137992
rect 265802 137980 265808 137992
rect 265860 137980 265866 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 15838 137952 15844 137964
rect 3292 137924 15844 137952
rect 3292 137912 3298 137924
rect 15838 137912 15844 137924
rect 15896 137912 15902 137964
rect 231486 137912 231492 137964
rect 231544 137952 231550 137964
rect 259454 137952 259460 137964
rect 231544 137924 259460 137952
rect 231544 137912 231550 137924
rect 259454 137912 259460 137924
rect 259512 137912 259518 137964
rect 282822 137912 282828 137964
rect 282880 137952 282886 137964
rect 295610 137952 295616 137964
rect 282880 137924 295616 137952
rect 282880 137912 282886 137924
rect 295610 137912 295616 137924
rect 295668 137912 295674 137964
rect 231762 137844 231768 137896
rect 231820 137884 231826 137896
rect 256694 137884 256700 137896
rect 231820 137856 256700 137884
rect 231820 137844 231826 137856
rect 256694 137844 256700 137856
rect 256752 137844 256758 137896
rect 249334 137232 249340 137284
rect 249392 137272 249398 137284
rect 265250 137272 265256 137284
rect 249392 137244 265256 137272
rect 249392 137232 249398 137244
rect 265250 137232 265256 137244
rect 265308 137232 265314 137284
rect 236638 136688 236644 136740
rect 236696 136728 236702 136740
rect 265710 136728 265716 136740
rect 236696 136700 265716 136728
rect 236696 136688 236702 136700
rect 265710 136688 265716 136700
rect 265768 136688 265774 136740
rect 192570 136620 192576 136672
rect 192628 136660 192634 136672
rect 213914 136660 213920 136672
rect 192628 136632 213920 136660
rect 192628 136620 192634 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 229922 136620 229928 136672
rect 229980 136660 229986 136672
rect 265802 136660 265808 136672
rect 229980 136632 265808 136660
rect 229980 136620 229986 136632
rect 265802 136620 265808 136632
rect 265860 136620 265866 136672
rect 231762 136552 231768 136604
rect 231820 136592 231826 136604
rect 254026 136592 254032 136604
rect 231820 136564 254032 136592
rect 231820 136552 231826 136564
rect 254026 136552 254032 136564
rect 254084 136552 254090 136604
rect 282730 136552 282736 136604
rect 282788 136592 282794 136604
rect 309226 136592 309232 136604
rect 282788 136564 309232 136592
rect 282788 136552 282794 136564
rect 309226 136552 309232 136564
rect 309284 136552 309290 136604
rect 231670 136484 231676 136536
rect 231728 136524 231734 136536
rect 243722 136524 243728 136536
rect 231728 136496 243728 136524
rect 231728 136484 231734 136496
rect 243722 136484 243728 136496
rect 243780 136484 243786 136536
rect 282822 136484 282828 136536
rect 282880 136524 282886 136536
rect 292666 136524 292672 136536
rect 282880 136496 292672 136524
rect 282880 136484 282886 136496
rect 292666 136484 292672 136496
rect 292724 136484 292730 136536
rect 260190 135396 260196 135448
rect 260248 135436 260254 135448
rect 265158 135436 265164 135448
rect 260248 135408 265164 135436
rect 260248 135396 260254 135408
rect 265158 135396 265164 135408
rect 265216 135396 265222 135448
rect 203610 135328 203616 135380
rect 203668 135368 203674 135380
rect 214006 135368 214012 135380
rect 203668 135340 214012 135368
rect 203668 135328 203674 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 243538 135328 243544 135380
rect 243596 135368 243602 135380
rect 265802 135368 265808 135380
rect 243596 135340 265808 135368
rect 243596 135328 243602 135340
rect 265802 135328 265808 135340
rect 265860 135328 265866 135380
rect 185670 135260 185676 135312
rect 185728 135300 185734 135312
rect 213914 135300 213920 135312
rect 185728 135272 213920 135300
rect 185728 135260 185734 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 229738 135260 229744 135312
rect 229796 135300 229802 135312
rect 265986 135300 265992 135312
rect 229796 135272 265992 135300
rect 229796 135260 229802 135272
rect 265986 135260 265992 135272
rect 266044 135260 266050 135312
rect 231762 135192 231768 135244
rect 231820 135232 231826 135244
rect 261478 135232 261484 135244
rect 231820 135204 261484 135232
rect 231820 135192 231826 135204
rect 261478 135192 261484 135204
rect 261536 135192 261542 135244
rect 282730 135192 282736 135244
rect 282788 135232 282794 135244
rect 310514 135232 310520 135244
rect 282788 135204 310520 135232
rect 282788 135192 282794 135204
rect 310514 135192 310520 135204
rect 310572 135192 310578 135244
rect 231670 135124 231676 135176
rect 231728 135164 231734 135176
rect 254578 135164 254584 135176
rect 231728 135136 254584 135164
rect 231728 135124 231734 135136
rect 254578 135124 254584 135136
rect 254636 135124 254642 135176
rect 282822 135124 282828 135176
rect 282880 135164 282886 135176
rect 294046 135164 294052 135176
rect 282880 135136 294052 135164
rect 282880 135124 282886 135136
rect 294046 135124 294052 135136
rect 294104 135124 294110 135176
rect 230750 134172 230756 134224
rect 230808 134212 230814 134224
rect 238110 134212 238116 134224
rect 230808 134184 238116 134212
rect 230808 134172 230814 134184
rect 238110 134172 238116 134184
rect 238168 134172 238174 134224
rect 261662 134036 261668 134088
rect 261720 134076 261726 134088
rect 265802 134076 265808 134088
rect 261720 134048 265808 134076
rect 261720 134036 261726 134048
rect 265802 134036 265808 134048
rect 265860 134036 265866 134088
rect 177482 133968 177488 134020
rect 177540 134008 177546 134020
rect 214006 134008 214012 134020
rect 177540 133980 214012 134008
rect 177540 133968 177546 133980
rect 214006 133968 214012 133980
rect 214064 133968 214070 134020
rect 262950 133968 262956 134020
rect 263008 134008 263014 134020
rect 265250 134008 265256 134020
rect 263008 133980 265256 134008
rect 263008 133968 263014 133980
rect 265250 133968 265256 133980
rect 265308 133968 265314 134020
rect 173158 133900 173164 133952
rect 173216 133940 173222 133952
rect 213914 133940 213920 133952
rect 173216 133912 213920 133940
rect 173216 133900 173222 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 254670 133900 254676 133952
rect 254728 133940 254734 133952
rect 264422 133940 264428 133952
rect 254728 133912 264428 133940
rect 254728 133900 254734 133912
rect 264422 133900 264428 133912
rect 264480 133900 264486 133952
rect 231762 133832 231768 133884
rect 231820 133872 231826 133884
rect 262858 133872 262864 133884
rect 231820 133844 262864 133872
rect 231820 133832 231826 133844
rect 262858 133832 262864 133844
rect 262916 133832 262922 133884
rect 281902 133832 281908 133884
rect 281960 133872 281966 133884
rect 313366 133872 313372 133884
rect 281960 133844 313372 133872
rect 281960 133832 281966 133844
rect 313366 133832 313372 133844
rect 313424 133832 313430 133884
rect 231670 133764 231676 133816
rect 231728 133804 231734 133816
rect 261754 133804 261760 133816
rect 231728 133776 261760 133804
rect 231728 133764 231734 133776
rect 261754 133764 261760 133776
rect 261812 133764 261818 133816
rect 263042 132608 263048 132660
rect 263100 132648 263106 132660
rect 265618 132648 265624 132660
rect 263100 132620 265624 132648
rect 263100 132608 263106 132620
rect 265618 132608 265624 132620
rect 265676 132608 265682 132660
rect 230750 132404 230756 132456
rect 230808 132444 230814 132456
rect 257338 132444 257344 132456
rect 230808 132416 257344 132444
rect 230808 132404 230814 132416
rect 257338 132404 257344 132416
rect 257396 132404 257402 132456
rect 231486 132336 231492 132388
rect 231544 132376 231550 132388
rect 246390 132376 246396 132388
rect 231544 132348 246396 132376
rect 231544 132336 231550 132348
rect 246390 132336 246396 132348
rect 246448 132336 246454 132388
rect 282822 132336 282828 132388
rect 282880 132376 282886 132388
rect 303890 132376 303896 132388
rect 282880 132348 303896 132376
rect 282880 132336 282886 132348
rect 303890 132336 303896 132348
rect 303948 132336 303954 132388
rect 231762 132268 231768 132320
rect 231820 132308 231826 132320
rect 244918 132308 244924 132320
rect 231820 132280 244924 132308
rect 231820 132268 231826 132280
rect 244918 132268 244924 132280
rect 244976 132268 244982 132320
rect 246666 131724 246672 131776
rect 246724 131764 246730 131776
rect 265526 131764 265532 131776
rect 246724 131736 265532 131764
rect 246724 131724 246730 131736
rect 265526 131724 265532 131736
rect 265584 131724 265590 131776
rect 191190 131180 191196 131232
rect 191248 131220 191254 131232
rect 214006 131220 214012 131232
rect 191248 131192 214012 131220
rect 191248 131180 191254 131192
rect 214006 131180 214012 131192
rect 214064 131180 214070 131232
rect 175918 131112 175924 131164
rect 175976 131152 175982 131164
rect 213914 131152 213920 131164
rect 175976 131124 213920 131152
rect 175976 131112 175982 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 246482 131112 246488 131164
rect 246540 131152 246546 131164
rect 265710 131152 265716 131164
rect 246540 131124 265716 131152
rect 246540 131112 246546 131124
rect 265710 131112 265716 131124
rect 265768 131112 265774 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 258902 131084 258908 131096
rect 231820 131056 258908 131084
rect 231820 131044 231826 131056
rect 258902 131044 258908 131056
rect 258960 131044 258966 131096
rect 231394 130976 231400 131028
rect 231452 131016 231458 131028
rect 242434 131016 242440 131028
rect 231452 130988 242440 131016
rect 231452 130976 231458 130988
rect 242434 130976 242440 130988
rect 242492 130976 242498 131028
rect 231486 130908 231492 130960
rect 231544 130948 231550 130960
rect 239674 130948 239680 130960
rect 231544 130920 239680 130948
rect 231544 130908 231550 130920
rect 239674 130908 239680 130920
rect 239732 130908 239738 130960
rect 282270 130432 282276 130484
rect 282328 130472 282334 130484
rect 288710 130472 288716 130484
rect 282328 130444 288716 130472
rect 282328 130432 282334 130444
rect 288710 130432 288716 130444
rect 288768 130432 288774 130484
rect 281718 130092 281724 130144
rect 281776 130132 281782 130144
rect 285858 130132 285864 130144
rect 281776 130104 285864 130132
rect 281776 130092 281782 130104
rect 285858 130092 285864 130104
rect 285916 130092 285922 130144
rect 257430 129820 257436 129872
rect 257488 129860 257494 129872
rect 261294 129860 261300 129872
rect 257488 129832 261300 129860
rect 257488 129820 257494 129832
rect 261294 129820 261300 129832
rect 261352 129820 261358 129872
rect 174538 129752 174544 129804
rect 174596 129792 174602 129804
rect 213914 129792 213920 129804
rect 174596 129764 213920 129792
rect 174596 129752 174602 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 239490 129752 239496 129804
rect 239548 129792 239554 129804
rect 264422 129792 264428 129804
rect 239548 129764 264428 129792
rect 239548 129752 239554 129764
rect 264422 129752 264428 129764
rect 264480 129752 264486 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 256234 129724 256240 129736
rect 231820 129696 256240 129724
rect 231820 129684 231826 129696
rect 256234 129684 256240 129696
rect 256292 129684 256298 129736
rect 231670 129616 231676 129668
rect 231728 129656 231734 129668
rect 239766 129656 239772 129668
rect 231728 129628 239772 129656
rect 231728 129616 231734 129628
rect 239766 129616 239772 129628
rect 239824 129616 239830 129668
rect 282822 129208 282828 129260
rect 282880 129248 282886 129260
rect 288526 129248 288532 129260
rect 282880 129220 288532 129248
rect 282880 129208 282886 129220
rect 288526 129208 288532 129220
rect 288584 129208 288590 129260
rect 256050 128460 256056 128512
rect 256108 128500 256114 128512
rect 264422 128500 264428 128512
rect 256108 128472 264428 128500
rect 256108 128460 256114 128472
rect 264422 128460 264428 128472
rect 264480 128460 264486 128512
rect 247770 128392 247776 128444
rect 247828 128432 247834 128444
rect 265802 128432 265808 128444
rect 247828 128404 265808 128432
rect 247828 128392 247834 128404
rect 265802 128392 265808 128404
rect 265860 128392 265866 128444
rect 171962 128324 171968 128376
rect 172020 128364 172026 128376
rect 213914 128364 213920 128376
rect 172020 128336 213920 128364
rect 172020 128324 172026 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 235350 128324 235356 128376
rect 235408 128364 235414 128376
rect 265342 128364 265348 128376
rect 235408 128336 265348 128364
rect 235408 128324 235414 128336
rect 265342 128324 265348 128336
rect 265400 128324 265406 128376
rect 230750 128256 230756 128308
rect 230808 128296 230814 128308
rect 250530 128296 250536 128308
rect 230808 128268 250536 128296
rect 230808 128256 230814 128268
rect 250530 128256 250536 128268
rect 250588 128256 250594 128308
rect 231762 128188 231768 128240
rect 231820 128228 231826 128240
rect 249058 128228 249064 128240
rect 231820 128200 249064 128228
rect 231820 128188 231826 128200
rect 249058 128188 249064 128200
rect 249116 128188 249122 128240
rect 231670 128120 231676 128172
rect 231728 128160 231734 128172
rect 243630 128160 243636 128172
rect 231728 128132 243636 128160
rect 231728 128120 231734 128132
rect 243630 128120 243636 128132
rect 243688 128120 243694 128172
rect 281902 127916 281908 127968
rect 281960 127956 281966 127968
rect 285766 127956 285772 127968
rect 281960 127928 285772 127956
rect 281960 127916 281966 127928
rect 285766 127916 285772 127928
rect 285824 127916 285830 127968
rect 250438 127032 250444 127084
rect 250496 127072 250502 127084
rect 265342 127072 265348 127084
rect 250496 127044 265348 127072
rect 250496 127032 250502 127044
rect 265342 127032 265348 127044
rect 265400 127032 265406 127084
rect 192478 126964 192484 127016
rect 192536 127004 192542 127016
rect 213914 127004 213920 127016
rect 192536 126976 213920 127004
rect 192536 126964 192542 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 249150 126964 249156 127016
rect 249208 127004 249214 127016
rect 264422 127004 264428 127016
rect 249208 126976 264428 127004
rect 249208 126964 249214 126976
rect 264422 126964 264428 126976
rect 264480 126964 264486 127016
rect 231762 126896 231768 126948
rect 231820 126936 231826 126948
rect 246298 126936 246304 126948
rect 231820 126908 246304 126936
rect 231820 126896 231826 126908
rect 246298 126896 246304 126908
rect 246356 126896 246362 126948
rect 282822 126896 282828 126948
rect 282880 126936 282886 126948
rect 302234 126936 302240 126948
rect 282880 126908 302240 126936
rect 282880 126896 282886 126908
rect 302234 126896 302240 126908
rect 302292 126896 302298 126948
rect 467098 126896 467104 126948
rect 467156 126936 467162 126948
rect 580166 126936 580172 126948
rect 467156 126908 580172 126936
rect 467156 126896 467162 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 231578 125808 231584 125860
rect 231636 125848 231642 125860
rect 234062 125848 234068 125860
rect 231636 125820 234068 125848
rect 231636 125808 231642 125820
rect 234062 125808 234068 125820
rect 234120 125808 234126 125860
rect 256234 125740 256240 125792
rect 256292 125780 256298 125792
rect 265710 125780 265716 125792
rect 256292 125752 265716 125780
rect 256292 125740 256298 125752
rect 265710 125740 265716 125752
rect 265768 125740 265774 125792
rect 180334 125672 180340 125724
rect 180392 125712 180398 125724
rect 214006 125712 214012 125724
rect 180392 125684 214012 125712
rect 180392 125672 180398 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 253290 125672 253296 125724
rect 253348 125712 253354 125724
rect 265802 125712 265808 125724
rect 253348 125684 265808 125712
rect 253348 125672 253354 125684
rect 265802 125672 265808 125684
rect 265860 125672 265866 125724
rect 166258 125604 166264 125656
rect 166316 125644 166322 125656
rect 213914 125644 213920 125656
rect 166316 125616 213920 125644
rect 166316 125604 166322 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 238110 125604 238116 125656
rect 238168 125644 238174 125656
rect 265618 125644 265624 125656
rect 238168 125616 265624 125644
rect 238168 125604 238174 125616
rect 265618 125604 265624 125616
rect 265676 125604 265682 125656
rect 231486 125536 231492 125588
rect 231544 125576 231550 125588
rect 255958 125576 255964 125588
rect 231544 125548 255964 125576
rect 231544 125536 231550 125548
rect 255958 125536 255964 125548
rect 256016 125536 256022 125588
rect 282730 125536 282736 125588
rect 282788 125576 282794 125588
rect 303706 125576 303712 125588
rect 282788 125548 303712 125576
rect 282788 125536 282794 125548
rect 303706 125536 303712 125548
rect 303764 125536 303770 125588
rect 231762 125468 231768 125520
rect 231820 125508 231826 125520
rect 240778 125508 240784 125520
rect 231820 125480 240784 125508
rect 231820 125468 231826 125480
rect 240778 125468 240784 125480
rect 240836 125468 240842 125520
rect 282822 125468 282828 125520
rect 282880 125508 282886 125520
rect 290090 125508 290096 125520
rect 282880 125480 290096 125508
rect 282880 125468 282886 125480
rect 290090 125468 290096 125480
rect 290148 125468 290154 125520
rect 230658 124856 230664 124908
rect 230716 124896 230722 124908
rect 246574 124896 246580 124908
rect 230716 124868 246580 124896
rect 230716 124856 230722 124868
rect 246574 124856 246580 124868
rect 246632 124856 246638 124908
rect 261478 124312 261484 124364
rect 261536 124352 261542 124364
rect 265526 124352 265532 124364
rect 261536 124324 265532 124352
rect 261536 124312 261542 124324
rect 265526 124312 265532 124324
rect 265584 124312 265590 124364
rect 200758 124244 200764 124296
rect 200816 124284 200822 124296
rect 213914 124284 213920 124296
rect 200816 124256 213920 124284
rect 200816 124244 200822 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 251818 124244 251824 124296
rect 251876 124284 251882 124296
rect 265802 124284 265808 124296
rect 251876 124256 265808 124284
rect 251876 124244 251882 124256
rect 265802 124244 265808 124256
rect 265860 124244 265866 124296
rect 60642 124176 60648 124228
rect 60700 124216 60706 124228
rect 65518 124216 65524 124228
rect 60700 124188 65524 124216
rect 60700 124176 60706 124188
rect 65518 124176 65524 124188
rect 65576 124176 65582 124228
rect 170674 124176 170680 124228
rect 170732 124216 170738 124228
rect 214006 124216 214012 124228
rect 170732 124188 214012 124216
rect 170732 124176 170738 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 244918 124176 244924 124228
rect 244976 124216 244982 124228
rect 265894 124216 265900 124228
rect 244976 124188 265900 124216
rect 244976 124176 244982 124188
rect 265894 124176 265900 124188
rect 265952 124176 265958 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 242158 124148 242164 124160
rect 231820 124120 242164 124148
rect 231820 124108 231826 124120
rect 242158 124108 242164 124120
rect 242216 124108 242222 124160
rect 281994 123972 282000 124024
rect 282052 124012 282058 124024
rect 284570 124012 284576 124024
rect 282052 123984 284576 124012
rect 282052 123972 282058 123984
rect 284570 123972 284576 123984
rect 284628 123972 284634 124024
rect 170398 123428 170404 123480
rect 170456 123468 170462 123480
rect 202230 123468 202236 123480
rect 170456 123440 202236 123468
rect 170456 123428 170462 123440
rect 202230 123428 202236 123440
rect 202288 123428 202294 123480
rect 231394 123428 231400 123480
rect 231452 123468 231458 123480
rect 263134 123468 263140 123480
rect 231452 123440 263140 123468
rect 231452 123428 231458 123440
rect 263134 123428 263140 123440
rect 263192 123428 263198 123480
rect 260098 122952 260104 123004
rect 260156 122992 260162 123004
rect 264422 122992 264428 123004
rect 260156 122964 264428 122992
rect 260156 122952 260162 122964
rect 264422 122952 264428 122964
rect 264480 122952 264486 123004
rect 173250 122884 173256 122936
rect 173308 122924 173314 122936
rect 214006 122924 214012 122936
rect 173308 122896 214012 122924
rect 173308 122884 173314 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 262858 122884 262864 122936
rect 262916 122924 262922 122936
rect 265802 122924 265808 122936
rect 262916 122896 265808 122924
rect 262916 122884 262922 122896
rect 265802 122884 265808 122896
rect 265860 122884 265866 122936
rect 62022 122816 62028 122868
rect 62080 122856 62086 122868
rect 66070 122856 66076 122868
rect 62080 122828 66076 122856
rect 62080 122816 62086 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 167822 122816 167828 122868
rect 167880 122856 167886 122868
rect 213914 122856 213920 122868
rect 167880 122828 213920 122856
rect 167880 122816 167886 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 232498 122816 232504 122868
rect 232556 122856 232562 122868
rect 265894 122856 265900 122868
rect 232556 122828 265900 122856
rect 232556 122816 232562 122828
rect 265894 122816 265900 122828
rect 265952 122816 265958 122868
rect 230934 122748 230940 122800
rect 230992 122788 230998 122800
rect 258718 122788 258724 122800
rect 230992 122760 258724 122788
rect 230992 122748 230998 122760
rect 258718 122748 258724 122760
rect 258776 122748 258782 122800
rect 282086 122748 282092 122800
rect 282144 122788 282150 122800
rect 304994 122788 305000 122800
rect 282144 122760 305000 122788
rect 282144 122748 282150 122760
rect 304994 122748 305000 122760
rect 305052 122748 305058 122800
rect 231762 122680 231768 122732
rect 231820 122720 231826 122732
rect 246666 122720 246672 122732
rect 231820 122692 246672 122720
rect 231820 122680 231826 122692
rect 246666 122680 246672 122692
rect 246724 122680 246730 122732
rect 282822 122680 282828 122732
rect 282880 122720 282886 122732
rect 291286 122720 291292 122732
rect 282880 122692 291292 122720
rect 282880 122680 282886 122692
rect 291286 122680 291292 122692
rect 291344 122680 291350 122732
rect 231486 122612 231492 122664
rect 231544 122652 231550 122664
rect 241054 122652 241060 122664
rect 231544 122624 241060 122652
rect 231544 122612 231550 122624
rect 241054 122612 241060 122624
rect 241112 122612 241118 122664
rect 258902 121592 258908 121644
rect 258960 121632 258966 121644
rect 264422 121632 264428 121644
rect 258960 121604 264428 121632
rect 258960 121592 258966 121604
rect 264422 121592 264428 121604
rect 264480 121592 264486 121644
rect 184382 121524 184388 121576
rect 184440 121564 184446 121576
rect 214006 121564 214012 121576
rect 184440 121536 214012 121564
rect 184440 121524 184446 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 257338 121524 257344 121576
rect 257396 121564 257402 121576
rect 265894 121564 265900 121576
rect 257396 121536 265900 121564
rect 257396 121524 257402 121536
rect 265894 121524 265900 121536
rect 265952 121524 265958 121576
rect 177574 121456 177580 121508
rect 177632 121496 177638 121508
rect 213914 121496 213920 121508
rect 177632 121468 213920 121496
rect 177632 121456 177638 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 240778 121456 240784 121508
rect 240836 121496 240842 121508
rect 265802 121496 265808 121508
rect 240836 121468 265808 121496
rect 240836 121456 240842 121468
rect 265802 121456 265808 121468
rect 265860 121456 265866 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 253382 121428 253388 121440
rect 231820 121400 253388 121428
rect 231820 121388 231826 121400
rect 253382 121388 253388 121400
rect 253440 121388 253446 121440
rect 282730 121388 282736 121440
rect 282788 121428 282794 121440
rect 300946 121428 300952 121440
rect 282788 121400 300952 121428
rect 282788 121388 282794 121400
rect 300946 121388 300952 121400
rect 301004 121388 301010 121440
rect 231302 121320 231308 121372
rect 231360 121360 231366 121372
rect 247678 121360 247684 121372
rect 231360 121332 247684 121360
rect 231360 121320 231366 121332
rect 247678 121320 247684 121332
rect 247736 121320 247742 121372
rect 282822 121320 282828 121372
rect 282880 121360 282886 121372
rect 299566 121360 299572 121372
rect 282880 121332 299572 121360
rect 282880 121320 282886 121332
rect 299566 121320 299572 121332
rect 299624 121320 299630 121372
rect 231486 121252 231492 121304
rect 231544 121292 231550 121304
rect 242342 121292 242348 121304
rect 231544 121264 242348 121292
rect 231544 121252 231550 121264
rect 242342 121252 242348 121264
rect 242400 121252 242406 121304
rect 254578 120232 254584 120284
rect 254636 120272 254642 120284
rect 265802 120272 265808 120284
rect 254636 120244 265808 120272
rect 254636 120232 254642 120244
rect 265802 120232 265808 120244
rect 265860 120232 265866 120284
rect 178770 120164 178776 120216
rect 178828 120204 178834 120216
rect 214006 120204 214012 120216
rect 178828 120176 214012 120204
rect 178828 120164 178834 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 249058 120164 249064 120216
rect 249116 120204 249122 120216
rect 265894 120204 265900 120216
rect 249116 120176 265900 120204
rect 249116 120164 249122 120176
rect 265894 120164 265900 120176
rect 265952 120164 265958 120216
rect 173434 120096 173440 120148
rect 173492 120136 173498 120148
rect 213914 120136 213920 120148
rect 173492 120108 213920 120136
rect 173492 120096 173498 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 242434 120096 242440 120148
rect 242492 120136 242498 120148
rect 265986 120136 265992 120148
rect 242492 120108 265992 120136
rect 242492 120096 242498 120108
rect 265986 120096 265992 120108
rect 266044 120096 266050 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 247862 120068 247868 120080
rect 231820 120040 247868 120068
rect 231820 120028 231826 120040
rect 247862 120028 247868 120040
rect 247920 120028 247926 120080
rect 282822 120028 282828 120080
rect 282880 120068 282886 120080
rect 306466 120068 306472 120080
rect 282880 120040 306472 120068
rect 282880 120028 282886 120040
rect 306466 120028 306472 120040
rect 306524 120028 306530 120080
rect 231302 119960 231308 120012
rect 231360 120000 231366 120012
rect 245010 120000 245016 120012
rect 231360 119972 245016 120000
rect 231360 119960 231366 119972
rect 245010 119960 245016 119972
rect 245068 119960 245074 120012
rect 177298 119348 177304 119400
rect 177356 119388 177362 119400
rect 195330 119388 195336 119400
rect 177356 119360 195336 119388
rect 177356 119348 177362 119360
rect 195330 119348 195336 119360
rect 195388 119348 195394 119400
rect 238386 119348 238392 119400
rect 238444 119388 238450 119400
rect 265526 119388 265532 119400
rect 238444 119360 265532 119388
rect 238444 119348 238450 119360
rect 265526 119348 265532 119360
rect 265584 119348 265590 119400
rect 177666 118804 177672 118856
rect 177724 118844 177730 118856
rect 213914 118844 213920 118856
rect 177724 118816 213920 118844
rect 177724 118804 177730 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 246298 118804 246304 118856
rect 246356 118844 246362 118856
rect 265526 118844 265532 118856
rect 246356 118816 265532 118844
rect 246356 118804 246362 118816
rect 265526 118804 265532 118816
rect 265584 118804 265590 118856
rect 209222 118736 209228 118788
rect 209280 118776 209286 118788
rect 214006 118776 214012 118788
rect 209280 118748 214012 118776
rect 209280 118736 209286 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 247678 118736 247684 118788
rect 247736 118776 247742 118788
rect 265618 118776 265624 118788
rect 247736 118748 265624 118776
rect 247736 118736 247742 118748
rect 265618 118736 265624 118748
rect 265676 118736 265682 118788
rect 231394 118600 231400 118652
rect 231452 118640 231458 118652
rect 256142 118640 256148 118652
rect 231452 118612 256148 118640
rect 231452 118600 231458 118612
rect 256142 118600 256148 118612
rect 256200 118600 256206 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 296806 118640 296812 118652
rect 282880 118612 296812 118640
rect 282880 118600 282886 118612
rect 296806 118600 296812 118612
rect 296864 118600 296870 118652
rect 281902 118532 281908 118584
rect 281960 118572 281966 118584
rect 284386 118572 284392 118584
rect 281960 118544 284392 118572
rect 281960 118532 281966 118544
rect 284386 118532 284392 118544
rect 284444 118532 284450 118584
rect 231394 117784 231400 117836
rect 231452 117824 231458 117836
rect 235626 117824 235632 117836
rect 231452 117796 235632 117824
rect 231452 117784 231458 117796
rect 235626 117784 235632 117796
rect 235684 117784 235690 117836
rect 255958 117444 255964 117496
rect 256016 117484 256022 117496
rect 265986 117484 265992 117496
rect 256016 117456 265992 117484
rect 256016 117444 256022 117456
rect 265986 117444 265992 117456
rect 266044 117444 266050 117496
rect 210418 117376 210424 117428
rect 210476 117416 210482 117428
rect 214006 117416 214012 117428
rect 210476 117388 214012 117416
rect 210476 117376 210482 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 246390 117376 246396 117428
rect 246448 117416 246454 117428
rect 265894 117416 265900 117428
rect 246448 117388 265900 117416
rect 246448 117376 246454 117388
rect 265894 117376 265900 117388
rect 265952 117376 265958 117428
rect 207658 117308 207664 117360
rect 207716 117348 207722 117360
rect 213914 117348 213920 117360
rect 207716 117320 213920 117348
rect 207716 117308 207722 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 235258 117308 235264 117360
rect 235316 117348 235322 117360
rect 265158 117348 265164 117360
rect 235316 117320 265164 117348
rect 235316 117308 235322 117320
rect 265158 117308 265164 117320
rect 265216 117308 265222 117360
rect 230658 117240 230664 117292
rect 230716 117280 230722 117292
rect 245102 117280 245108 117292
rect 230716 117252 245108 117280
rect 230716 117240 230722 117252
rect 245102 117240 245108 117252
rect 245160 117240 245166 117292
rect 282178 117240 282184 117292
rect 282236 117280 282242 117292
rect 306650 117280 306656 117292
rect 282236 117252 306656 117280
rect 282236 117240 282242 117252
rect 306650 117240 306656 117252
rect 306708 117240 306714 117292
rect 231486 117172 231492 117224
rect 231544 117212 231550 117224
rect 239582 117212 239588 117224
rect 231544 117184 239588 117212
rect 231544 117172 231550 117184
rect 239582 117172 239588 117184
rect 239640 117172 239646 117224
rect 282822 117172 282828 117224
rect 282880 117212 282886 117224
rect 305086 117212 305092 117224
rect 282880 117184 305092 117212
rect 282880 117172 282886 117184
rect 305086 117172 305092 117184
rect 305144 117172 305150 117224
rect 231118 117104 231124 117156
rect 231176 117144 231182 117156
rect 233970 117144 233976 117156
rect 231176 117116 233976 117144
rect 231176 117104 231182 117116
rect 233970 117104 233976 117116
rect 234028 117104 234034 117156
rect 169662 116560 169668 116612
rect 169720 116600 169726 116612
rect 203518 116600 203524 116612
rect 169720 116572 203524 116600
rect 169720 116560 169726 116572
rect 203518 116560 203524 116572
rect 203576 116560 203582 116612
rect 258994 116084 259000 116136
rect 259052 116124 259058 116136
rect 265526 116124 265532 116136
rect 259052 116096 265532 116124
rect 259052 116084 259058 116096
rect 265526 116084 265532 116096
rect 265584 116084 265590 116136
rect 181530 116016 181536 116068
rect 181588 116056 181594 116068
rect 214006 116056 214012 116068
rect 181588 116028 214012 116056
rect 181588 116016 181594 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 245010 116016 245016 116068
rect 245068 116056 245074 116068
rect 265618 116056 265624 116068
rect 245068 116028 265624 116056
rect 245068 116016 245074 116028
rect 265618 116016 265624 116028
rect 265676 116016 265682 116068
rect 169294 115948 169300 116000
rect 169352 115988 169358 116000
rect 213914 115988 213920 116000
rect 169352 115960 213920 115988
rect 169352 115948 169358 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 234062 115948 234068 116000
rect 234120 115988 234126 116000
rect 264422 115988 264428 116000
rect 234120 115960 264428 115988
rect 234120 115948 234126 115960
rect 264422 115948 264428 115960
rect 264480 115948 264486 116000
rect 281718 115880 281724 115932
rect 281776 115920 281782 115932
rect 302418 115920 302424 115932
rect 281776 115892 302424 115920
rect 281776 115880 281782 115892
rect 302418 115880 302424 115892
rect 302476 115880 302482 115932
rect 282086 115812 282092 115864
rect 282144 115852 282150 115864
rect 298738 115852 298744 115864
rect 282144 115824 298744 115852
rect 282144 115812 282150 115824
rect 298738 115812 298744 115824
rect 298796 115812 298802 115864
rect 231210 115472 231216 115524
rect 231268 115512 231274 115524
rect 238018 115512 238024 115524
rect 231268 115484 238024 115512
rect 231268 115472 231274 115484
rect 238018 115472 238024 115484
rect 238076 115472 238082 115524
rect 230566 115200 230572 115252
rect 230624 115240 230630 115252
rect 259086 115240 259092 115252
rect 230624 115212 259092 115240
rect 230624 115200 230630 115212
rect 259086 115200 259092 115212
rect 259144 115200 259150 115252
rect 260282 114588 260288 114640
rect 260340 114628 260346 114640
rect 265434 114628 265440 114640
rect 260340 114600 265440 114628
rect 260340 114588 260346 114600
rect 265434 114588 265440 114600
rect 265492 114588 265498 114640
rect 172054 114520 172060 114572
rect 172112 114560 172118 114572
rect 213914 114560 213920 114572
rect 172112 114532 213920 114560
rect 172112 114520 172118 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 243630 114520 243636 114572
rect 243688 114560 243694 114572
rect 265618 114560 265624 114572
rect 243688 114532 265624 114560
rect 243688 114520 243694 114532
rect 265618 114520 265624 114532
rect 265676 114520 265682 114572
rect 231762 114452 231768 114504
rect 231820 114492 231826 114504
rect 240962 114492 240968 114504
rect 231820 114464 240968 114492
rect 231820 114452 231826 114464
rect 240962 114452 240968 114464
rect 241020 114452 241026 114504
rect 282270 114452 282276 114504
rect 282328 114492 282334 114504
rect 303798 114492 303804 114504
rect 282328 114464 303804 114492
rect 282328 114452 282334 114464
rect 303798 114452 303804 114464
rect 303856 114452 303862 114504
rect 231486 114384 231492 114436
rect 231544 114424 231550 114436
rect 239398 114424 239404 114436
rect 231544 114396 239404 114424
rect 231544 114384 231550 114396
rect 239398 114384 239404 114396
rect 239456 114384 239462 114436
rect 282638 114384 282644 114436
rect 282696 114424 282702 114436
rect 292574 114424 292580 114436
rect 282696 114396 292580 114424
rect 282696 114384 282702 114396
rect 292574 114384 292580 114396
rect 292632 114384 292638 114436
rect 168190 113636 168196 113688
rect 168248 113676 168254 113688
rect 173342 113676 173348 113688
rect 168248 113648 173348 113676
rect 168248 113636 168254 113648
rect 173342 113636 173348 113648
rect 173400 113636 173406 113688
rect 250622 113296 250628 113348
rect 250680 113336 250686 113348
rect 265526 113336 265532 113348
rect 250680 113308 265532 113336
rect 250680 113296 250686 113308
rect 265526 113296 265532 113308
rect 265584 113296 265590 113348
rect 188522 113228 188528 113280
rect 188580 113268 188586 113280
rect 213914 113268 213920 113280
rect 188580 113240 213920 113268
rect 188580 113228 188586 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 242342 113228 242348 113280
rect 242400 113268 242406 113280
rect 265434 113268 265440 113280
rect 242400 113240 265440 113268
rect 242400 113228 242406 113240
rect 265434 113228 265440 113240
rect 265492 113228 265498 113280
rect 174814 113160 174820 113212
rect 174872 113200 174878 113212
rect 214006 113200 214012 113212
rect 174872 113172 214012 113200
rect 174872 113160 174878 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 229830 113160 229836 113212
rect 229888 113200 229894 113212
rect 265894 113200 265900 113212
rect 229888 113172 265900 113200
rect 229888 113160 229894 113172
rect 265894 113160 265900 113172
rect 265952 113160 265958 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 258810 113132 258816 113144
rect 231820 113104 258816 113132
rect 231820 113092 231826 113104
rect 258810 113092 258816 113104
rect 258868 113092 258874 113144
rect 282086 113092 282092 113144
rect 282144 113132 282150 113144
rect 295334 113132 295340 113144
rect 282144 113104 295340 113132
rect 282144 113092 282150 113104
rect 295334 113092 295340 113104
rect 295392 113092 295398 113144
rect 231670 112820 231676 112872
rect 231728 112860 231734 112872
rect 238202 112860 238208 112872
rect 231728 112832 238208 112860
rect 231728 112820 231734 112832
rect 238202 112820 238208 112832
rect 238260 112820 238266 112872
rect 231118 112412 231124 112464
rect 231176 112452 231182 112464
rect 243814 112452 243820 112464
rect 231176 112424 243820 112452
rect 231176 112412 231182 112424
rect 243814 112412 243820 112424
rect 243872 112412 243878 112464
rect 258718 111936 258724 111988
rect 258776 111976 258782 111988
rect 265618 111976 265624 111988
rect 258776 111948 265624 111976
rect 258776 111936 258782 111948
rect 265618 111936 265624 111948
rect 265676 111936 265682 111988
rect 169202 111868 169208 111920
rect 169260 111908 169266 111920
rect 214006 111908 214012 111920
rect 169260 111880 214012 111908
rect 169260 111868 169266 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 253382 111868 253388 111920
rect 253440 111908 253446 111920
rect 265894 111908 265900 111920
rect 253440 111880 265900 111908
rect 253440 111868 253446 111880
rect 265894 111868 265900 111880
rect 265952 111868 265958 111920
rect 166350 111800 166356 111852
rect 166408 111840 166414 111852
rect 213914 111840 213920 111852
rect 166408 111812 213920 111840
rect 166408 111800 166414 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 239398 111800 239404 111852
rect 239456 111840 239462 111852
rect 265526 111840 265532 111852
rect 239456 111812 265532 111840
rect 239456 111800 239462 111812
rect 265526 111800 265532 111812
rect 265584 111800 265590 111852
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 11698 111772 11704 111784
rect 3476 111744 11704 111772
rect 3476 111732 3482 111744
rect 11698 111732 11704 111744
rect 11756 111732 11762 111784
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 169110 111772 169116 111784
rect 168340 111744 169116 111772
rect 168340 111732 168346 111744
rect 169110 111732 169116 111744
rect 169168 111732 169174 111784
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 264330 111772 264336 111784
rect 231820 111744 264336 111772
rect 231820 111732 231826 111744
rect 264330 111732 264336 111744
rect 264388 111732 264394 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 298094 111772 298100 111784
rect 282880 111744 298100 111772
rect 282880 111732 282886 111744
rect 298094 111732 298100 111744
rect 298152 111732 298158 111784
rect 231670 111664 231676 111716
rect 231728 111704 231734 111716
rect 236914 111704 236920 111716
rect 231728 111676 236920 111704
rect 231728 111664 231734 111676
rect 236914 111664 236920 111676
rect 236972 111664 236978 111716
rect 230934 111120 230940 111172
rect 230992 111160 230998 111172
rect 235442 111160 235448 111172
rect 230992 111132 235448 111160
rect 230992 111120 230998 111132
rect 235442 111120 235448 111132
rect 235500 111120 235506 111172
rect 238202 110576 238208 110628
rect 238260 110616 238266 110628
rect 265894 110616 265900 110628
rect 238260 110588 265900 110616
rect 238260 110576 238266 110588
rect 265894 110576 265900 110588
rect 265952 110576 265958 110628
rect 191282 110508 191288 110560
rect 191340 110548 191346 110560
rect 214006 110548 214012 110560
rect 191340 110520 214012 110548
rect 191340 110508 191346 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 256142 110508 256148 110560
rect 256200 110548 256206 110560
rect 265158 110548 265164 110560
rect 256200 110520 265164 110548
rect 256200 110508 256206 110520
rect 265158 110508 265164 110520
rect 265216 110508 265222 110560
rect 178862 110440 178868 110492
rect 178920 110480 178926 110492
rect 213914 110480 213920 110492
rect 178920 110452 213920 110480
rect 178920 110440 178926 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 231670 110372 231676 110424
rect 231728 110412 231734 110424
rect 260466 110412 260472 110424
rect 231728 110384 260472 110412
rect 231728 110372 231734 110384
rect 260466 110372 260472 110384
rect 260524 110372 260530 110424
rect 282822 110372 282828 110424
rect 282880 110412 282886 110424
rect 291194 110412 291200 110424
rect 282880 110384 291200 110412
rect 282880 110372 282886 110384
rect 291194 110372 291200 110384
rect 291252 110372 291258 110424
rect 231762 110304 231768 110356
rect 231820 110344 231826 110356
rect 253198 110344 253204 110356
rect 231820 110316 253204 110344
rect 231820 110304 231826 110316
rect 253198 110304 253204 110316
rect 253256 110304 253262 110356
rect 231670 109692 231676 109744
rect 231728 109732 231734 109744
rect 236822 109732 236828 109744
rect 231728 109704 236828 109732
rect 231728 109692 231734 109704
rect 236822 109692 236828 109704
rect 236880 109692 236886 109744
rect 260374 109148 260380 109200
rect 260432 109188 260438 109200
rect 265986 109188 265992 109200
rect 260432 109160 265992 109188
rect 260432 109148 260438 109160
rect 265986 109148 265992 109160
rect 266044 109148 266050 109200
rect 188430 109080 188436 109132
rect 188488 109120 188494 109132
rect 213914 109120 213920 109132
rect 188488 109092 213920 109120
rect 188488 109080 188494 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 257614 109080 257620 109132
rect 257672 109120 257678 109132
rect 265894 109120 265900 109132
rect 257672 109092 265900 109120
rect 257672 109080 257678 109092
rect 265894 109080 265900 109092
rect 265952 109080 265958 109132
rect 169110 109012 169116 109064
rect 169168 109052 169174 109064
rect 214006 109052 214012 109064
rect 169168 109024 214012 109052
rect 169168 109012 169174 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 243722 109012 243728 109064
rect 243780 109052 243786 109064
rect 265526 109052 265532 109064
rect 243780 109024 265532 109052
rect 243780 109012 243786 109024
rect 265526 109012 265532 109024
rect 265584 109012 265590 109064
rect 167914 108944 167920 108996
rect 167972 108984 167978 108996
rect 174630 108984 174636 108996
rect 167972 108956 174636 108984
rect 167972 108944 167978 108956
rect 174630 108944 174636 108956
rect 174688 108944 174694 108996
rect 231670 108944 231676 108996
rect 231728 108984 231734 108996
rect 250714 108984 250720 108996
rect 231728 108956 250720 108984
rect 231728 108944 231734 108956
rect 250714 108944 250720 108956
rect 250772 108944 250778 108996
rect 282822 108944 282828 108996
rect 282880 108984 282886 108996
rect 310606 108984 310612 108996
rect 282880 108956 310612 108984
rect 282880 108944 282886 108956
rect 310606 108944 310612 108956
rect 310664 108944 310670 108996
rect 231762 108876 231768 108928
rect 231820 108916 231826 108928
rect 245194 108916 245200 108928
rect 231820 108888 245200 108916
rect 231820 108876 231826 108888
rect 245194 108876 245200 108888
rect 245252 108876 245258 108928
rect 231578 108400 231584 108452
rect 231636 108440 231642 108452
rect 234154 108440 234160 108452
rect 231636 108412 234160 108440
rect 231636 108400 231642 108412
rect 234154 108400 234160 108412
rect 234212 108400 234218 108452
rect 238294 107856 238300 107908
rect 238352 107896 238358 107908
rect 265894 107896 265900 107908
rect 238352 107868 265900 107896
rect 238352 107856 238358 107868
rect 265894 107856 265900 107868
rect 265952 107856 265958 107908
rect 250530 107788 250536 107840
rect 250588 107828 250594 107840
rect 265986 107828 265992 107840
rect 250588 107800 265992 107828
rect 250588 107788 250594 107800
rect 265986 107788 265992 107800
rect 266044 107788 266050 107840
rect 178954 107720 178960 107772
rect 179012 107760 179018 107772
rect 214006 107760 214012 107772
rect 179012 107732 214012 107760
rect 179012 107720 179018 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 245102 107720 245108 107772
rect 245160 107760 245166 107772
rect 264514 107760 264520 107772
rect 245160 107732 264520 107760
rect 245160 107720 245166 107732
rect 264514 107720 264520 107732
rect 264572 107720 264578 107772
rect 174722 107652 174728 107704
rect 174780 107692 174786 107704
rect 213914 107692 213920 107704
rect 174780 107664 213920 107692
rect 174780 107652 174786 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 261754 107652 261760 107704
rect 261812 107692 261818 107704
rect 265342 107692 265348 107704
rect 261812 107664 265348 107692
rect 261812 107652 261818 107664
rect 265342 107652 265348 107664
rect 265400 107652 265406 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 257522 107624 257528 107636
rect 231820 107596 257528 107624
rect 231820 107584 231826 107596
rect 257522 107584 257528 107596
rect 257580 107584 257586 107636
rect 231486 107108 231492 107160
rect 231544 107148 231550 107160
rect 233878 107148 233884 107160
rect 231544 107120 233884 107148
rect 231544 107108 231550 107120
rect 233878 107108 233884 107120
rect 233936 107108 233942 107160
rect 230750 106632 230756 106684
rect 230808 106672 230814 106684
rect 235534 106672 235540 106684
rect 230808 106644 235540 106672
rect 230808 106632 230814 106644
rect 235534 106632 235540 106644
rect 235592 106632 235598 106684
rect 240962 106428 240968 106480
rect 241020 106468 241026 106480
rect 265894 106468 265900 106480
rect 241020 106440 265900 106468
rect 241020 106428 241026 106440
rect 265894 106428 265900 106440
rect 265952 106428 265958 106480
rect 170398 106360 170404 106412
rect 170456 106400 170462 106412
rect 214006 106400 214012 106412
rect 170456 106372 214012 106400
rect 170456 106360 170462 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 249242 106360 249248 106412
rect 249300 106400 249306 106412
rect 265986 106400 265992 106412
rect 249300 106372 265992 106400
rect 249300 106360 249306 106372
rect 265986 106360 265992 106372
rect 266044 106360 266050 106412
rect 167914 106292 167920 106344
rect 167972 106332 167978 106344
rect 213914 106332 213920 106344
rect 167972 106304 213920 106332
rect 167972 106292 167978 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 231486 106224 231492 106276
rect 231544 106264 231550 106276
rect 261570 106264 261576 106276
rect 231544 106236 261576 106264
rect 231544 106224 231550 106236
rect 261570 106224 261576 106236
rect 261628 106224 261634 106276
rect 231762 106156 231768 106208
rect 231820 106196 231826 106208
rect 242250 106196 242256 106208
rect 231820 106168 242256 106196
rect 231820 106156 231826 106168
rect 242250 106156 242256 106168
rect 242308 106156 242314 106208
rect 282822 105068 282828 105120
rect 282880 105108 282886 105120
rect 287238 105108 287244 105120
rect 282880 105080 287244 105108
rect 282880 105068 282886 105080
rect 287238 105068 287244 105080
rect 287296 105068 287302 105120
rect 263134 105000 263140 105052
rect 263192 105040 263198 105052
rect 265250 105040 265256 105052
rect 263192 105012 265256 105040
rect 263192 105000 263198 105012
rect 265250 105000 265256 105012
rect 265308 105000 265314 105052
rect 210602 104932 210608 104984
rect 210660 104972 210666 104984
rect 214006 104972 214012 104984
rect 210660 104944 214012 104972
rect 210660 104932 210666 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 253474 104932 253480 104984
rect 253532 104972 253538 104984
rect 265894 104972 265900 104984
rect 253532 104944 265900 104972
rect 253532 104932 253538 104944
rect 265894 104932 265900 104944
rect 265952 104932 265958 104984
rect 176102 104864 176108 104916
rect 176160 104904 176166 104916
rect 213914 104904 213920 104916
rect 176160 104876 213920 104904
rect 176160 104864 176166 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 242158 104864 242164 104916
rect 242216 104904 242222 104916
rect 265618 104904 265624 104916
rect 242216 104876 265624 104904
rect 242216 104864 242222 104876
rect 265618 104864 265624 104876
rect 265676 104864 265682 104916
rect 230566 104796 230572 104848
rect 230624 104836 230630 104848
rect 232590 104836 232596 104848
rect 230624 104808 232596 104836
rect 230624 104796 230630 104808
rect 232590 104796 232596 104808
rect 232648 104796 232654 104848
rect 230474 104116 230480 104168
rect 230532 104156 230538 104168
rect 254762 104156 254768 104168
rect 230532 104128 254768 104156
rect 230532 104116 230538 104128
rect 254762 104116 254768 104128
rect 254820 104116 254826 104168
rect 258810 103980 258816 104032
rect 258868 104020 258874 104032
rect 265618 104020 265624 104032
rect 258868 103992 265624 104020
rect 258868 103980 258874 103992
rect 265618 103980 265624 103992
rect 265676 103980 265682 104032
rect 247862 103572 247868 103624
rect 247920 103612 247926 103624
rect 265986 103612 265992 103624
rect 247920 103584 265992 103612
rect 247920 103572 247926 103584
rect 265986 103572 265992 103584
rect 266044 103572 266050 103624
rect 206462 103504 206468 103556
rect 206520 103544 206526 103556
rect 213914 103544 213920 103556
rect 206520 103516 213920 103544
rect 206520 103504 206526 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 233970 103504 233976 103556
rect 234028 103544 234034 103556
rect 265894 103544 265900 103556
rect 234028 103516 265900 103544
rect 234028 103504 234034 103516
rect 265894 103504 265900 103516
rect 265952 103504 265958 103556
rect 231578 102756 231584 102808
rect 231636 102796 231642 102808
rect 250806 102796 250812 102808
rect 231636 102768 250812 102796
rect 231636 102756 231642 102768
rect 250806 102756 250812 102768
rect 250864 102756 250870 102808
rect 257522 102280 257528 102332
rect 257580 102320 257586 102332
rect 265342 102320 265348 102332
rect 257580 102292 265348 102320
rect 257580 102280 257586 102292
rect 265342 102280 265348 102292
rect 265400 102280 265406 102332
rect 232590 102212 232596 102264
rect 232648 102252 232654 102264
rect 232648 102224 232912 102252
rect 232648 102212 232654 102224
rect 211890 102144 211896 102196
rect 211948 102184 211954 102196
rect 213914 102184 213920 102196
rect 211948 102156 213920 102184
rect 211948 102144 211954 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 230934 102144 230940 102196
rect 230992 102184 230998 102196
rect 232774 102184 232780 102196
rect 230992 102156 232780 102184
rect 230992 102144 230998 102156
rect 232774 102144 232780 102156
rect 232832 102144 232838 102196
rect 232884 102184 232912 102224
rect 236914 102212 236920 102264
rect 236972 102252 236978 102264
rect 265526 102252 265532 102264
rect 236972 102224 265532 102252
rect 236972 102212 236978 102224
rect 265526 102212 265532 102224
rect 265584 102212 265590 102264
rect 265618 102184 265624 102196
rect 232884 102156 265624 102184
rect 265618 102144 265624 102156
rect 265676 102144 265682 102196
rect 230566 102076 230572 102128
rect 230624 102116 230630 102128
rect 264606 102116 264612 102128
rect 230624 102088 264612 102116
rect 230624 102076 230630 102088
rect 264606 102076 264612 102088
rect 264664 102076 264670 102128
rect 230750 101940 230756 101992
rect 230808 101980 230814 101992
rect 232682 101980 232688 101992
rect 230808 101952 232688 101980
rect 230808 101940 230814 101952
rect 232682 101940 232688 101952
rect 232740 101940 232746 101992
rect 231670 101396 231676 101448
rect 231728 101436 231734 101448
rect 252094 101436 252100 101448
rect 231728 101408 252100 101436
rect 231728 101396 231734 101408
rect 252094 101396 252100 101408
rect 252152 101396 252158 101448
rect 250714 100852 250720 100904
rect 250772 100892 250778 100904
rect 265894 100892 265900 100904
rect 250772 100864 265900 100892
rect 250772 100852 250778 100864
rect 265894 100852 265900 100864
rect 265952 100852 265958 100904
rect 210510 100784 210516 100836
rect 210568 100824 210574 100836
rect 214006 100824 214012 100836
rect 210568 100796 214012 100824
rect 210568 100784 210574 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 252002 100784 252008 100836
rect 252060 100824 252066 100836
rect 265986 100824 265992 100836
rect 252060 100796 265992 100824
rect 252060 100784 252066 100796
rect 265986 100784 265992 100796
rect 266044 100784 266050 100836
rect 200850 100716 200856 100768
rect 200908 100756 200914 100768
rect 213914 100756 213920 100768
rect 200908 100728 213920 100756
rect 200908 100716 200914 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 231486 100648 231492 100700
rect 231544 100688 231550 100700
rect 253566 100688 253572 100700
rect 231544 100660 253572 100688
rect 231544 100648 231550 100660
rect 253566 100648 253572 100660
rect 253624 100648 253630 100700
rect 471238 100648 471244 100700
rect 471296 100688 471302 100700
rect 580166 100688 580172 100700
rect 471296 100660 580172 100688
rect 471296 100648 471302 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 231762 100580 231768 100632
rect 231820 100620 231826 100632
rect 249334 100620 249340 100632
rect 231820 100592 249340 100620
rect 231820 100580 231826 100592
rect 249334 100580 249340 100592
rect 249392 100580 249398 100632
rect 254762 99492 254768 99544
rect 254820 99532 254826 99544
rect 265894 99532 265900 99544
rect 254820 99504 265900 99532
rect 254820 99492 254826 99504
rect 265894 99492 265900 99504
rect 265952 99492 265958 99544
rect 253198 99424 253204 99476
rect 253256 99464 253262 99476
rect 265618 99464 265624 99476
rect 253256 99436 265624 99464
rect 253256 99424 253262 99436
rect 265618 99424 265624 99436
rect 265676 99424 265682 99476
rect 166534 99356 166540 99408
rect 166592 99396 166598 99408
rect 213914 99396 213920 99408
rect 166592 99368 213920 99396
rect 166592 99356 166598 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 246574 99356 246580 99408
rect 246632 99396 246638 99408
rect 265158 99396 265164 99408
rect 246632 99368 265164 99396
rect 246632 99356 246638 99368
rect 265158 99356 265164 99368
rect 265216 99356 265222 99408
rect 231762 99288 231768 99340
rect 231820 99328 231826 99340
rect 267090 99328 267096 99340
rect 231820 99300 267096 99328
rect 231820 99288 231826 99300
rect 267090 99288 267096 99300
rect 267148 99288 267154 99340
rect 231486 98608 231492 98660
rect 231544 98648 231550 98660
rect 238386 98648 238392 98660
rect 231544 98620 238392 98648
rect 231544 98608 231550 98620
rect 238386 98608 238392 98620
rect 238444 98608 238450 98660
rect 166442 98064 166448 98116
rect 166500 98104 166506 98116
rect 214006 98104 214012 98116
rect 166500 98076 214012 98104
rect 166500 98064 166506 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 242250 98064 242256 98116
rect 242308 98104 242314 98116
rect 261202 98104 261208 98116
rect 242308 98076 261208 98104
rect 242308 98064 242314 98076
rect 261202 98064 261208 98076
rect 261260 98064 261266 98116
rect 164878 97996 164884 98048
rect 164936 98036 164942 98048
rect 213914 98036 213920 98048
rect 164936 98008 213920 98036
rect 164936 97996 164942 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 238018 97996 238024 98048
rect 238076 98036 238082 98048
rect 264606 98036 264612 98048
rect 238076 98008 264612 98036
rect 238076 97996 238082 98008
rect 264606 97996 264612 98008
rect 264664 97996 264670 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 14458 97968 14464 97980
rect 3476 97940 14464 97968
rect 3476 97928 3482 97940
rect 14458 97928 14464 97940
rect 14516 97928 14522 97980
rect 236822 96704 236828 96756
rect 236880 96744 236886 96756
rect 265986 96744 265992 96756
rect 236880 96716 265992 96744
rect 236880 96704 236886 96716
rect 265986 96704 265992 96716
rect 266044 96704 266050 96756
rect 231118 96636 231124 96688
rect 231176 96676 231182 96688
rect 265342 96676 265348 96688
rect 231176 96648 265348 96676
rect 231176 96636 231182 96648
rect 265342 96636 265348 96648
rect 265400 96636 265406 96688
rect 209130 96568 209136 96620
rect 209188 96608 209194 96620
rect 229094 96608 229100 96620
rect 209188 96580 229100 96608
rect 209188 96568 209194 96580
rect 229094 96568 229100 96580
rect 229152 96608 229158 96620
rect 230566 96608 230572 96620
rect 229152 96580 230572 96608
rect 229152 96568 229158 96580
rect 230566 96568 230572 96580
rect 230624 96568 230630 96620
rect 189718 96364 189724 96416
rect 189776 96404 189782 96416
rect 281626 96404 281632 96416
rect 189776 96376 281632 96404
rect 189776 96364 189782 96376
rect 281626 96364 281632 96376
rect 281684 96364 281690 96416
rect 231762 95888 231768 95940
rect 231820 95928 231826 95940
rect 268010 95928 268016 95940
rect 231820 95900 268016 95928
rect 231820 95888 231826 95900
rect 268010 95888 268016 95900
rect 268068 95888 268074 95940
rect 228358 95208 228364 95260
rect 228416 95248 228422 95260
rect 265526 95248 265532 95260
rect 228416 95220 265532 95248
rect 228416 95208 228422 95220
rect 265526 95208 265532 95220
rect 265584 95208 265590 95260
rect 184198 95140 184204 95192
rect 184256 95180 184262 95192
rect 281534 95180 281540 95192
rect 184256 95152 281540 95180
rect 184256 95140 184262 95152
rect 281534 95140 281540 95152
rect 281592 95140 281598 95192
rect 199378 95072 199384 95124
rect 199436 95112 199442 95124
rect 281718 95112 281724 95124
rect 199436 95084 281724 95112
rect 199436 95072 199442 95084
rect 281718 95072 281724 95084
rect 281776 95072 281782 95124
rect 216122 95004 216128 95056
rect 216180 95044 216186 95056
rect 279418 95044 279424 95056
rect 216180 95016 279424 95044
rect 216180 95004 216186 95016
rect 279418 95004 279424 95016
rect 279476 95004 279482 95056
rect 222838 94460 222844 94512
rect 222896 94500 222902 94512
rect 267182 94500 267188 94512
rect 222896 94472 267188 94500
rect 222896 94460 222902 94472
rect 267182 94460 267188 94472
rect 267240 94460 267246 94512
rect 133138 94120 133144 94172
rect 133196 94160 133202 94172
rect 171870 94160 171876 94172
rect 133196 94132 171876 94160
rect 133196 94120 133202 94132
rect 171870 94120 171876 94132
rect 171928 94120 171934 94172
rect 120626 94052 120632 94104
rect 120684 94092 120690 94104
rect 167822 94092 167828 94104
rect 120684 94064 167828 94092
rect 120684 94052 120690 94064
rect 167822 94052 167828 94064
rect 167880 94052 167886 94104
rect 104342 93984 104348 94036
rect 104400 94024 104406 94036
rect 174814 94024 174820 94036
rect 104400 93996 174820 94024
rect 104400 93984 104406 93996
rect 174814 93984 174820 93996
rect 174872 93984 174878 94036
rect 116670 93916 116676 93968
rect 116728 93956 116734 93968
rect 192570 93956 192576 93968
rect 116728 93928 192576 93956
rect 116728 93916 116734 93928
rect 192570 93916 192576 93928
rect 192628 93916 192634 93968
rect 94958 93848 94964 93900
rect 95016 93888 95022 93900
rect 178954 93888 178960 93900
rect 95016 93860 178960 93888
rect 95016 93848 95022 93860
rect 178954 93848 178960 93860
rect 179012 93848 179018 93900
rect 230566 93848 230572 93900
rect 230624 93888 230630 93900
rect 234154 93888 234160 93900
rect 230624 93860 234160 93888
rect 230624 93848 230630 93860
rect 234154 93848 234160 93860
rect 234212 93848 234218 93900
rect 268010 93780 268016 93832
rect 268068 93820 268074 93832
rect 276934 93820 276940 93832
rect 268068 93792 276940 93820
rect 268068 93780 268074 93792
rect 276934 93780 276940 93792
rect 276992 93780 276998 93832
rect 234154 93712 234160 93764
rect 234212 93752 234218 93764
rect 270954 93752 270960 93764
rect 234212 93724 270960 93752
rect 234212 93712 234218 93724
rect 270954 93712 270960 93724
rect 271012 93712 271018 93764
rect 151722 93440 151728 93492
rect 151780 93480 151786 93492
rect 167638 93480 167644 93492
rect 151780 93452 167644 93480
rect 151780 93440 151786 93452
rect 167638 93440 167644 93452
rect 167696 93440 167702 93492
rect 122098 93372 122104 93424
rect 122156 93412 122162 93424
rect 170582 93412 170588 93424
rect 122156 93384 170588 93412
rect 122156 93372 122162 93384
rect 170582 93372 170588 93384
rect 170640 93372 170646 93424
rect 115842 93304 115848 93356
rect 115900 93344 115906 93356
rect 173434 93344 173440 93356
rect 115900 93316 173440 93344
rect 115900 93304 115906 93316
rect 173434 93304 173440 93316
rect 173492 93304 173498 93356
rect 107746 93236 107752 93288
rect 107804 93276 107810 93288
rect 169294 93276 169300 93288
rect 107804 93248 169300 93276
rect 107804 93236 107810 93248
rect 169294 93236 169300 93248
rect 169352 93236 169358 93288
rect 85666 93168 85672 93220
rect 85724 93208 85730 93220
rect 164878 93208 164884 93220
rect 85724 93180 164884 93208
rect 85724 93168 85730 93180
rect 164878 93168 164884 93180
rect 164936 93168 164942 93220
rect 129734 93100 129740 93152
rect 129792 93140 129798 93152
rect 214558 93140 214564 93152
rect 129792 93112 214564 93140
rect 129792 93100 129798 93112
rect 214558 93100 214564 93112
rect 214616 93100 214622 93152
rect 217226 93100 217232 93152
rect 217284 93140 217290 93152
rect 277394 93140 277400 93152
rect 217284 93112 277400 93140
rect 217284 93100 217290 93112
rect 277394 93100 277400 93112
rect 277452 93100 277458 93152
rect 230474 92488 230480 92540
rect 230532 92528 230538 92540
rect 233878 92528 233884 92540
rect 230532 92500 233884 92528
rect 230532 92488 230538 92500
rect 233878 92488 233884 92500
rect 233936 92488 233942 92540
rect 114462 92420 114468 92472
rect 114520 92460 114526 92472
rect 203610 92460 203616 92472
rect 114520 92432 203616 92460
rect 114520 92420 114526 92432
rect 203610 92420 203616 92432
rect 203668 92420 203674 92472
rect 105722 92352 105728 92404
rect 105780 92392 105786 92404
rect 191190 92392 191196 92404
rect 105780 92364 191196 92392
rect 105780 92352 105786 92364
rect 191190 92352 191196 92364
rect 191248 92352 191254 92404
rect 120258 92284 120264 92336
rect 120316 92324 120322 92336
rect 181438 92324 181444 92336
rect 120316 92296 181444 92324
rect 120316 92284 120322 92296
rect 181438 92284 181444 92296
rect 181496 92284 181502 92336
rect 123202 92216 123208 92268
rect 123260 92256 123266 92268
rect 176010 92256 176016 92268
rect 123260 92228 176016 92256
rect 123260 92216 123266 92228
rect 176010 92216 176016 92228
rect 176068 92216 176074 92268
rect 106826 92148 106832 92200
rect 106884 92188 106890 92200
rect 129734 92188 129740 92200
rect 106884 92160 129740 92188
rect 106884 92148 106890 92160
rect 129734 92148 129740 92160
rect 129792 92148 129798 92200
rect 134426 92148 134432 92200
rect 134484 92188 134490 92200
rect 167730 92188 167736 92200
rect 134484 92160 167736 92188
rect 134484 92148 134490 92160
rect 167730 92148 167736 92160
rect 167788 92148 167794 92200
rect 152090 92080 152096 92132
rect 152148 92120 152154 92132
rect 171778 92120 171784 92132
rect 152148 92092 171784 92120
rect 152148 92080 152154 92092
rect 171778 92080 171784 92092
rect 171836 92080 171842 92132
rect 188338 91740 188344 91792
rect 188396 91780 188402 91792
rect 276014 91780 276020 91792
rect 188396 91752 276020 91780
rect 188396 91740 188402 91752
rect 276014 91740 276020 91752
rect 276072 91740 276078 91792
rect 99282 91264 99288 91316
rect 99340 91304 99346 91316
rect 106918 91304 106924 91316
rect 99340 91276 106924 91304
rect 99340 91264 99346 91276
rect 106918 91264 106924 91276
rect 106976 91264 106982 91316
rect 100018 91196 100024 91248
rect 100076 91236 100082 91248
rect 123478 91236 123484 91248
rect 100076 91208 123484 91236
rect 100076 91196 100082 91208
rect 123478 91196 123484 91208
rect 123536 91196 123542 91248
rect 88058 91128 88064 91180
rect 88116 91168 88122 91180
rect 120074 91168 120080 91180
rect 88116 91140 120080 91168
rect 88116 91128 88122 91140
rect 120074 91128 120080 91140
rect 120132 91128 120138 91180
rect 85114 91060 85120 91112
rect 85172 91100 85178 91112
rect 133138 91100 133144 91112
rect 85172 91072 133144 91100
rect 85172 91060 85178 91072
rect 133138 91060 133144 91072
rect 133196 91060 133202 91112
rect 67542 90992 67548 91044
rect 67600 91032 67606 91044
rect 214650 91032 214656 91044
rect 67600 91004 214656 91032
rect 67600 90992 67606 91004
rect 214650 90992 214656 91004
rect 214708 90992 214714 91044
rect 180242 90924 180248 90976
rect 180300 90964 180306 90976
rect 280246 90964 280252 90976
rect 180300 90936 280252 90964
rect 180300 90924 180306 90936
rect 280246 90924 280252 90936
rect 280304 90924 280310 90976
rect 120074 90856 120080 90908
rect 120132 90896 120138 90908
rect 214834 90896 214840 90908
rect 120132 90868 214840 90896
rect 120132 90856 120138 90868
rect 214834 90856 214840 90868
rect 214892 90856 214898 90908
rect 124122 90788 124128 90840
rect 124180 90828 124186 90840
rect 170674 90828 170680 90840
rect 124180 90800 170680 90828
rect 124180 90788 124186 90800
rect 170674 90788 170680 90800
rect 170732 90788 170738 90840
rect 125410 90720 125416 90772
rect 125468 90760 125474 90772
rect 166258 90760 166264 90772
rect 125468 90732 166264 90760
rect 125468 90720 125474 90732
rect 166258 90720 166264 90732
rect 166316 90720 166322 90772
rect 109678 90652 109684 90704
rect 109736 90692 109742 90704
rect 181530 90692 181536 90704
rect 109736 90664 181536 90692
rect 109736 90652 109742 90664
rect 181530 90652 181536 90664
rect 181588 90652 181594 90704
rect 67358 89632 67364 89684
rect 67416 89672 67422 89684
rect 210510 89672 210516 89684
rect 67416 89644 210516 89672
rect 67416 89632 67422 89644
rect 210510 89632 210516 89644
rect 210568 89632 210574 89684
rect 126882 89564 126888 89616
rect 126940 89604 126946 89616
rect 195422 89604 195428 89616
rect 126940 89576 195428 89604
rect 126940 89564 126946 89576
rect 195422 89564 195428 89576
rect 195480 89564 195486 89616
rect 101858 89496 101864 89548
rect 101916 89536 101922 89548
rect 169202 89536 169208 89548
rect 101916 89508 169208 89536
rect 101916 89496 101922 89508
rect 169202 89496 169208 89508
rect 169260 89496 169266 89548
rect 112714 89428 112720 89480
rect 112772 89468 112778 89480
rect 177666 89468 177672 89480
rect 112772 89440 177672 89468
rect 112772 89428 112778 89440
rect 177666 89428 177672 89440
rect 177724 89428 177730 89480
rect 119522 89360 119528 89412
rect 119580 89400 119586 89412
rect 170490 89400 170496 89412
rect 119580 89372 170496 89400
rect 119580 89360 119586 89372
rect 170490 89360 170496 89372
rect 170548 89360 170554 89412
rect 136266 89292 136272 89344
rect 136324 89332 136330 89344
rect 187142 89332 187148 89344
rect 136324 89304 187148 89332
rect 136324 89292 136330 89304
rect 187142 89292 187148 89304
rect 187200 89292 187206 89344
rect 196710 88952 196716 89004
rect 196768 88992 196774 89004
rect 265802 88992 265808 89004
rect 196768 88964 265808 88992
rect 196768 88952 196774 88964
rect 265802 88952 265808 88964
rect 265860 88952 265866 89004
rect 89070 88272 89076 88324
rect 89128 88312 89134 88324
rect 166534 88312 166540 88324
rect 89128 88284 166540 88312
rect 89128 88272 89134 88284
rect 166534 88272 166540 88284
rect 166592 88272 166598 88324
rect 122834 88204 122840 88256
rect 122892 88244 122898 88256
rect 200758 88244 200764 88256
rect 122892 88216 200764 88244
rect 122892 88204 122898 88216
rect 200758 88204 200764 88216
rect 200816 88204 200822 88256
rect 107102 88136 107108 88188
rect 107160 88176 107166 88188
rect 172054 88176 172060 88188
rect 107160 88148 172060 88176
rect 107160 88136 107166 88148
rect 172054 88136 172060 88148
rect 172112 88136 172118 88188
rect 151538 88068 151544 88120
rect 151596 88108 151602 88120
rect 211798 88108 211804 88120
rect 151596 88080 211804 88108
rect 151596 88068 151602 88080
rect 211798 88068 211804 88080
rect 211856 88068 211862 88120
rect 118234 88000 118240 88052
rect 118292 88040 118298 88052
rect 177574 88040 177580 88052
rect 118292 88012 177580 88040
rect 118292 88000 118298 88012
rect 177574 88000 177580 88012
rect 177632 88000 177638 88052
rect 129458 87932 129464 87984
rect 129516 87972 129522 87984
rect 182818 87972 182824 87984
rect 129516 87944 182824 87972
rect 129516 87932 129522 87944
rect 182818 87932 182824 87944
rect 182876 87932 182882 87984
rect 105722 86912 105728 86964
rect 105780 86952 105786 86964
rect 213454 86952 213460 86964
rect 105780 86924 213460 86952
rect 105780 86912 105786 86924
rect 213454 86912 213460 86924
rect 213512 86912 213518 86964
rect 90634 86844 90640 86896
rect 90692 86884 90698 86896
rect 176102 86884 176108 86896
rect 90692 86856 176108 86884
rect 90692 86844 90698 86856
rect 176102 86844 176108 86856
rect 176160 86844 176166 86896
rect 119706 86776 119712 86828
rect 119764 86816 119770 86828
rect 184382 86816 184388 86828
rect 119764 86788 184388 86816
rect 119764 86776 119770 86788
rect 184382 86776 184388 86788
rect 184440 86776 184446 86828
rect 151722 86708 151728 86760
rect 151780 86748 151786 86760
rect 196802 86748 196808 86760
rect 151780 86720 196808 86748
rect 151780 86708 151786 86720
rect 196802 86708 196808 86720
rect 196860 86708 196866 86760
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 35158 85524 35164 85536
rect 3200 85496 35164 85524
rect 3200 85484 3206 85496
rect 35158 85484 35164 85496
rect 35216 85484 35222 85536
rect 67634 85484 67640 85536
rect 67692 85524 67698 85536
rect 216214 85524 216220 85536
rect 67692 85496 216220 85524
rect 67692 85484 67698 85496
rect 216214 85484 216220 85496
rect 216272 85484 216278 85536
rect 67726 85416 67732 85468
rect 67784 85456 67790 85468
rect 214742 85456 214748 85468
rect 67784 85428 214748 85456
rect 67784 85416 67790 85428
rect 214742 85416 214748 85428
rect 214800 85416 214806 85468
rect 91922 85348 91928 85400
rect 91980 85388 91986 85400
rect 167914 85388 167920 85400
rect 91980 85360 167920 85388
rect 91980 85348 91986 85360
rect 167914 85348 167920 85360
rect 167972 85348 167978 85400
rect 111058 85280 111064 85332
rect 111116 85320 111122 85332
rect 177482 85320 177488 85332
rect 111116 85292 177488 85320
rect 111116 85280 111122 85292
rect 177482 85280 177488 85292
rect 177540 85280 177546 85332
rect 130746 85212 130752 85264
rect 130804 85252 130810 85264
rect 189810 85252 189816 85264
rect 130804 85224 189816 85252
rect 130804 85212 130810 85224
rect 189810 85212 189816 85224
rect 189868 85212 189874 85264
rect 122282 85144 122288 85196
rect 122340 85184 122346 85196
rect 173250 85184 173256 85196
rect 122340 85156 173256 85184
rect 122340 85144 122346 85156
rect 173250 85144 173256 85156
rect 173308 85144 173314 85196
rect 75822 84124 75828 84176
rect 75880 84164 75886 84176
rect 216674 84164 216680 84176
rect 75880 84136 216680 84164
rect 75880 84124 75886 84136
rect 216674 84124 216680 84136
rect 216732 84124 216738 84176
rect 103330 84056 103336 84108
rect 103388 84096 103394 84108
rect 188522 84096 188528 84108
rect 103388 84068 188528 84096
rect 103388 84056 103394 84068
rect 188522 84056 188528 84068
rect 188580 84056 188586 84108
rect 117222 83988 117228 84040
rect 117280 84028 117286 84040
rect 178770 84028 178776 84040
rect 117280 84000 178776 84028
rect 117280 83988 117286 84000
rect 178770 83988 178776 84000
rect 178828 83988 178834 84040
rect 126790 83920 126796 83972
rect 126848 83960 126854 83972
rect 180334 83960 180340 83972
rect 126848 83932 180340 83960
rect 126848 83920 126854 83932
rect 180334 83920 180340 83932
rect 180392 83920 180398 83972
rect 180150 83444 180156 83496
rect 180208 83484 180214 83496
rect 265894 83484 265900 83496
rect 180208 83456 265900 83484
rect 180208 83444 180214 83456
rect 265894 83444 265900 83456
rect 265952 83444 265958 83496
rect 110230 82764 110236 82816
rect 110288 82804 110294 82816
rect 210418 82804 210424 82816
rect 110288 82776 210424 82804
rect 110288 82764 110294 82776
rect 210418 82764 210424 82776
rect 210476 82764 210482 82816
rect 114462 82696 114468 82748
rect 114520 82736 114526 82748
rect 213362 82736 213368 82748
rect 114520 82708 213368 82736
rect 114520 82696 114526 82708
rect 213362 82696 213368 82708
rect 213420 82696 213426 82748
rect 97902 82628 97908 82680
rect 97960 82668 97966 82680
rect 169110 82668 169116 82680
rect 97960 82640 169116 82668
rect 97960 82628 97966 82640
rect 169110 82628 169116 82640
rect 169168 82628 169174 82680
rect 103422 82560 103428 82612
rect 103480 82600 103486 82612
rect 174538 82600 174544 82612
rect 103480 82572 174544 82600
rect 103480 82560 103486 82572
rect 174538 82560 174544 82572
rect 174596 82560 174602 82612
rect 125502 82492 125508 82544
rect 125560 82532 125566 82544
rect 169018 82532 169024 82544
rect 125560 82504 169024 82532
rect 125560 82492 125566 82504
rect 169018 82492 169024 82504
rect 169076 82492 169082 82544
rect 111702 81336 111708 81388
rect 111760 81376 111766 81388
rect 207658 81376 207664 81388
rect 111760 81348 207664 81376
rect 111760 81336 111766 81348
rect 207658 81336 207664 81348
rect 207716 81336 207722 81388
rect 93762 81268 93768 81320
rect 93820 81308 93826 81320
rect 170398 81308 170404 81320
rect 93820 81280 170404 81308
rect 93820 81268 93826 81280
rect 170398 81268 170404 81280
rect 170456 81268 170462 81320
rect 104802 81200 104808 81252
rect 104860 81240 104866 81252
rect 175918 81240 175924 81252
rect 104860 81212 175924 81240
rect 104860 81200 104866 81212
rect 175918 81200 175924 81212
rect 175976 81200 175982 81252
rect 100570 81132 100576 81184
rect 100628 81172 100634 81184
rect 166350 81172 166356 81184
rect 100628 81144 166356 81172
rect 100628 81132 100634 81144
rect 166350 81132 166356 81144
rect 166408 81132 166414 81184
rect 126698 81064 126704 81116
rect 126756 81104 126762 81116
rect 184290 81104 184296 81116
rect 126756 81076 184296 81104
rect 126756 81064 126762 81076
rect 184290 81064 184296 81076
rect 184348 81064 184354 81116
rect 180058 80656 180064 80708
rect 180116 80696 180122 80708
rect 287054 80696 287060 80708
rect 180116 80668 287060 80696
rect 180116 80656 180122 80668
rect 287054 80656 287060 80668
rect 287112 80656 287118 80708
rect 115750 79976 115756 80028
rect 115808 80016 115814 80028
rect 209222 80016 209228 80028
rect 115808 79988 209228 80016
rect 115808 79976 115814 79988
rect 209222 79976 209228 79988
rect 209280 79976 209286 80028
rect 86862 79908 86868 79960
rect 86920 79948 86926 79960
rect 166442 79948 166448 79960
rect 86920 79920 166448 79948
rect 86920 79908 86926 79920
rect 166442 79908 166448 79920
rect 166500 79908 166506 79960
rect 95142 79840 95148 79892
rect 95200 79880 95206 79892
rect 174722 79880 174728 79892
rect 95200 79852 174728 79880
rect 95200 79840 95206 79852
rect 174722 79840 174728 79852
rect 174780 79840 174786 79892
rect 99190 79772 99196 79824
rect 99248 79812 99254 79824
rect 171962 79812 171968 79824
rect 99248 79784 171968 79812
rect 99248 79772 99254 79784
rect 171962 79772 171968 79784
rect 172020 79772 172026 79824
rect 113082 79704 113088 79756
rect 113140 79744 113146 79756
rect 185670 79744 185676 79756
rect 113140 79716 185676 79744
rect 113140 79704 113146 79716
rect 185670 79704 185676 79716
rect 185728 79704 185734 79756
rect 96522 78616 96528 78668
rect 96580 78656 96586 78668
rect 188430 78656 188436 78668
rect 96580 78628 188436 78656
rect 96580 78616 96586 78628
rect 188430 78616 188436 78628
rect 188488 78616 188494 78668
rect 128262 78548 128268 78600
rect 128320 78588 128326 78600
rect 213270 78588 213276 78600
rect 128320 78560 213276 78588
rect 128320 78548 128326 78560
rect 213270 78548 213276 78560
rect 213328 78548 213334 78600
rect 123478 78480 123484 78532
rect 123536 78520 123542 78532
rect 191282 78520 191288 78532
rect 123536 78492 191288 78520
rect 123536 78480 123542 78492
rect 191282 78480 191288 78492
rect 191340 78480 191346 78532
rect 110322 78412 110328 78464
rect 110380 78452 110386 78464
rect 173158 78452 173164 78464
rect 110380 78424 173164 78452
rect 110380 78412 110386 78424
rect 173158 78412 173164 78424
rect 173216 78412 173222 78464
rect 133138 77188 133144 77240
rect 133196 77228 133202 77240
rect 200850 77228 200856 77240
rect 133196 77200 200856 77228
rect 133196 77188 133202 77200
rect 200850 77188 200856 77200
rect 200908 77188 200914 77240
rect 118694 76576 118700 76628
rect 118752 76616 118758 76628
rect 256234 76616 256240 76628
rect 118752 76588 256240 76616
rect 118752 76576 118758 76588
rect 256234 76576 256240 76588
rect 256292 76576 256298 76628
rect 4154 76508 4160 76560
rect 4212 76548 4218 76560
rect 228358 76548 228364 76560
rect 4212 76520 228364 76548
rect 4212 76508 4218 76520
rect 228358 76508 228364 76520
rect 228416 76508 228422 76560
rect 106918 75828 106924 75880
rect 106976 75868 106982 75880
rect 192478 75868 192484 75880
rect 106976 75840 192484 75868
rect 106976 75828 106982 75840
rect 192478 75828 192484 75840
rect 192536 75828 192542 75880
rect 99098 75760 99104 75812
rect 99156 75800 99162 75812
rect 178862 75800 178868 75812
rect 99156 75772 178868 75800
rect 99156 75760 99162 75772
rect 178862 75760 178868 75772
rect 178920 75760 178926 75812
rect 67634 75216 67640 75268
rect 67692 75256 67698 75268
rect 263042 75256 263048 75268
rect 67692 75228 263048 75256
rect 67692 75216 67698 75228
rect 263042 75216 263048 75228
rect 263100 75216 263106 75268
rect 64690 75148 64696 75200
rect 64748 75188 64754 75200
rect 281534 75188 281540 75200
rect 64748 75160 281540 75188
rect 64748 75148 64754 75160
rect 281534 75148 281540 75160
rect 281592 75148 281598 75200
rect 124214 73856 124220 73908
rect 124272 73896 124278 73908
rect 230014 73896 230020 73908
rect 124272 73868 230020 73896
rect 124272 73856 124278 73868
rect 230014 73856 230020 73868
rect 230072 73856 230078 73908
rect 64598 73788 64604 73840
rect 64656 73828 64662 73840
rect 269114 73828 269120 73840
rect 64656 73800 269120 73828
rect 64656 73788 64662 73800
rect 269114 73788 269120 73800
rect 269172 73788 269178 73840
rect 80054 72428 80060 72480
rect 80112 72468 80118 72480
rect 242434 72468 242440 72480
rect 80112 72440 242440 72468
rect 80112 72428 80118 72440
rect 242434 72428 242440 72440
rect 242492 72428 242498 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 47578 71720 47584 71732
rect 3476 71692 47584 71720
rect 3476 71680 3482 71692
rect 47578 71680 47584 71692
rect 47636 71680 47642 71732
rect 74534 71068 74540 71120
rect 74592 71108 74598 71120
rect 261662 71108 261668 71120
rect 74592 71080 261668 71108
rect 74592 71068 74598 71080
rect 261662 71068 261668 71080
rect 261720 71068 261726 71120
rect 64414 71000 64420 71052
rect 64472 71040 64478 71052
rect 273254 71040 273260 71052
rect 64472 71012 273260 71040
rect 64472 71000 64478 71012
rect 273254 71000 273260 71012
rect 273312 71000 273318 71052
rect 77294 69640 77300 69692
rect 77352 69680 77358 69692
rect 254670 69680 254676 69692
rect 77352 69652 254676 69680
rect 77352 69640 77358 69652
rect 254670 69640 254676 69652
rect 254728 69640 254734 69692
rect 81434 68348 81440 68400
rect 81492 68388 81498 68400
rect 262950 68388 262956 68400
rect 81492 68360 262956 68388
rect 81492 68348 81498 68360
rect 262950 68348 262956 68360
rect 263008 68348 263014 68400
rect 46934 68280 46940 68332
rect 46992 68320 46998 68332
rect 236914 68320 236920 68332
rect 46992 68292 236920 68320
rect 46992 68280 46998 68292
rect 236914 68280 236920 68292
rect 236972 68280 236978 68332
rect 85574 66920 85580 66972
rect 85632 66960 85638 66972
rect 260190 66960 260196 66972
rect 85632 66932 260196 66960
rect 85632 66920 85638 66932
rect 260190 66920 260196 66932
rect 260248 66920 260254 66972
rect 53834 66852 53840 66904
rect 53892 66892 53898 66904
rect 247862 66892 247868 66904
rect 53892 66864 247868 66892
rect 53892 66852 53898 66864
rect 247862 66852 247868 66864
rect 247920 66852 247926 66904
rect 88334 65560 88340 65612
rect 88392 65600 88398 65612
rect 243538 65600 243544 65612
rect 88392 65572 243544 65600
rect 88392 65560 88398 65572
rect 243538 65560 243544 65572
rect 243596 65560 243602 65612
rect 64874 65492 64880 65544
rect 64932 65532 64938 65544
rect 253474 65532 253480 65544
rect 64932 65504 253480 65532
rect 64932 65492 64938 65504
rect 253474 65492 253480 65504
rect 253532 65492 253538 65544
rect 69014 64132 69020 64184
rect 69072 64172 69078 64184
rect 263134 64172 263140 64184
rect 69072 64144 263140 64172
rect 69072 64132 69078 64144
rect 263134 64132 263140 64144
rect 263192 64132 263198 64184
rect 75914 62772 75920 62824
rect 75972 62812 75978 62824
rect 249242 62812 249248 62824
rect 75972 62784 249248 62812
rect 75972 62772 75978 62784
rect 249242 62772 249248 62784
rect 249300 62772 249306 62824
rect 60734 61412 60740 61464
rect 60792 61452 60798 61464
rect 246482 61452 246488 61464
rect 60792 61424 246488 61452
rect 60792 61412 60798 61424
rect 246482 61412 246488 61424
rect 246540 61412 246546 61464
rect 78674 61344 78680 61396
rect 78732 61384 78738 61396
rect 264514 61384 264520 61396
rect 78732 61356 264520 61384
rect 78732 61344 78738 61356
rect 264514 61344 264520 61356
rect 264572 61344 264578 61396
rect 358078 60664 358084 60716
rect 358136 60704 358142 60716
rect 580166 60704 580172 60716
rect 358136 60676 580172 60704
rect 358136 60664 358142 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 82814 60052 82820 60104
rect 82872 60092 82878 60104
rect 238294 60092 238300 60104
rect 82872 60064 238300 60092
rect 82872 60052 82878 60064
rect 238294 60052 238300 60064
rect 238352 60052 238358 60104
rect 49694 59984 49700 60036
rect 49752 60024 49758 60036
rect 257430 60024 257436 60036
rect 49752 59996 257436 60024
rect 49752 59984 49758 59996
rect 257430 59984 257436 59996
rect 257488 59984 257494 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 53098 59344 53104 59356
rect 3108 59316 53104 59344
rect 3108 59304 3114 59316
rect 53098 59304 53104 59316
rect 53156 59304 53162 59356
rect 85666 58692 85672 58744
rect 85724 58732 85730 58744
rect 245102 58732 245108 58744
rect 85724 58704 245108 58732
rect 85724 58692 85730 58704
rect 245102 58692 245108 58704
rect 245160 58692 245166 58744
rect 52454 58624 52460 58676
rect 52512 58664 52518 58676
rect 265710 58664 265716 58676
rect 52512 58636 265716 58664
rect 52512 58624 52518 58636
rect 265710 58624 265716 58636
rect 265768 58624 265774 58676
rect 89714 57264 89720 57316
rect 89772 57304 89778 57316
rect 261754 57304 261760 57316
rect 89772 57276 261760 57304
rect 89772 57264 89778 57276
rect 261754 57264 261760 57276
rect 261812 57264 261818 57316
rect 9674 57196 9680 57248
rect 9732 57236 9738 57248
rect 253290 57236 253296 57248
rect 9732 57208 253296 57236
rect 9732 57196 9738 57208
rect 253290 57196 253296 57208
rect 253348 57196 253354 57248
rect 96614 55904 96620 55956
rect 96672 55944 96678 55956
rect 257614 55944 257620 55956
rect 96672 55916 257620 55944
rect 96672 55904 96678 55916
rect 257614 55904 257620 55916
rect 257672 55904 257678 55956
rect 41414 55836 41420 55888
rect 41472 55876 41478 55888
rect 234062 55876 234068 55888
rect 41472 55848 234068 55876
rect 41472 55836 41478 55848
rect 234062 55836 234068 55848
rect 234120 55836 234126 55888
rect 100754 54544 100760 54596
rect 100812 54584 100818 54596
rect 260374 54584 260380 54596
rect 100812 54556 260380 54584
rect 100812 54544 100818 54556
rect 260374 54544 260380 54556
rect 260432 54544 260438 54596
rect 34514 54476 34520 54528
rect 34572 54516 34578 54528
rect 243630 54516 243636 54528
rect 34572 54488 243636 54516
rect 34572 54476 34578 54488
rect 243630 54476 243636 54488
rect 243688 54476 243694 54528
rect 103514 53116 103520 53168
rect 103572 53156 103578 53168
rect 243722 53156 243728 53168
rect 103572 53128 243728 53156
rect 103572 53116 103578 53128
rect 243722 53116 243728 53128
rect 243780 53116 243786 53168
rect 30374 53048 30380 53100
rect 30432 53088 30438 53100
rect 260282 53088 260288 53100
rect 30432 53060 260288 53088
rect 30432 53048 30438 53060
rect 260282 53048 260288 53060
rect 260340 53048 260346 53100
rect 107654 51688 107660 51740
rect 107712 51728 107718 51740
rect 238202 51728 238208 51740
rect 107712 51700 238208 51728
rect 107712 51688 107718 51700
rect 238202 51688 238208 51700
rect 238260 51688 238266 51740
rect 106274 50396 106280 50448
rect 106332 50436 106338 50448
rect 229922 50436 229928 50448
rect 106332 50408 229928 50436
rect 106332 50396 106338 50408
rect 229922 50396 229928 50408
rect 229980 50396 229986 50448
rect 16574 50328 16580 50380
rect 16632 50368 16638 50380
rect 246574 50368 246580 50380
rect 16632 50340 246580 50368
rect 16632 50328 16638 50340
rect 246574 50328 246580 50340
rect 246632 50328 246638 50380
rect 118786 49036 118792 49088
rect 118844 49076 118850 49088
rect 253382 49076 253388 49088
rect 118844 49048 253388 49076
rect 118844 49036 118850 49048
rect 253382 49036 253388 49048
rect 253440 49036 253446 49088
rect 17954 48968 17960 49020
rect 18012 49008 18018 49020
rect 242342 49008 242348 49020
rect 18012 48980 242348 49008
rect 18012 48968 18018 48980
rect 242342 48968 242348 48980
rect 242400 48968 242406 49020
rect 110414 47608 110420 47660
rect 110472 47648 110478 47660
rect 256142 47648 256148 47660
rect 110472 47620 256148 47648
rect 110472 47608 110478 47620
rect 256142 47608 256148 47620
rect 256200 47608 256206 47660
rect 22094 47540 22100 47592
rect 22152 47580 22158 47592
rect 250622 47580 250628 47592
rect 22152 47552 250628 47580
rect 22152 47540 22158 47552
rect 250622 47540 250628 47552
rect 250680 47540 250686 47592
rect 177390 46860 177396 46912
rect 177448 46900 177454 46912
rect 580166 46900 580172 46912
rect 177448 46872 580172 46900
rect 177448 46860 177454 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 122834 46248 122840 46300
rect 122892 46288 122898 46300
rect 238110 46288 238116 46300
rect 122892 46260 238116 46288
rect 122892 46248 122898 46260
rect 238110 46248 238116 46260
rect 238168 46248 238174 46300
rect 86954 46180 86960 46232
rect 87012 46220 87018 46232
rect 258902 46220 258908 46232
rect 87012 46192 258908 46220
rect 87012 46180 87018 46192
rect 258902 46180 258908 46192
rect 258960 46180 258966 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 40678 45540 40684 45552
rect 3476 45512 40684 45540
rect 3476 45500 3482 45512
rect 40678 45500 40684 45512
rect 40736 45500 40742 45552
rect 113174 44888 113180 44940
rect 113232 44928 113238 44940
rect 240870 44928 240876 44940
rect 113232 44900 240876 44928
rect 113232 44888 113238 44900
rect 240870 44888 240876 44900
rect 240928 44888 240934 44940
rect 48314 44820 48320 44872
rect 48372 44860 48378 44872
rect 258994 44860 259000 44872
rect 48372 44832 259000 44860
rect 48372 44820 48378 44832
rect 258994 44820 259000 44832
rect 259052 44820 259058 44872
rect 20714 43392 20720 43444
rect 20772 43432 20778 43444
rect 254762 43432 254768 43444
rect 20772 43404 254768 43432
rect 20772 43392 20778 43404
rect 254762 43392 254768 43404
rect 254820 43392 254826 43444
rect 35894 42100 35900 42152
rect 35952 42140 35958 42152
rect 235350 42140 235356 42152
rect 35952 42112 235356 42140
rect 35952 42100 35958 42112
rect 235350 42100 235356 42112
rect 235408 42100 235414 42152
rect 26234 42032 26240 42084
rect 26292 42072 26298 42084
rect 250714 42072 250720 42084
rect 26292 42044 250720 42072
rect 26292 42032 26298 42044
rect 250714 42032 250720 42044
rect 250772 42032 250778 42084
rect 28994 40672 29000 40724
rect 29052 40712 29058 40724
rect 252002 40712 252008 40724
rect 29052 40684 252008 40712
rect 29052 40672 29058 40684
rect 252002 40672 252008 40684
rect 252060 40672 252066 40724
rect 45554 39380 45560 39432
rect 45612 39420 45618 39432
rect 239490 39420 239496 39432
rect 45612 39392 239496 39420
rect 45612 39380 45618 39392
rect 239490 39380 239496 39392
rect 239548 39380 239554 39432
rect 35986 39312 35992 39364
rect 36044 39352 36050 39364
rect 257522 39352 257528 39364
rect 36044 39324 257528 39352
rect 36044 39312 36050 39324
rect 257522 39312 257528 39324
rect 257580 39312 257586 39364
rect 40034 37952 40040 38004
rect 40092 37992 40098 38004
rect 261570 37992 261576 38004
rect 40092 37964 261576 37992
rect 40092 37952 40098 37964
rect 261570 37952 261576 37964
rect 261628 37952 261634 38004
rect 31754 37884 31760 37936
rect 31812 37924 31818 37936
rect 256050 37924 256056 37936
rect 31812 37896 256056 37924
rect 31812 37884 31818 37896
rect 256050 37884 256056 37896
rect 256108 37884 256114 37936
rect 2774 36592 2780 36644
rect 2832 36632 2838 36644
rect 236822 36632 236828 36644
rect 2832 36604 236828 36632
rect 2832 36592 2838 36604
rect 236822 36592 236828 36604
rect 236880 36592 236886 36644
rect 37182 36524 37188 36576
rect 37240 36564 37246 36576
rect 280154 36564 280160 36576
rect 37240 36536 280160 36564
rect 37240 36524 37246 36536
rect 280154 36524 280160 36536
rect 280212 36524 280218 36576
rect 44174 35232 44180 35284
rect 44232 35272 44238 35284
rect 232590 35272 232596 35284
rect 44232 35244 232596 35272
rect 44232 35232 44238 35244
rect 232590 35232 232596 35244
rect 232648 35232 232654 35284
rect 27706 35164 27712 35216
rect 27764 35204 27770 35216
rect 247770 35204 247776 35216
rect 27764 35176 247776 35204
rect 27764 35164 27770 35176
rect 247770 35164 247776 35176
rect 247828 35164 247834 35216
rect 93854 33804 93860 33856
rect 93912 33844 93918 33856
rect 250530 33844 250536 33856
rect 93912 33816 250536 33844
rect 93912 33804 93918 33816
rect 250530 33804 250536 33816
rect 250588 33804 250594 33856
rect 44266 33736 44272 33788
rect 44324 33776 44330 33788
rect 245010 33776 245016 33788
rect 44324 33748 245016 33776
rect 44324 33736 44330 33748
rect 245010 33736 245016 33748
rect 245068 33736 245074 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 51718 33096 51724 33108
rect 3568 33068 51724 33096
rect 3568 33056 3574 33068
rect 51718 33056 51724 33068
rect 51776 33056 51782 33108
rect 187050 33056 187056 33108
rect 187108 33096 187114 33108
rect 580166 33096 580172 33108
rect 187108 33068 580172 33096
rect 187108 33056 187114 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 109034 32444 109040 32496
rect 109092 32484 109098 32496
rect 261478 32484 261484 32496
rect 109092 32456 261484 32484
rect 109092 32444 109098 32456
rect 261478 32444 261484 32456
rect 261536 32444 261542 32496
rect 51074 32376 51080 32428
rect 51132 32416 51138 32428
rect 233970 32416 233976 32428
rect 51132 32388 233976 32416
rect 51132 32376 51138 32388
rect 233970 32376 233976 32388
rect 234028 32376 234034 32428
rect 114554 31016 114560 31068
rect 114612 31056 114618 31068
rect 264422 31056 264428 31068
rect 114612 31028 264428 31056
rect 114612 31016 114618 31028
rect 264422 31016 264428 31028
rect 264480 31016 264486 31068
rect 71774 29656 71780 29708
rect 71832 29696 71838 29708
rect 240962 29696 240968 29708
rect 71832 29668 240968 29696
rect 71832 29656 71838 29668
rect 240962 29656 240968 29668
rect 241020 29656 241026 29708
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 249150 29628 249156 29640
rect 19392 29600 249156 29628
rect 19392 29588 19398 29600
rect 249150 29588 249156 29600
rect 249208 29588 249214 29640
rect 57974 28296 57980 28348
rect 58032 28336 58038 28348
rect 258810 28336 258816 28348
rect 58032 28308 258816 28336
rect 58032 28296 58038 28308
rect 258810 28296 258816 28308
rect 258868 28296 258874 28348
rect 23474 28228 23480 28280
rect 23532 28268 23538 28280
rect 250438 28268 250444 28280
rect 23532 28240 250444 28268
rect 23532 28228 23538 28240
rect 250438 28228 250444 28240
rect 250496 28228 250502 28280
rect 110506 26936 110512 26988
rect 110564 26976 110570 26988
rect 251910 26976 251916 26988
rect 110564 26948 251916 26976
rect 110564 26936 110570 26948
rect 251910 26936 251916 26948
rect 251968 26936 251974 26988
rect 6914 26868 6920 26920
rect 6972 26908 6978 26920
rect 242250 26908 242256 26920
rect 6972 26880 242256 26908
rect 6972 26868 6978 26880
rect 242250 26868 242256 26880
rect 242308 26868 242314 26920
rect 120074 25508 120080 25560
rect 120132 25548 120138 25560
rect 236730 25548 236736 25560
rect 120132 25520 236736 25548
rect 120132 25508 120138 25520
rect 236730 25508 236736 25520
rect 236788 25508 236794 25560
rect 102134 22856 102140 22908
rect 102192 22896 102198 22908
rect 236638 22896 236644 22908
rect 102192 22868 236644 22896
rect 102192 22856 102198 22868
rect 236638 22856 236644 22868
rect 236696 22856 236702 22908
rect 63402 22788 63408 22840
rect 63460 22828 63466 22840
rect 284386 22828 284392 22840
rect 63460 22800 284392 22828
rect 63460 22788 63466 22800
rect 284386 22788 284392 22800
rect 284444 22788 284450 22840
rect 14 22720 20 22772
rect 72 22760 78 22772
rect 230474 22760 230480 22772
rect 72 22732 230480 22760
rect 72 22720 78 22732
rect 230474 22720 230480 22732
rect 230532 22720 230538 22772
rect 52546 21428 52552 21480
rect 52604 21468 52610 21480
rect 246390 21468 246396 21480
rect 52604 21440 246396 21468
rect 52604 21428 52610 21440
rect 246390 21428 246396 21440
rect 246448 21428 246454 21480
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 253198 21400 253204 21412
rect 11112 21372 253204 21400
rect 11112 21360 11118 21372
rect 253198 21360 253204 21372
rect 253256 21360 253262 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 29638 20652 29644 20664
rect 3476 20624 29644 20652
rect 3476 20612 3482 20624
rect 29638 20612 29644 20624
rect 29696 20612 29702 20664
rect 195330 20000 195336 20052
rect 195388 20040 195394 20052
rect 271874 20040 271880 20052
rect 195388 20012 271880 20040
rect 195388 20000 195394 20012
rect 271874 20000 271880 20012
rect 271932 20000 271938 20052
rect 97994 19932 98000 19984
rect 98052 19972 98058 19984
rect 260098 19972 260104 19984
rect 98052 19944 260104 19972
rect 98052 19932 98058 19944
rect 260098 19932 260104 19944
rect 260156 19932 260162 19984
rect 206370 18708 206376 18760
rect 206428 18748 206434 18760
rect 285674 18748 285680 18760
rect 206428 18720 285680 18748
rect 206428 18708 206434 18720
rect 285674 18708 285680 18720
rect 285732 18708 285738 18760
rect 104894 18640 104900 18692
rect 104952 18680 104958 18692
rect 222838 18680 222844 18692
rect 104952 18652 222844 18680
rect 104952 18640 104958 18652
rect 222838 18640 222844 18652
rect 222896 18640 222902 18692
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 239398 18612 239404 18624
rect 8352 18584 239404 18612
rect 8352 18572 8358 18584
rect 239398 18572 239404 18584
rect 239456 18572 239462 18624
rect 196618 17348 196624 17400
rect 196676 17388 196682 17400
rect 241514 17388 241520 17400
rect 196676 17360 241520 17388
rect 196676 17348 196682 17360
rect 241514 17348 241520 17360
rect 241572 17348 241578 17400
rect 77386 17280 77392 17332
rect 77444 17320 77450 17332
rect 249058 17320 249064 17332
rect 77444 17292 249064 17320
rect 77444 17280 77450 17292
rect 249058 17280 249064 17292
rect 249116 17280 249122 17332
rect 55214 17212 55220 17264
rect 55272 17252 55278 17264
rect 255958 17252 255964 17264
rect 55272 17224 255964 17252
rect 55272 17212 55278 17224
rect 255958 17212 255964 17224
rect 256016 17212 256022 17264
rect 204898 15988 204904 16040
rect 204956 16028 204962 16040
rect 276106 16028 276112 16040
rect 204956 16000 276112 16028
rect 204956 15988 204962 16000
rect 276106 15988 276112 16000
rect 276164 15988 276170 16040
rect 122282 15920 122288 15972
rect 122340 15960 122346 15972
rect 258718 15960 258724 15972
rect 122340 15932 258724 15960
rect 122340 15920 122346 15932
rect 258718 15920 258724 15932
rect 258776 15920 258782 15972
rect 69842 15852 69848 15904
rect 69900 15892 69906 15904
rect 247678 15892 247684 15904
rect 69900 15864 247684 15892
rect 69900 15852 69906 15864
rect 247678 15852 247684 15864
rect 247736 15852 247742 15904
rect 202138 14560 202144 14612
rect 202196 14600 202202 14612
rect 268378 14600 268384 14612
rect 202196 14572 268384 14600
rect 202196 14560 202202 14572
rect 268378 14560 268384 14572
rect 268436 14560 268442 14612
rect 102226 14492 102232 14544
rect 102284 14532 102290 14544
rect 232498 14532 232504 14544
rect 102284 14504 232504 14532
rect 102284 14492 102290 14504
rect 232498 14492 232504 14504
rect 232556 14492 232562 14544
rect 33594 14424 33600 14476
rect 33652 14464 33658 14476
rect 264330 14464 264336 14476
rect 33652 14436 264336 14464
rect 33652 14424 33658 14436
rect 264330 14424 264336 14436
rect 264388 14424 264394 14476
rect 197998 13200 198004 13252
rect 198056 13240 198062 13252
rect 261754 13240 261760 13252
rect 198056 13212 261760 13240
rect 198056 13200 198062 13212
rect 261754 13200 261760 13212
rect 261812 13200 261818 13252
rect 63218 13132 63224 13184
rect 63276 13172 63282 13184
rect 246298 13172 246304 13184
rect 63276 13144 246304 13172
rect 63276 13132 63282 13144
rect 246298 13132 246304 13144
rect 246356 13132 246362 13184
rect 13538 13064 13544 13116
rect 13596 13104 13602 13116
rect 229830 13104 229836 13116
rect 13596 13076 229836 13104
rect 13596 13064 13602 13076
rect 229830 13064 229836 13076
rect 229888 13064 229894 13116
rect 199470 11772 199476 11824
rect 199528 11812 199534 11824
rect 292574 11812 292580 11824
rect 199528 11784 292580 11812
rect 199528 11772 199534 11784
rect 292574 11772 292580 11784
rect 292632 11772 292638 11824
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 265618 11744 265624 11756
rect 15988 11716 265624 11744
rect 15988 11704 15994 11716
rect 265618 11704 265624 11716
rect 265676 11704 265682 11756
rect 91554 10344 91560 10396
rect 91612 10384 91618 10396
rect 257338 10384 257344 10396
rect 91612 10356 257344 10384
rect 91612 10344 91618 10356
rect 257338 10344 257344 10356
rect 257396 10344 257402 10396
rect 25314 10276 25320 10328
rect 25372 10316 25378 10328
rect 238018 10316 238024 10328
rect 25372 10288 238024 10316
rect 25372 10276 25378 10288
rect 238018 10276 238024 10288
rect 238076 10276 238082 10328
rect 198090 9120 198096 9172
rect 198148 9160 198154 9172
rect 262950 9160 262956 9172
rect 198148 9132 262956 9160
rect 198148 9120 198154 9132
rect 262950 9120 262956 9132
rect 263008 9120 263014 9172
rect 39666 9052 39672 9104
rect 39724 9092 39730 9104
rect 132954 9092 132960 9104
rect 39724 9064 132960 9092
rect 39724 9052 39730 9064
rect 132954 9052 132960 9064
rect 133012 9052 133018 9104
rect 203518 9052 203524 9104
rect 203576 9092 203582 9104
rect 271230 9092 271236 9104
rect 203576 9064 271236 9092
rect 203576 9052 203582 9064
rect 271230 9052 271236 9064
rect 271288 9052 271294 9104
rect 95142 8984 95148 9036
rect 95200 9024 95206 9036
rect 262858 9024 262864 9036
rect 95200 8996 262864 9024
rect 95200 8984 95206 8996
rect 262858 8984 262864 8996
rect 262916 8984 262922 9036
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 231118 8956 231124 8968
rect 11204 8928 231124 8956
rect 11204 8916 11210 8928
rect 231118 8916 231124 8928
rect 231176 8916 231182 8968
rect 34422 7692 34428 7744
rect 34480 7732 34486 7744
rect 136450 7732 136456 7744
rect 34480 7704 136456 7732
rect 34480 7692 34486 7704
rect 136450 7692 136456 7704
rect 136508 7692 136514 7744
rect 191098 7692 191104 7744
rect 191156 7732 191162 7744
rect 239306 7732 239312 7744
rect 191156 7704 239312 7732
rect 191156 7692 191162 7704
rect 239306 7692 239312 7704
rect 239364 7692 239370 7744
rect 112806 7624 112812 7676
rect 112864 7664 112870 7676
rect 244918 7664 244924 7676
rect 112864 7636 244924 7664
rect 112864 7624 112870 7636
rect 244918 7624 244924 7636
rect 244976 7624 244982 7676
rect 66714 7556 66720 7608
rect 66772 7596 66778 7608
rect 264238 7596 264244 7608
rect 66772 7568 264244 7596
rect 66772 7556 66778 7568
rect 264238 7556 264244 7568
rect 264296 7556 264302 7608
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 4798 6644 4804 6656
rect 3016 6616 4804 6644
rect 3016 6604 3022 6616
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 204990 6332 204996 6384
rect 205048 6372 205054 6384
rect 260650 6372 260656 6384
rect 205048 6344 260656 6372
rect 205048 6332 205054 6344
rect 260650 6332 260656 6344
rect 260708 6332 260714 6384
rect 44082 6264 44088 6316
rect 44140 6304 44146 6316
rect 129366 6304 129372 6316
rect 44140 6276 129372 6304
rect 44140 6264 44146 6276
rect 129366 6264 129372 6276
rect 129424 6264 129430 6316
rect 206278 6264 206284 6316
rect 206336 6304 206342 6316
rect 283098 6304 283104 6316
rect 206336 6276 283104 6304
rect 206336 6264 206342 6276
rect 283098 6264 283104 6276
rect 283156 6264 283162 6316
rect 59630 6196 59636 6248
rect 59688 6236 59694 6248
rect 235258 6236 235264 6248
rect 59688 6208 235264 6236
rect 59688 6196 59694 6208
rect 235258 6196 235264 6208
rect 235316 6196 235322 6248
rect 73798 6128 73804 6180
rect 73856 6168 73862 6180
rect 254578 6168 254584 6180
rect 73856 6140 254584 6168
rect 73856 6128 73862 6140
rect 254578 6128 254584 6140
rect 254636 6128 254642 6180
rect 193858 4972 193864 5024
rect 193916 5012 193922 5024
rect 244090 5012 244096 5024
rect 193916 4984 244096 5012
rect 193916 4972 193922 4984
rect 244090 4972 244096 4984
rect 244148 4972 244154 5024
rect 213178 4904 213184 4956
rect 213236 4944 213242 4956
rect 264146 4944 264152 4956
rect 213236 4916 264152 4944
rect 213236 4904 213242 4916
rect 264146 4904 264152 4916
rect 264204 4904 264210 4956
rect 96246 4836 96252 4888
rect 96304 4876 96310 4888
rect 229738 4876 229744 4888
rect 96304 4848 229744 4876
rect 96304 4836 96310 4848
rect 229738 4836 229744 4848
rect 229796 4836 229802 4888
rect 62022 4768 62028 4820
rect 62080 4808 62086 4820
rect 242158 4808 242164 4820
rect 62080 4780 242164 4808
rect 62080 4768 62086 4780
rect 242158 4768 242164 4780
rect 242216 4768 242222 4820
rect 216030 3680 216036 3732
rect 216088 3720 216094 3732
rect 242894 3720 242900 3732
rect 216088 3692 242900 3720
rect 216088 3680 216094 3692
rect 242894 3680 242900 3692
rect 242952 3680 242958 3732
rect 209038 3612 209044 3664
rect 209096 3652 209102 3664
rect 247586 3652 247592 3664
rect 209096 3624 247592 3652
rect 209096 3612 209102 3624
rect 247586 3612 247592 3624
rect 247644 3612 247650 3664
rect 266998 3612 267004 3664
rect 267056 3652 267062 3664
rect 285398 3652 285404 3664
rect 267056 3624 285404 3652
rect 267056 3612 267062 3624
rect 285398 3612 285404 3624
rect 285456 3612 285462 3664
rect 332686 3612 332692 3664
rect 332744 3652 332750 3664
rect 333882 3652 333888 3664
rect 332744 3624 333888 3652
rect 332744 3612 332750 3624
rect 333882 3612 333888 3624
rect 333940 3612 333946 3664
rect 52454 3544 52460 3596
rect 52512 3584 52518 3596
rect 53374 3584 53380 3596
rect 52512 3556 53380 3584
rect 52512 3544 52518 3556
rect 53374 3544 53380 3556
rect 53432 3544 53438 3596
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 78214 3584 78220 3596
rect 77352 3556 78220 3584
rect 77352 3544 77358 3556
rect 78214 3544 78220 3556
rect 78272 3544 78278 3596
rect 99834 3544 99840 3596
rect 99892 3584 99898 3596
rect 99892 3556 103514 3584
rect 99892 3544 99898 3556
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 98638 3516 98644 3528
rect 6512 3488 98644 3516
rect 6512 3476 6518 3488
rect 98638 3476 98644 3488
rect 98696 3476 98702 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 103486 3516 103514 3556
rect 110414 3544 110420 3596
rect 110472 3584 110478 3596
rect 111610 3584 111616 3596
rect 110472 3556 111616 3584
rect 110472 3544 110478 3556
rect 111610 3544 111616 3556
rect 111668 3544 111674 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 173894 3584 173900 3596
rect 125928 3556 173900 3584
rect 125928 3544 125934 3556
rect 173894 3544 173900 3556
rect 173952 3544 173958 3596
rect 202230 3544 202236 3596
rect 202288 3584 202294 3596
rect 267734 3584 267740 3596
rect 202288 3556 267740 3584
rect 202288 3544 202294 3556
rect 267734 3544 267740 3556
rect 267792 3544 267798 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 276750 3584 276756 3596
rect 276072 3556 276756 3584
rect 276072 3544 276078 3556
rect 276750 3544 276756 3556
rect 276808 3544 276814 3596
rect 316126 3544 316132 3596
rect 316184 3584 316190 3596
rect 317322 3584 317328 3596
rect 316184 3556 317328 3584
rect 316184 3544 316190 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 335998 3544 336004 3596
rect 336056 3544 336062 3596
rect 196710 3516 196716 3528
rect 103486 3488 196716 3516
rect 196710 3476 196716 3488
rect 196768 3476 196774 3528
rect 215938 3476 215944 3528
rect 215996 3516 216002 3528
rect 290182 3516 290188 3528
rect 215996 3488 290188 3516
rect 215996 3476 216002 3488
rect 290182 3476 290188 3488
rect 290240 3476 290246 3528
rect 324406 3476 324412 3528
rect 324464 3516 324470 3528
rect 325602 3516 325608 3528
rect 324464 3488 325608 3516
rect 324464 3476 324470 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 331858 3476 331864 3528
rect 331916 3516 331922 3528
rect 332686 3516 332692 3528
rect 331916 3488 332692 3516
rect 331916 3476 331922 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 38378 3408 38384 3460
rect 38436 3448 38442 3460
rect 180150 3448 180156 3460
rect 38436 3420 180156 3448
rect 38436 3408 38442 3420
rect 180150 3408 180156 3420
rect 180208 3408 180214 3460
rect 195238 3408 195244 3460
rect 195296 3448 195302 3460
rect 274818 3448 274824 3460
rect 195296 3420 274824 3448
rect 195296 3408 195302 3420
rect 274818 3408 274824 3420
rect 274876 3408 274882 3460
rect 336016 3448 336044 3544
rect 340966 3476 340972 3528
rect 341024 3516 341030 3528
rect 342162 3516 342168 3528
rect 341024 3488 342168 3516
rect 341024 3476 341030 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 349246 3476 349252 3528
rect 349304 3516 349310 3528
rect 350442 3516 350448 3528
rect 349304 3488 350448 3516
rect 349304 3476 349310 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 336016 3420 349292 3448
rect 349264 3392 349292 3420
rect 233878 3340 233884 3392
rect 233936 3380 233942 3392
rect 235810 3380 235816 3392
rect 233936 3352 235816 3380
rect 233936 3340 233942 3352
rect 235810 3340 235816 3352
rect 235868 3340 235874 3392
rect 309870 3340 309876 3392
rect 309928 3380 309934 3392
rect 311434 3380 311440 3392
rect 309928 3352 311440 3380
rect 309928 3340 309934 3352
rect 311434 3340 311440 3352
rect 311492 3340 311498 3392
rect 349246 3340 349252 3392
rect 349304 3340 349310 3392
rect 322198 3000 322204 3052
rect 322256 3040 322262 3052
rect 324406 3040 324412 3052
rect 322256 3012 324412 3040
rect 322256 3000 322262 3012
rect 324406 3000 324412 3012
rect 324464 3000 324470 3052
rect 186958 2184 186964 2236
rect 187016 2224 187022 2236
rect 265342 2224 265348 2236
rect 187016 2196 265348 2224
rect 187016 2184 187022 2196
rect 265342 2184 265348 2196
rect 265400 2184 265406 2236
rect 116394 2116 116400 2168
rect 116452 2156 116458 2168
rect 251818 2156 251824 2168
rect 116452 2128 251824 2156
rect 116452 2116 116458 2128
rect 251818 2116 251824 2128
rect 251876 2116 251882 2168
rect 84470 2048 84476 2100
rect 84528 2088 84534 2100
rect 240778 2088 240784 2100
rect 84528 2060 240784 2088
rect 84528 2048 84534 2060
rect 240778 2048 240784 2060
rect 240836 2048 240842 2100
rect 307754 824 307760 876
rect 307812 864 307818 876
rect 309042 864 309048 876
rect 307812 836 309048 864
rect 307812 824 307818 836
rect 309042 824 309048 836
rect 309100 824 309106 876
<< via1 >>
rect 201500 703196 201552 703248
rect 202788 703196 202840 703248
rect 95148 703128 95200 703180
rect 332508 703128 332560 703180
rect 116584 703060 116636 703112
rect 397460 703060 397512 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 76564 702992 76616 703044
rect 364984 702992 365036 703044
rect 104808 702924 104860 702976
rect 413652 702924 413704 702976
rect 113088 702856 113140 702908
rect 462320 702856 462372 702908
rect 75184 702788 75236 702840
rect 429844 702788 429896 702840
rect 110328 702720 110380 702772
rect 478512 702720 478564 702772
rect 115848 702652 115900 702704
rect 494796 702652 494848 702704
rect 111708 702584 111760 702636
rect 559656 702584 559708 702636
rect 79324 702516 79376 702568
rect 527180 702516 527232 702568
rect 68928 702448 68980 702500
rect 543464 702448 543516 702500
rect 8116 700340 8168 700392
rect 85580 700340 85632 700392
rect 97264 700340 97316 700392
rect 154120 700340 154172 700392
rect 155224 700340 155276 700392
rect 218980 700340 219032 700392
rect 62028 700272 62080 700324
rect 235172 700272 235224 700324
rect 24308 698912 24360 698964
rect 106280 698912 106332 698964
rect 57888 697552 57940 697604
rect 170312 697552 170364 697604
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 69020 696940 69072 696992
rect 580172 696940 580224 696992
rect 122748 683136 122800 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 57980 670692 58032 670744
rect 83464 670692 83516 670744
rect 580172 670692 580224 670744
rect 3516 658112 3568 658164
rect 7564 658112 7616 658164
rect 129004 643084 129056 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 3516 618264 3568 618316
rect 87604 618264 87656 618316
rect 411904 616836 411956 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 35164 605820 35216 605872
rect 68836 596776 68888 596828
rect 136640 596776 136692 596828
rect 78036 595416 78088 595468
rect 266360 595416 266412 595468
rect 40040 591268 40092 591320
rect 55864 591268 55916 591320
rect 111616 590656 111668 590708
rect 580172 590656 580224 590708
rect 68468 589908 68520 589960
rect 97264 589908 97316 589960
rect 7564 588548 7616 588600
rect 87328 588548 87380 588600
rect 87604 587868 87656 587920
rect 95240 587868 95292 587920
rect 81716 587800 81768 587852
rect 83464 587800 83516 587852
rect 3424 587120 3476 587172
rect 53840 587120 53892 587172
rect 88340 587120 88392 587172
rect 111800 587120 111852 587172
rect 133236 587120 133288 587172
rect 155224 587120 155276 587172
rect 94136 586780 94188 586832
rect 117504 586780 117556 586832
rect 91560 586712 91612 586764
rect 123116 586712 123168 586764
rect 94872 586644 94924 586696
rect 127072 586644 127124 586696
rect 46848 586576 46900 586628
rect 85120 586576 85172 586628
rect 90272 586576 90324 586628
rect 124312 586576 124364 586628
rect 41236 586508 41288 586560
rect 80612 586508 80664 586560
rect 98736 586508 98788 586560
rect 133236 586508 133288 586560
rect 69112 585760 69164 585812
rect 282920 585760 282972 585812
rect 54484 585352 54536 585404
rect 76564 585352 76616 585404
rect 95240 585352 95292 585404
rect 95884 585352 95936 585404
rect 118700 585352 118752 585404
rect 52184 585284 52236 585336
rect 78036 585284 78088 585336
rect 95148 585284 95200 585336
rect 122840 585284 122892 585336
rect 34244 585216 34296 585268
rect 72240 585216 72292 585268
rect 92296 585216 92348 585268
rect 125600 585216 125652 585268
rect 46756 585148 46808 585200
rect 85580 585148 85632 585200
rect 87328 585148 87380 585200
rect 87512 585148 87564 585200
rect 121460 585148 121512 585200
rect 103152 584400 103204 584452
rect 104808 584400 104860 584452
rect 116308 584400 116360 584452
rect 37004 584060 37056 584112
rect 75460 584060 75512 584112
rect 77852 584060 77904 584112
rect 79324 584060 79376 584112
rect 59268 583992 59320 584044
rect 101312 583992 101364 584044
rect 113180 583992 113232 584044
rect 53564 583924 53616 583976
rect 75092 583924 75144 583976
rect 101864 583924 101916 583976
rect 114560 583924 114612 583976
rect 57704 583856 57756 583908
rect 81440 583856 81492 583908
rect 81716 583856 81768 583908
rect 88984 583856 89036 583908
rect 100760 583856 100812 583908
rect 105544 583856 105596 583908
rect 118792 583856 118844 583908
rect 61752 583788 61804 583840
rect 87696 583788 87748 583840
rect 96528 583788 96580 583840
rect 110696 583788 110748 583840
rect 69204 583720 69256 583772
rect 73344 583720 73396 583772
rect 97448 583720 97500 583772
rect 124220 583720 124272 583772
rect 60004 582972 60056 583024
rect 71872 582972 71924 583024
rect 100760 582972 100812 583024
rect 124496 582972 124548 583024
rect 11704 582700 11756 582752
rect 107660 582700 107712 582752
rect 55128 582632 55180 582684
rect 78680 582632 78732 582684
rect 56324 582564 56376 582616
rect 81900 582564 81952 582616
rect 89628 582564 89680 582616
rect 118976 582564 119028 582616
rect 52092 582496 52144 582548
rect 79324 582496 79376 582548
rect 99288 582496 99340 582548
rect 129740 582496 129792 582548
rect 103888 582428 103940 582480
rect 116124 582428 116176 582480
rect 68744 582360 68796 582412
rect 386328 582360 386380 582412
rect 70400 581680 70452 581732
rect 70952 581680 71004 581732
rect 43812 581272 43864 581324
rect 67640 581272 67692 581324
rect 59084 581204 59136 581256
rect 70400 581204 70452 581256
rect 57796 581136 57848 581188
rect 82728 581748 82780 581800
rect 104992 581748 105044 581800
rect 111984 581748 112036 581800
rect 76748 581680 76800 581732
rect 100576 581680 100628 581732
rect 50804 581068 50856 581120
rect 35624 581000 35676 581052
rect 70492 581000 70544 581052
rect 104440 581680 104492 581732
rect 123024 581068 123076 581120
rect 121552 581000 121604 581052
rect 39948 580252 40000 580304
rect 67916 580252 67968 580304
rect 3240 579708 3292 579760
rect 7564 579708 7616 579760
rect 108948 579640 109000 579692
rect 120172 579640 120224 579692
rect 106740 578892 106792 578944
rect 121644 578892 121696 578944
rect 59176 578280 59228 578332
rect 67640 578280 67692 578332
rect 108856 578280 108908 578332
rect 117320 578280 117372 578332
rect 108948 578212 109000 578264
rect 134064 578212 134116 578264
rect 108212 578144 108264 578196
rect 111708 578144 111760 578196
rect 386328 578144 386380 578196
rect 579804 578144 579856 578196
rect 63224 576852 63276 576904
rect 67640 576852 67692 576904
rect 108948 575560 109000 575612
rect 126244 575560 126296 575612
rect 34428 575492 34480 575544
rect 67640 575492 67692 575544
rect 108856 575492 108908 575544
rect 129832 575492 129884 575544
rect 64604 574132 64656 574184
rect 67732 574132 67784 574184
rect 53748 574064 53800 574116
rect 67640 574064 67692 574116
rect 108948 573996 109000 574048
rect 121920 573996 121972 574048
rect 121920 573316 121972 573368
rect 122748 573316 122800 573368
rect 131764 573316 131816 573368
rect 108948 572840 109000 572892
rect 113364 572840 113416 572892
rect 64696 572772 64748 572824
rect 67732 572772 67784 572824
rect 107844 572772 107896 572824
rect 110512 572772 110564 572824
rect 61844 572704 61896 572756
rect 67640 572704 67692 572756
rect 105636 572296 105688 572348
rect 109224 572296 109276 572348
rect 66168 571548 66220 571600
rect 68284 571548 68336 571600
rect 108948 571344 109000 571396
rect 128360 571344 128412 571396
rect 108856 569984 108908 570036
rect 132500 569984 132552 570036
rect 39304 569916 39356 569968
rect 67640 569916 67692 569968
rect 108948 569916 109000 569968
rect 135352 569916 135404 569968
rect 64788 568624 64840 568676
rect 67640 568624 67692 568676
rect 108948 568556 109000 568608
rect 120080 568556 120132 568608
rect 108948 567536 109000 567588
rect 114652 567536 114704 567588
rect 66076 567196 66128 567248
rect 67640 567196 67692 567248
rect 108948 567196 109000 567248
rect 115940 567196 115992 567248
rect 108856 565904 108908 565956
rect 117412 565904 117464 565956
rect 3424 565836 3476 565888
rect 22744 565836 22796 565888
rect 108948 565836 109000 565888
rect 125876 565836 125928 565888
rect 65984 564476 66036 564528
rect 67732 564476 67784 564528
rect 49608 564408 49660 564460
rect 67640 564408 67692 564460
rect 108948 564408 109000 564460
rect 131028 564408 131080 564460
rect 413284 564408 413336 564460
rect 108948 563728 109000 563780
rect 110328 563728 110380 563780
rect 136824 563728 136876 563780
rect 126244 563660 126296 563712
rect 580172 563660 580224 563712
rect 61936 563116 61988 563168
rect 67640 563116 67692 563168
rect 48136 563048 48188 563100
rect 67732 563048 67784 563100
rect 60740 562980 60792 563032
rect 62028 562980 62080 563032
rect 67640 562980 67692 563032
rect 52276 562300 52328 562352
rect 60740 562300 60792 562352
rect 107660 560328 107712 560380
rect 120264 560328 120316 560380
rect 50988 560260 51040 560312
rect 67640 560260 67692 560312
rect 108948 560260 109000 560312
rect 139492 560260 139544 560312
rect 128636 559512 128688 559564
rect 201500 559512 201552 559564
rect 108856 558968 108908 559020
rect 128636 558968 128688 559020
rect 45468 558900 45520 558952
rect 67640 558900 67692 558952
rect 108948 558900 109000 558952
rect 138112 558900 138164 558952
rect 108580 558016 108632 558068
rect 111892 558016 111944 558068
rect 62764 557540 62816 557592
rect 67640 557540 67692 557592
rect 108948 556520 109000 556572
rect 113272 556520 113324 556572
rect 53656 556248 53708 556300
rect 67732 556248 67784 556300
rect 43904 556180 43956 556232
rect 67640 556180 67692 556232
rect 57888 556112 57940 556164
rect 67732 556112 67784 556164
rect 48228 555432 48280 555484
rect 57888 555432 57940 555484
rect 35716 554752 35768 554804
rect 67640 554752 67692 554804
rect 109224 554752 109276 554804
rect 115204 554752 115256 554804
rect 3148 554684 3200 554736
rect 11704 554684 11756 554736
rect 108948 554004 109000 554056
rect 111616 554004 111668 554056
rect 133972 554004 134024 554056
rect 57244 553392 57296 553444
rect 67640 553392 67692 553444
rect 108948 553392 109000 553444
rect 127256 553392 127308 553444
rect 129004 553392 129056 553444
rect 50896 552032 50948 552084
rect 67640 552032 67692 552084
rect 108948 552032 109000 552084
rect 136640 552032 136692 552084
rect 42708 550604 42760 550656
rect 67640 550604 67692 550656
rect 108948 550604 109000 550656
rect 131120 550604 131172 550656
rect 63408 549312 63460 549364
rect 67640 549312 67692 549364
rect 108948 549312 109000 549364
rect 139400 549312 139452 549364
rect 44088 549244 44140 549296
rect 67732 549244 67784 549296
rect 108856 549244 108908 549296
rect 140964 549244 141016 549296
rect 67272 549108 67324 549160
rect 68376 549108 68428 549160
rect 107844 548360 107896 548412
rect 110604 548360 110656 548412
rect 107660 548224 107712 548276
rect 107844 548224 107896 548276
rect 41144 547884 41196 547936
rect 67640 547884 67692 547936
rect 133788 547136 133840 547188
rect 299480 547136 299532 547188
rect 63316 546524 63368 546576
rect 67732 546524 67784 546576
rect 109684 546524 109736 546576
rect 133144 546524 133196 546576
rect 133788 546524 133840 546576
rect 60648 546456 60700 546508
rect 67640 546456 67692 546508
rect 108948 546456 109000 546508
rect 142344 546456 142396 546508
rect 37188 545708 37240 545760
rect 68744 545708 68796 545760
rect 108948 545708 109000 545760
rect 115848 545708 115900 545760
rect 124404 545708 124456 545760
rect 108948 545096 109000 545148
rect 135444 545096 135496 545148
rect 22744 544348 22796 544400
rect 33140 544348 33192 544400
rect 108948 544348 109000 544400
rect 113088 544348 113140 544400
rect 136732 544348 136784 544400
rect 38568 543804 38620 543856
rect 67732 543804 67784 543856
rect 33140 543736 33192 543788
rect 34336 543736 34388 543788
rect 67640 543736 67692 543788
rect 60556 542444 60608 542496
rect 67640 542444 67692 542496
rect 49424 542376 49476 542428
rect 68928 542376 68980 542428
rect 108948 542376 109000 542428
rect 142160 542376 142212 542428
rect 109776 541628 109828 541680
rect 580264 541628 580316 541680
rect 62028 540948 62080 541000
rect 67640 540948 67692 541000
rect 108948 540948 109000 541000
rect 140780 540948 140832 541000
rect 41328 539656 41380 539708
rect 60004 539656 60056 539708
rect 37096 539588 37148 539640
rect 67640 539588 67692 539640
rect 4804 539520 4856 539572
rect 99012 539520 99064 539572
rect 57980 539452 58032 539504
rect 91284 539452 91336 539504
rect 99196 539044 99248 539096
rect 111984 539044 112036 539096
rect 99012 538976 99064 539028
rect 122932 538976 122984 539028
rect 95148 538908 95200 538960
rect 121644 538908 121696 538960
rect 61752 538840 61804 538892
rect 83004 538840 83056 538892
rect 88064 538840 88116 538892
rect 122104 538840 122156 538892
rect 411904 538840 411956 538892
rect 413284 538840 413336 538892
rect 580908 538840 580960 538892
rect 57520 538568 57572 538620
rect 57980 538568 58032 538620
rect 7564 538160 7616 538212
rect 98368 538160 98420 538212
rect 103520 538160 103572 538212
rect 109684 538160 109736 538212
rect 60004 538092 60056 538144
rect 73896 538092 73948 538144
rect 94504 538092 94556 538144
rect 104716 538092 104768 538144
rect 102232 537752 102284 537804
rect 127164 537752 127216 537804
rect 95792 537684 95844 537736
rect 121736 537684 121788 537736
rect 59084 537616 59136 537668
rect 69756 537616 69808 537668
rect 85488 537616 85540 537668
rect 98644 537616 98696 537668
rect 102876 537616 102928 537668
rect 132592 537616 132644 537668
rect 52368 537548 52420 537600
rect 82912 537548 82964 537600
rect 98368 537548 98420 537600
rect 128544 537548 128596 537600
rect 57796 537480 57848 537532
rect 74724 537480 74776 537532
rect 80336 537412 80388 537464
rect 81440 537412 81492 537464
rect 116584 537480 116636 537532
rect 83464 536800 83516 536852
rect 84844 536800 84896 536852
rect 35164 536732 35216 536784
rect 106096 536732 106148 536784
rect 111800 536528 111852 536580
rect 114744 536528 114796 536580
rect 38476 536052 38528 536104
rect 71320 536052 71372 536104
rect 106096 536052 106148 536104
rect 134156 536052 134208 536104
rect 71044 534964 71096 535016
rect 79692 534964 79744 535016
rect 101956 534964 102008 535016
rect 107936 534964 107988 535016
rect 56416 534896 56468 534948
rect 75184 534896 75236 534948
rect 97816 534896 97868 534948
rect 116124 534896 116176 534948
rect 42616 534828 42668 534880
rect 73252 534828 73304 534880
rect 89996 534828 90048 534880
rect 111984 534828 112036 534880
rect 50712 534760 50764 534812
rect 83556 534760 83608 534812
rect 95056 534760 95108 534812
rect 121552 534760 121604 534812
rect 45284 534692 45336 534744
rect 78404 534692 78456 534744
rect 93860 534692 93912 534744
rect 125784 534692 125836 534744
rect 97080 532176 97132 532228
rect 109224 532176 109276 532228
rect 93768 532108 93820 532160
rect 117504 532108 117556 532160
rect 87420 532040 87472 532092
rect 111800 532040 111852 532092
rect 92572 531972 92624 532024
rect 121644 531972 121696 532024
rect 49332 529252 49384 529304
rect 71964 529252 72016 529304
rect 46572 529184 46624 529236
rect 77116 529184 77168 529236
rect 3148 528504 3200 528556
rect 106924 528572 106976 528624
rect 116216 528572 116268 528624
rect 39764 525784 39816 525836
rect 68928 525716 68980 525768
rect 579804 525716 579856 525768
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 58624 512184 58676 512236
rect 59176 512184 59228 512236
rect 59176 511980 59228 512032
rect 580172 511912 580224 511964
rect 84200 500216 84252 500268
rect 117504 500216 117556 500268
rect 96436 497632 96488 497684
rect 118884 497632 118936 497684
rect 57612 497564 57664 497616
rect 77760 497564 77812 497616
rect 86776 497564 86828 497616
rect 117596 497564 117648 497616
rect 45376 497496 45428 497548
rect 72608 497496 72660 497548
rect 4804 497428 4856 497480
rect 91284 497496 91336 497548
rect 124220 497496 124272 497548
rect 135260 497496 135312 497548
rect 92572 497428 92624 497480
rect 133236 497428 133288 497480
rect 138020 497428 138072 497480
rect 118792 496748 118844 496800
rect 119068 496748 119120 496800
rect 56232 496204 56284 496256
rect 81440 496204 81492 496256
rect 89628 496136 89680 496188
rect 123116 496136 123168 496188
rect 124220 496136 124272 496188
rect 56324 496068 56376 496120
rect 75828 496068 75880 496120
rect 81440 496068 81492 496120
rect 88064 496068 88116 496120
rect 127072 496068 127124 496120
rect 133880 496068 133932 496120
rect 81440 495456 81492 495508
rect 110420 495456 110472 495508
rect 52092 494844 52144 494896
rect 73252 494844 73304 494896
rect 98644 494844 98696 494896
rect 112076 494844 112128 494896
rect 49516 494776 49568 494828
rect 74724 494776 74776 494828
rect 76104 494776 76156 494828
rect 82912 494776 82964 494828
rect 118792 494844 118844 494896
rect 3516 494708 3568 494760
rect 82820 494708 82872 494760
rect 97724 494708 97776 494760
rect 102140 494708 102192 494760
rect 95792 494640 95844 494692
rect 114560 494708 114612 494760
rect 123208 494776 123260 494828
rect 118792 494708 118844 494760
rect 118976 494708 119028 494760
rect 130016 494708 130068 494760
rect 85488 494368 85540 494420
rect 89628 494368 89680 494420
rect 80980 494096 81032 494148
rect 121460 494096 121512 494148
rect 41236 494028 41288 494080
rect 74540 494028 74592 494080
rect 76656 494028 76708 494080
rect 120356 494028 120408 494080
rect 82820 493960 82872 494012
rect 83556 493960 83608 494012
rect 124312 493960 124364 494012
rect 130108 493960 130160 494012
rect 129740 493892 129792 493944
rect 131212 493892 131264 493944
rect 90272 493416 90324 493468
rect 110696 493416 110748 493468
rect 54760 493348 54812 493400
rect 59268 493348 59320 493400
rect 68008 493348 68060 493400
rect 91928 493348 91980 493400
rect 95148 493348 95200 493400
rect 116032 493348 116084 493400
rect 43996 493280 44048 493332
rect 50804 493280 50856 493332
rect 70308 493280 70360 493332
rect 93216 493280 93268 493332
rect 129740 493280 129792 493332
rect 57704 492872 57756 492924
rect 75000 492872 75052 492924
rect 46848 492600 46900 492652
rect 52092 492804 52144 492856
rect 79324 492804 79376 492856
rect 59268 492736 59320 492788
rect 90272 492736 90324 492788
rect 92480 492736 92532 492788
rect 93768 492736 93820 492788
rect 114560 492736 114612 492788
rect 54944 492668 54996 492720
rect 57244 492600 57296 492652
rect 580356 492668 580408 492720
rect 87420 492600 87472 492652
rect 92480 492600 92532 492652
rect 46664 492464 46716 492516
rect 48044 492464 48096 492516
rect 93308 492124 93360 492176
rect 102232 492124 102284 492176
rect 53288 492056 53340 492108
rect 54484 492056 54536 492108
rect 70032 492056 70084 492108
rect 97908 492056 97960 492108
rect 111064 492056 111116 492108
rect 53472 491988 53524 492040
rect 55128 491988 55180 492040
rect 72240 491988 72292 492040
rect 97080 491988 97132 492040
rect 116308 491988 116360 492040
rect 48044 491920 48096 491972
rect 78036 491920 78088 491972
rect 81624 491920 81676 491972
rect 83004 491920 83056 491972
rect 113456 491920 113508 491972
rect 143540 491920 143592 491972
rect 96436 491784 96488 491836
rect 97908 491784 97960 491836
rect 68008 491648 68060 491700
rect 71136 491648 71188 491700
rect 86408 491580 86460 491632
rect 100668 491580 100720 491632
rect 82268 491512 82320 491564
rect 109132 491512 109184 491564
rect 52184 491444 52236 491496
rect 71780 491444 71832 491496
rect 89996 491376 90048 491428
rect 92848 491376 92900 491428
rect 99656 491376 99708 491428
rect 118792 491376 118844 491428
rect 119068 491376 119120 491428
rect 46756 491308 46808 491360
rect 80060 491308 80112 491360
rect 100668 491240 100720 491292
rect 125600 491240 125652 491292
rect 109132 491172 109184 491224
rect 123116 491172 123168 491224
rect 124496 491172 124548 491224
rect 125508 491172 125560 491224
rect 101864 491104 101916 491156
rect 109316 491104 109368 491156
rect 60372 490764 60424 490816
rect 86132 490764 86184 490816
rect 54852 490696 54904 490748
rect 83464 490696 83516 490748
rect 47952 490628 48004 490680
rect 79048 490628 79100 490680
rect 88984 490628 89036 490680
rect 101312 490628 101364 490680
rect 35808 490560 35860 490612
rect 37004 490560 37056 490612
rect 69756 490560 69808 490612
rect 94136 490560 94188 490612
rect 95056 490560 95108 490612
rect 109684 490560 109736 490612
rect 125508 490560 125560 490612
rect 580264 490560 580316 490612
rect 125600 490288 125652 490340
rect 127072 490288 127124 490340
rect 86960 489880 87012 489932
rect 101864 489880 101916 489932
rect 118792 489880 118844 489932
rect 124312 489880 124364 489932
rect 69848 489812 69900 489864
rect 70860 489812 70912 489864
rect 98736 489812 98788 489864
rect 99288 489812 99340 489864
rect 101312 489812 101364 489864
rect 122840 489812 122892 489864
rect 104256 489744 104308 489796
rect 118700 489744 118752 489796
rect 110328 489676 110380 489728
rect 113180 489676 113232 489728
rect 103336 488452 103388 488504
rect 117320 488452 117372 488504
rect 103428 488384 103480 488436
rect 109040 488384 109092 488436
rect 114468 488384 114520 488436
rect 123024 488384 123076 488436
rect 53564 487840 53616 487892
rect 59176 487840 59228 487892
rect 109040 487840 109092 487892
rect 116124 487840 116176 487892
rect 117320 487840 117372 487892
rect 125692 487840 125744 487892
rect 56508 487772 56560 487824
rect 67640 487772 67692 487824
rect 103520 487772 103572 487824
rect 134064 487772 134116 487824
rect 145012 487772 145064 487824
rect 59176 487160 59228 487212
rect 67732 487160 67784 487212
rect 34244 485732 34296 485784
rect 35164 485732 35216 485784
rect 67640 485800 67692 485852
rect 102324 485052 102376 485104
rect 112168 485052 112220 485104
rect 65892 484576 65944 484628
rect 68744 484576 68796 484628
rect 55036 484304 55088 484356
rect 57336 484304 57388 484356
rect 67640 484372 67692 484424
rect 113088 484372 113140 484424
rect 128452 484372 128504 484424
rect 102324 483624 102376 483676
rect 125600 483624 125652 483676
rect 126244 483624 126296 483676
rect 35624 482944 35676 482996
rect 64144 482944 64196 482996
rect 67640 483012 67692 483064
rect 102416 482944 102468 482996
rect 131764 482944 131816 482996
rect 146484 483012 146536 483064
rect 43812 482876 43864 482928
rect 68100 482876 68152 482928
rect 102324 482876 102376 482928
rect 106372 482876 106424 482928
rect 107476 482876 107528 482928
rect 107476 482264 107528 482316
rect 118792 482264 118844 482316
rect 102416 481584 102468 481636
rect 113364 481584 113416 481636
rect 120172 481584 120224 481636
rect 102324 481516 102376 481568
rect 110512 481516 110564 481568
rect 111708 481516 111760 481568
rect 111708 480904 111760 480956
rect 118700 480904 118752 480956
rect 55036 480224 55088 480276
rect 58624 480224 58676 480276
rect 39856 480156 39908 480208
rect 68560 480224 68612 480276
rect 102324 480156 102376 480208
rect 128360 480156 128412 480208
rect 58624 480088 58676 480140
rect 67640 480088 67692 480140
rect 63224 480020 63276 480072
rect 67732 480020 67784 480072
rect 128360 479476 128412 479528
rect 151912 479476 151964 479528
rect 61752 478864 61804 478916
rect 63224 478864 63276 478916
rect 111708 478252 111760 478304
rect 116032 478252 116084 478304
rect 107476 477572 107528 477624
rect 107844 477572 107896 477624
rect 102416 477504 102468 477556
rect 116032 477504 116084 477556
rect 100668 477436 100720 477488
rect 114652 477436 114704 477488
rect 108396 476144 108448 476196
rect 109224 476144 109276 476196
rect 39672 476076 39724 476128
rect 67640 476076 67692 476128
rect 102324 476076 102376 476128
rect 116032 476076 116084 476128
rect 102416 476008 102468 476060
rect 117412 476008 117464 476060
rect 117780 476008 117832 476060
rect 120080 476008 120132 476060
rect 102324 475940 102376 475992
rect 115940 475940 115992 475992
rect 99748 475668 99800 475720
rect 100760 475668 100812 475720
rect 53380 475328 53432 475380
rect 53748 475328 53800 475380
rect 67640 475328 67692 475380
rect 117780 475328 117832 475380
rect 132500 475328 132552 475380
rect 64696 474988 64748 475040
rect 67640 474988 67692 475040
rect 3424 474716 3476 474768
rect 7564 474716 7616 474768
rect 107384 474716 107436 474768
rect 107752 474716 107804 474768
rect 102324 474648 102376 474700
rect 125876 474648 125928 474700
rect 128360 474648 128412 474700
rect 61844 474308 61896 474360
rect 67640 474308 67692 474360
rect 102324 472744 102376 472796
rect 131120 472744 131172 472796
rect 103428 472676 103480 472728
rect 135168 472676 135220 472728
rect 102324 472608 102376 472660
rect 136824 472608 136876 472660
rect 140872 472608 140924 472660
rect 105544 472200 105596 472252
rect 110604 472200 110656 472252
rect 58992 471996 59044 472048
rect 66168 471996 66220 472048
rect 67640 471996 67692 472048
rect 67456 471928 67508 471980
rect 67732 471928 67784 471980
rect 102416 471928 102468 471980
rect 107384 471928 107436 471980
rect 135168 471248 135220 471300
rect 147772 471248 147824 471300
rect 107384 470976 107436 471028
rect 108304 470976 108356 471028
rect 30288 470568 30340 470620
rect 39304 470500 39356 470552
rect 67640 470568 67692 470620
rect 102784 470568 102836 470620
rect 139492 470568 139544 470620
rect 147772 470568 147824 470620
rect 580172 470568 580224 470620
rect 64788 470500 64840 470552
rect 66904 470500 66956 470552
rect 67732 470500 67784 470552
rect 42524 469820 42576 469872
rect 67180 469820 67232 469872
rect 67640 469820 67692 469872
rect 107016 469820 107068 469872
rect 121644 469820 121696 469872
rect 102324 469140 102376 469192
rect 120264 469140 120316 469192
rect 120264 468528 120316 468580
rect 129924 468528 129976 468580
rect 103520 468460 103572 468512
rect 138112 468460 138164 468512
rect 147680 468460 147732 468512
rect 64788 468120 64840 468172
rect 66076 468120 66128 468172
rect 67640 468120 67692 468172
rect 119988 467780 120040 467832
rect 123024 467780 123076 467832
rect 102784 466420 102836 466472
rect 102324 466352 102376 466404
rect 111892 466352 111944 466404
rect 112352 466352 112404 466404
rect 117228 466352 117280 466404
rect 128636 466352 128688 466404
rect 49608 465672 49660 465724
rect 67640 465672 67692 465724
rect 112352 465672 112404 465724
rect 119344 465672 119396 465724
rect 66168 465400 66220 465452
rect 67640 465400 67692 465452
rect 48044 464992 48096 465044
rect 49608 464992 49660 465044
rect 60464 464992 60516 465044
rect 61936 464992 61988 465044
rect 67732 464992 67784 465044
rect 102324 464992 102376 465044
rect 107476 464992 107528 465044
rect 142252 465060 142304 465112
rect 47860 464720 47912 464772
rect 48136 464720 48188 464772
rect 47860 464312 47912 464364
rect 67640 464312 67692 464364
rect 102416 463700 102468 463752
rect 113088 463700 113140 463752
rect 52000 463632 52052 463684
rect 52276 463632 52328 463684
rect 102324 463632 102376 463684
rect 115204 463632 115256 463684
rect 136824 463700 136876 463752
rect 52000 462952 52052 463004
rect 67640 462952 67692 463004
rect 3240 462340 3292 462392
rect 22744 462340 22796 462392
rect 102324 462272 102376 462324
rect 133972 462340 134024 462392
rect 102324 460912 102376 460964
rect 114652 460912 114704 460964
rect 50988 460232 51040 460284
rect 67640 460232 67692 460284
rect 115480 460232 115532 460284
rect 116216 460232 116268 460284
rect 126980 460232 127032 460284
rect 44456 460164 44508 460216
rect 45468 460164 45520 460216
rect 67732 460164 67784 460216
rect 102324 460164 102376 460216
rect 106188 460096 106240 460148
rect 115296 460096 115348 460148
rect 50804 459620 50856 459672
rect 50988 459620 51040 459672
rect 45468 459552 45520 459604
rect 62764 459552 62816 459604
rect 102876 459552 102928 459604
rect 67640 459484 67692 459536
rect 106188 459484 106240 459536
rect 136640 459484 136692 459536
rect 102324 459416 102376 459468
rect 115480 459416 115532 459468
rect 107752 458872 107804 458924
rect 142344 458872 142396 458924
rect 146392 458872 146444 458924
rect 34152 458804 34204 458856
rect 67272 458804 67324 458856
rect 103520 458804 103572 458856
rect 140964 458804 141016 458856
rect 149152 458804 149204 458856
rect 36912 458192 36964 458244
rect 44456 458192 44508 458244
rect 102416 458192 102468 458244
rect 115204 458192 115256 458244
rect 53656 458124 53708 458176
rect 68100 458124 68152 458176
rect 108488 458124 108540 458176
rect 114836 458124 114888 458176
rect 43904 457444 43956 457496
rect 67640 457444 67692 457496
rect 103520 457104 103572 457156
rect 107752 457104 107804 457156
rect 102232 455472 102284 455524
rect 105544 455472 105596 455524
rect 67640 455404 67692 455456
rect 102416 455404 102468 455456
rect 35716 455336 35768 455388
rect 40684 455336 40736 455388
rect 102232 455336 102284 455388
rect 107568 455336 107620 455388
rect 133788 455336 133840 455388
rect 139400 455336 139452 455388
rect 49608 454656 49660 454708
rect 54944 454656 54996 454708
rect 67732 454656 67784 454708
rect 48228 454044 48280 454096
rect 55128 454044 55180 454096
rect 67640 454044 67692 454096
rect 102232 453976 102284 454028
rect 124404 453976 124456 454028
rect 129832 453976 129884 454028
rect 102232 453364 102284 453416
rect 106096 453364 106148 453416
rect 50896 453296 50948 453348
rect 67640 453296 67692 453348
rect 34244 452616 34296 452668
rect 67732 452616 67784 452668
rect 68284 452616 68336 452668
rect 102232 452548 102284 452600
rect 136732 452548 136784 452600
rect 137100 452548 137152 452600
rect 42708 451868 42760 451920
rect 66996 451868 67048 451920
rect 103520 451868 103572 451920
rect 142160 451868 142212 451920
rect 150532 451868 150584 451920
rect 137100 451256 137152 451308
rect 142344 451256 142396 451308
rect 100852 450576 100904 450628
rect 105820 450576 105872 450628
rect 120080 450576 120132 450628
rect 107568 450508 107620 450560
rect 140780 450508 140832 450560
rect 44088 449828 44140 449880
rect 62764 449896 62816 449948
rect 67640 449896 67692 449948
rect 140780 449896 140832 449948
rect 143632 449896 143684 449948
rect 102416 449828 102468 449880
rect 107568 449828 107620 449880
rect 63408 449216 63460 449268
rect 67732 449216 67784 449268
rect 102140 449216 102192 449268
rect 107476 449216 107528 449268
rect 41144 449148 41196 449200
rect 67640 449148 67692 449200
rect 106188 449148 106240 449200
rect 134156 449148 134208 449200
rect 140780 449148 140832 449200
rect 107384 448604 107436 448656
rect 3148 448536 3200 448588
rect 46204 448536 46256 448588
rect 106924 448536 106976 448588
rect 107476 448536 107528 448588
rect 144920 448536 144972 448588
rect 61936 448468 61988 448520
rect 63316 448468 63368 448520
rect 67640 448468 67692 448520
rect 102140 448468 102192 448520
rect 106188 448468 106240 448520
rect 102416 448400 102468 448452
rect 107384 448400 107436 448452
rect 41144 447924 41196 447976
rect 42064 447924 42116 447976
rect 100024 447856 100076 447908
rect 112076 447856 112128 447908
rect 105728 447788 105780 447840
rect 118884 447788 118936 447840
rect 60648 445884 60700 445936
rect 64512 445884 64564 445936
rect 67640 445884 67692 445936
rect 102140 445816 102192 445868
rect 105544 445816 105596 445868
rect 37188 445680 37240 445732
rect 65524 445748 65576 445800
rect 67732 445748 67784 445800
rect 103520 445068 103572 445120
rect 133144 445136 133196 445188
rect 134064 445136 134116 445188
rect 38568 445000 38620 445052
rect 67640 445000 67692 445052
rect 102600 445000 102652 445052
rect 132592 445000 132644 445052
rect 136732 445000 136784 445052
rect 49424 444320 49476 444372
rect 67640 444320 67692 444372
rect 45192 443640 45244 443692
rect 49424 443640 49476 443692
rect 106096 443640 106148 443692
rect 117412 443640 117464 443692
rect 34336 443028 34388 443080
rect 37004 443028 37056 443080
rect 35716 442960 35768 443012
rect 38568 442960 38620 443012
rect 67732 442960 67784 443012
rect 39764 442892 39816 442944
rect 67640 442892 67692 442944
rect 102876 442824 102928 442876
rect 127164 442824 127216 442876
rect 127440 442824 127492 442876
rect 38568 442280 38620 442332
rect 39764 442280 39816 442332
rect 127440 442212 127492 442264
rect 143816 442212 143868 442264
rect 103336 441600 103388 441652
rect 139584 441600 139636 441652
rect 45376 440852 45428 440904
rect 69848 440648 69900 440700
rect 70400 440648 70452 440700
rect 72332 440648 72384 440700
rect 87696 440648 87748 440700
rect 88432 440648 88484 440700
rect 117596 440852 117648 440904
rect 62028 440308 62080 440360
rect 67548 440308 67600 440360
rect 67732 440308 67784 440360
rect 65984 440240 66036 440292
rect 71136 440240 71188 440292
rect 102876 440240 102928 440292
rect 138112 440240 138164 440292
rect 97448 440172 97500 440224
rect 98644 440172 98696 440224
rect 105728 440172 105780 440224
rect 57612 439492 57664 439544
rect 76012 439492 76064 439544
rect 77760 439492 77812 439544
rect 56232 439356 56284 439408
rect 57244 439356 57296 439408
rect 121920 439288 121972 439340
rect 122932 439288 122984 439340
rect 7564 439152 7616 439204
rect 96436 439152 96488 439204
rect 57244 439084 57296 439136
rect 80612 439084 80664 439136
rect 103060 439084 103112 439136
rect 136916 439084 136968 439136
rect 56416 439016 56468 439068
rect 74632 439016 74684 439068
rect 75828 439016 75880 439068
rect 97724 439016 97776 439068
rect 108396 439016 108448 439068
rect 41328 438948 41380 439000
rect 73896 438948 73948 439000
rect 88708 438948 88760 439000
rect 121552 438948 121604 439000
rect 72976 438880 73028 438932
rect 73436 438880 73488 438932
rect 93860 438880 93912 438932
rect 95148 438880 95200 438932
rect 22744 438812 22796 438864
rect 50712 438812 50764 438864
rect 96620 438880 96672 438932
rect 97724 438880 97776 438932
rect 108488 438880 108540 438932
rect 99656 438812 99708 438864
rect 121920 438812 121972 438864
rect 122196 438812 122248 438864
rect 45284 438744 45336 438796
rect 78404 438744 78456 438796
rect 99012 438744 99064 438796
rect 128544 438744 128596 438796
rect 46572 438676 46624 438728
rect 77116 438676 77168 438728
rect 96436 438676 96488 438728
rect 121736 438676 121788 438728
rect 59084 438608 59136 438660
rect 70032 438608 70084 438660
rect 93216 438608 93268 438660
rect 93768 438608 93820 438660
rect 107016 438608 107068 438660
rect 46204 438540 46256 438592
rect 99748 438540 99800 438592
rect 93676 438472 93728 438524
rect 102324 438472 102376 438524
rect 69388 438336 69440 438388
rect 71872 438336 71924 438388
rect 98368 438268 98420 438320
rect 99288 438268 99340 438320
rect 102232 438268 102284 438320
rect 65892 438200 65944 438252
rect 75184 438200 75236 438252
rect 50712 438132 50764 438184
rect 52184 438132 52236 438184
rect 83556 438132 83608 438184
rect 69296 437860 69348 437912
rect 70032 437860 70084 437912
rect 91100 437588 91152 437640
rect 92572 437588 92624 437640
rect 78404 437520 78456 437572
rect 80704 437520 80756 437572
rect 46572 437452 46624 437504
rect 46756 437452 46808 437504
rect 79048 437452 79100 437504
rect 80060 437452 80112 437504
rect 83648 437452 83700 437504
rect 84844 437452 84896 437504
rect 85028 437452 85080 437504
rect 86776 437452 86828 437504
rect 57520 437384 57572 437436
rect 91744 437384 91796 437436
rect 94504 437384 94556 437436
rect 125784 437384 125836 437436
rect 42616 437316 42668 437368
rect 73344 437316 73396 437368
rect 86224 437316 86276 437368
rect 100024 437316 100076 437368
rect 52368 437248 52420 437300
rect 82912 437248 82964 437300
rect 64144 436704 64196 436756
rect 75276 436704 75328 436756
rect 47952 436024 48004 436076
rect 80060 436024 80112 436076
rect 88248 436024 88300 436076
rect 111800 436024 111852 436076
rect 54852 435956 54904 436008
rect 83096 435956 83148 436008
rect 83648 435956 83700 436008
rect 60372 435888 60424 435940
rect 84200 435888 84252 435940
rect 85028 435888 85080 435940
rect 38476 434664 38528 434716
rect 71320 434664 71372 434716
rect 48964 433984 49016 434036
rect 76472 433984 76524 434036
rect 80704 431196 80756 431248
rect 580172 431196 580224 431248
rect 3424 429836 3476 429888
rect 100852 429836 100904 429888
rect 3516 422288 3568 422340
rect 48136 422288 48188 422340
rect 100668 422220 100720 422272
rect 124312 422220 124364 422272
rect 66996 419432 67048 419484
rect 67364 419432 67416 419484
rect 580172 419432 580224 419484
rect 56416 418752 56468 418804
rect 67364 418752 67416 418804
rect 91836 404336 91888 404388
rect 580172 404336 580224 404388
rect 108304 402364 108356 402416
rect 117596 402364 117648 402416
rect 96620 402296 96672 402348
rect 127164 402296 127216 402348
rect 88248 402228 88300 402280
rect 124312 402228 124364 402280
rect 108856 401616 108908 401668
rect 113456 401616 113508 401668
rect 74632 400188 74684 400240
rect 75276 400188 75328 400240
rect 162124 400188 162176 400240
rect 104164 399508 104216 399560
rect 138204 399508 138256 399560
rect 35164 399440 35216 399492
rect 75920 399440 75972 399492
rect 98644 399440 98696 399492
rect 135352 399440 135404 399492
rect 99380 398216 99432 398268
rect 118884 398216 118936 398268
rect 89628 398148 89680 398200
rect 122104 398148 122156 398200
rect 50988 398080 51040 398132
rect 99380 398080 99432 398132
rect 106924 398080 106976 398132
rect 141056 398080 141108 398132
rect 92480 397536 92532 397588
rect 92664 397536 92716 397588
rect 220084 397536 220136 397588
rect 3424 397468 3476 397520
rect 50988 397468 51040 397520
rect 65984 397468 66036 397520
rect 269764 397468 269816 397520
rect 46572 396856 46624 396908
rect 80060 396856 80112 396908
rect 105636 396856 105688 396908
rect 131304 396856 131356 396908
rect 53564 396788 53616 396840
rect 80704 396788 80756 396840
rect 91744 396788 91796 396840
rect 127256 396788 127308 396840
rect 46664 396720 46716 396772
rect 91928 396720 91980 396772
rect 93860 396720 93912 396772
rect 123116 396720 123168 396772
rect 53472 396040 53524 396092
rect 54484 396040 54536 396092
rect 84200 396040 84252 396092
rect 85120 396040 85172 396092
rect 166264 396040 166316 396092
rect 49516 395292 49568 395344
rect 88340 395292 88392 395344
rect 97908 395292 97960 395344
rect 121644 395292 121696 395344
rect 317420 395292 317472 395344
rect 70400 394952 70452 395004
rect 71136 394952 71188 395004
rect 39764 394884 39816 394936
rect 103704 394884 103756 394936
rect 104256 394884 104308 394936
rect 66076 394816 66128 394868
rect 142160 394816 142212 394868
rect 88340 394748 88392 394800
rect 170404 394748 170456 394800
rect 71136 394680 71188 394732
rect 214564 394680 214616 394732
rect 77944 394612 77996 394664
rect 91836 394612 91888 394664
rect 47860 394136 47912 394188
rect 56232 394136 56284 394188
rect 66076 394136 66128 394188
rect 52092 394068 52144 394120
rect 82912 394068 82964 394120
rect 47952 394000 48004 394052
rect 79324 394000 79376 394052
rect 43996 393932 44048 393984
rect 81440 393932 81492 393984
rect 87696 393932 87748 393984
rect 110420 393932 110472 393984
rect 43996 393456 44048 393508
rect 101404 393456 101456 393508
rect 81440 393388 81492 393440
rect 152004 393388 152056 393440
rect 75920 393320 75972 393372
rect 159364 393320 159416 393372
rect 110420 392776 110472 392828
rect 123208 392776 123260 392828
rect 96528 392708 96580 392760
rect 125876 392708 125928 392760
rect 57704 392640 57756 392692
rect 88432 392640 88484 392692
rect 96252 392640 96304 392692
rect 130016 392640 130068 392692
rect 140964 392640 141016 392692
rect 45284 392572 45336 392624
rect 78680 392572 78732 392624
rect 99288 392572 99340 392624
rect 135444 392572 135496 392624
rect 113088 392436 113140 392488
rect 114560 392436 114612 392488
rect 46848 392028 46900 392080
rect 92940 392028 92992 392080
rect 52276 391960 52328 392012
rect 110420 391960 110472 392012
rect 110972 391960 111024 392012
rect 111064 391960 111116 392012
rect 112076 391960 112128 392012
rect 113824 391960 113876 392012
rect 177304 391960 177356 392012
rect 60556 391484 60608 391536
rect 82820 391484 82872 391536
rect 54760 391348 54812 391400
rect 82820 391348 82872 391400
rect 100668 391348 100720 391400
rect 115388 391348 115440 391400
rect 60372 391280 60424 391332
rect 94504 391280 94556 391332
rect 102048 391280 102100 391332
rect 120356 391280 120408 391332
rect 41236 391212 41288 391264
rect 85948 391212 86000 391264
rect 94136 391212 94188 391264
rect 121460 391212 121512 391264
rect 147864 391212 147916 391264
rect 119344 390668 119396 390720
rect 124220 390668 124272 390720
rect 82912 390600 82964 390652
rect 83648 390600 83700 390652
rect 139400 390600 139452 390652
rect 82820 390532 82872 390584
rect 83004 390532 83056 390584
rect 143724 390532 143776 390584
rect 124128 389988 124180 390040
rect 135260 389988 135312 390040
rect 97448 389920 97500 389972
rect 130108 389920 130160 389972
rect 146300 389920 146352 389972
rect 53656 389852 53708 389904
rect 59268 389852 59320 389904
rect 104532 389852 104584 389904
rect 108948 389852 109000 389904
rect 131212 389852 131264 389904
rect 134156 389852 134208 389904
rect 49056 389784 49108 389836
rect 119344 389784 119396 389836
rect 106280 389240 106332 389292
rect 122840 389240 122892 389292
rect 124128 389240 124180 389292
rect 39856 389172 39908 389224
rect 71780 389172 71832 389224
rect 114376 389172 114428 389224
rect 142436 389172 142488 389224
rect 101404 389104 101456 389156
rect 103612 389104 103664 389156
rect 120632 389104 120684 389156
rect 127072 389104 127124 389156
rect 71872 388832 71924 388884
rect 72332 388832 72384 388884
rect 101864 388492 101916 388544
rect 113088 388492 113140 388544
rect 122288 388492 122340 388544
rect 57336 388424 57388 388476
rect 75828 388424 75880 388476
rect 107016 388424 107068 388476
rect 111708 388424 111760 388476
rect 124956 388424 125008 388476
rect 55036 388084 55088 388136
rect 69756 388084 69808 388136
rect 75184 388084 75236 388136
rect 75552 388084 75604 388136
rect 82452 388084 82504 388136
rect 109684 388084 109736 388136
rect 119344 388084 119396 388136
rect 59176 388016 59228 388068
rect 79324 388016 79376 388068
rect 100024 388016 100076 388068
rect 120632 388016 120684 388068
rect 56508 387948 56560 388000
rect 78036 387948 78088 388000
rect 91008 387948 91060 388000
rect 121920 387948 121972 388000
rect 25504 387880 25556 387932
rect 41236 387880 41288 387932
rect 72332 387880 72384 387932
rect 75828 387880 75880 387932
rect 113088 387880 113140 387932
rect 35808 387812 35860 387864
rect 80060 387812 80112 387864
rect 90272 387812 90324 387864
rect 98828 387812 98880 387864
rect 112076 387812 112128 387864
rect 188344 387812 188396 387864
rect 53748 387472 53800 387524
rect 56508 387472 56560 387524
rect 113088 387268 113140 387320
rect 132592 387268 132644 387320
rect 105544 387200 105596 387252
rect 131212 387200 131264 387252
rect 57612 387132 57664 387184
rect 74540 387132 74592 387184
rect 90916 387132 90968 387184
rect 125784 387132 125836 387184
rect 128636 387132 128688 387184
rect 143540 387132 143592 387184
rect 58900 387064 58952 387116
rect 90364 387064 90416 387116
rect 94872 387064 94924 387116
rect 108856 387064 108908 387116
rect 215944 387064 215996 387116
rect 52368 386452 52420 386504
rect 53472 386452 53524 386504
rect 80612 386452 80664 386504
rect 112904 386452 112956 386504
rect 128636 386452 128688 386504
rect 57888 386384 57940 386436
rect 87052 386384 87104 386436
rect 110328 386384 110380 386436
rect 136640 386384 136692 386436
rect 61752 386316 61804 386368
rect 68836 386316 68888 386368
rect 135260 386316 135312 386368
rect 138020 386316 138072 386368
rect 61660 385840 61712 385892
rect 73436 385840 73488 385892
rect 70308 385772 70360 385824
rect 83096 385772 83148 385824
rect 59084 385704 59136 385756
rect 56324 385636 56376 385688
rect 73436 385636 73488 385688
rect 112996 385704 113048 385756
rect 122932 385704 122984 385756
rect 82452 385636 82504 385688
rect 303620 385636 303672 385688
rect 86316 385568 86368 385620
rect 117320 385432 117372 385484
rect 117688 385432 117740 385484
rect 56508 385024 56560 385076
rect 77484 385296 77536 385348
rect 102600 385296 102652 385348
rect 107568 385296 107620 385348
rect 135260 385092 135312 385144
rect 133880 385024 133932 385076
rect 134616 385024 134668 385076
rect 117412 384888 117464 384940
rect 118240 384888 118292 384940
rect 121460 384888 121512 384940
rect 117412 384548 117464 384600
rect 34336 383664 34388 383716
rect 68744 383664 68796 383716
rect 116676 383664 116728 383716
rect 130016 383664 130068 383716
rect 116768 383596 116820 383648
rect 125692 383596 125744 383648
rect 121460 382916 121512 382968
rect 349252 382916 349304 382968
rect 44088 382236 44140 382288
rect 67732 382236 67784 382288
rect 62028 382168 62080 382220
rect 67640 382168 67692 382220
rect 117320 382168 117372 382220
rect 145012 382168 145064 382220
rect 145012 381488 145064 381540
rect 206284 381488 206336 381540
rect 64420 380808 64472 380860
rect 67456 380808 67508 380860
rect 117320 380808 117372 380860
rect 128452 380808 128504 380860
rect 64696 380740 64748 380792
rect 68008 380740 68060 380792
rect 50712 380672 50764 380724
rect 53380 380672 53432 380724
rect 67640 380672 67692 380724
rect 117688 380128 117740 380180
rect 126244 380128 126296 380180
rect 128452 379516 128504 379568
rect 129740 379516 129792 379568
rect 33048 378768 33100 378820
rect 47860 378768 47912 378820
rect 60280 378768 60332 378820
rect 70308 378768 70360 378820
rect 118608 378768 118660 378820
rect 125692 378768 125744 378820
rect 47860 378156 47912 378208
rect 48228 378156 48280 378208
rect 67640 378156 67692 378208
rect 124864 378156 124916 378208
rect 580172 378156 580224 378208
rect 58992 377408 59044 377460
rect 59176 377408 59228 377460
rect 67640 377408 67692 377460
rect 118608 377408 118660 377460
rect 121460 377408 121512 377460
rect 146484 377408 146536 377460
rect 66076 376660 66128 376712
rect 68376 376660 68428 376712
rect 118608 376048 118660 376100
rect 128452 376048 128504 376100
rect 49516 375980 49568 376032
rect 59176 375980 59228 376032
rect 118516 375980 118568 376032
rect 120172 375980 120224 376032
rect 143540 375980 143592 376032
rect 64696 375300 64748 375352
rect 66904 375300 66956 375352
rect 67640 375300 67692 375352
rect 118608 375300 118660 375352
rect 151912 375300 151964 375352
rect 153108 375300 153160 375352
rect 153108 374620 153160 374672
rect 202144 374620 202196 374672
rect 42524 373940 42576 373992
rect 66904 373940 66956 373992
rect 67732 374008 67784 374060
rect 117504 373328 117556 373380
rect 123852 373328 123904 373380
rect 118424 372580 118476 372632
rect 222936 372580 222988 372632
rect 3240 372512 3292 372564
rect 49056 372512 49108 372564
rect 64788 372512 64840 372564
rect 67640 372512 67692 372564
rect 119988 371900 120040 371952
rect 122932 371900 122984 371952
rect 63224 371220 63276 371272
rect 67456 371220 67508 371272
rect 67640 371220 67692 371272
rect 118608 371220 118660 371272
rect 273996 371220 274048 371272
rect 56232 369792 56284 369844
rect 67640 369792 67692 369844
rect 66168 369112 66220 369164
rect 67732 369112 67784 369164
rect 118976 368500 119028 368552
rect 127072 368500 127124 368552
rect 131672 368432 131724 368484
rect 132500 368432 132552 368484
rect 52000 367752 52052 367804
rect 61476 367752 61528 367804
rect 119344 367752 119396 367804
rect 128360 367752 128412 367804
rect 118608 367208 118660 367260
rect 119344 367208 119396 367260
rect 37188 367072 37240 367124
rect 60464 367072 60516 367124
rect 63408 367072 63460 367124
rect 67640 367072 67692 367124
rect 118516 367072 118568 367124
rect 131672 367072 131724 367124
rect 61384 367004 61436 367056
rect 67732 367004 67784 367056
rect 118608 367004 118660 367056
rect 131120 367004 131172 367056
rect 116032 366936 116084 366988
rect 122932 366936 122984 366988
rect 61476 366324 61528 366376
rect 67640 366324 67692 366376
rect 131120 365712 131172 365764
rect 132500 365712 132552 365764
rect 118700 365100 118752 365152
rect 140872 365100 140924 365152
rect 121552 365032 121604 365084
rect 147772 365032 147824 365084
rect 122932 364964 122984 365016
rect 580264 364964 580316 365016
rect 118608 364760 118660 364812
rect 121552 364760 121604 364812
rect 50804 363672 50856 363724
rect 67640 363672 67692 363724
rect 36912 363604 36964 363656
rect 67732 363604 67784 363656
rect 36912 362924 36964 362976
rect 37096 362924 37148 362976
rect 50620 362924 50672 362976
rect 50804 362924 50856 362976
rect 117964 362856 118016 362908
rect 151820 362856 151872 362908
rect 153108 362856 153160 362908
rect 34152 362176 34204 362228
rect 60740 362176 60792 362228
rect 118608 362176 118660 362228
rect 122104 362176 122156 362228
rect 139492 362176 139544 362228
rect 60740 361632 60792 361684
rect 61752 361632 61804 361684
rect 67640 361632 67692 361684
rect 43812 361564 43864 361616
rect 69204 361564 69256 361616
rect 43904 360816 43956 360868
rect 59176 360816 59228 360868
rect 116676 360272 116728 360324
rect 117228 360272 117280 360324
rect 45468 360136 45520 360188
rect 65616 360204 65668 360256
rect 67640 360204 67692 360256
rect 118608 360204 118660 360256
rect 120172 360204 120224 360256
rect 132684 360204 132736 360256
rect 118148 360136 118200 360188
rect 147680 360136 147732 360188
rect 120172 360068 120224 360120
rect 120724 360068 120776 360120
rect 129924 360068 129976 360120
rect 61476 359524 61528 359576
rect 61844 359524 61896 359576
rect 59176 359456 59228 359508
rect 67640 359456 67692 359508
rect 147680 359456 147732 359508
rect 198004 359456 198056 359508
rect 118608 358436 118660 358488
rect 124220 358436 124272 358488
rect 54852 358028 54904 358080
rect 55128 358028 55180 358080
rect 67640 358028 67692 358080
rect 3148 357416 3200 357468
rect 22744 357416 22796 357468
rect 40684 357348 40736 357400
rect 62856 357416 62908 357468
rect 67732 357416 67784 357468
rect 115296 357348 115348 357400
rect 117320 357348 117372 357400
rect 117688 357008 117740 357060
rect 121644 357008 121696 357060
rect 122196 356736 122248 356788
rect 128360 356736 128412 356788
rect 50896 356668 50948 356720
rect 60648 356668 60700 356720
rect 124956 356668 125008 356720
rect 325700 356668 325752 356720
rect 60648 356124 60700 356176
rect 67732 356124 67784 356176
rect 34152 356056 34204 356108
rect 69480 356056 69532 356108
rect 118608 355988 118660 356040
rect 142252 355988 142304 356040
rect 143448 355988 143500 356040
rect 63500 355308 63552 355360
rect 67640 355308 67692 355360
rect 143448 355308 143500 355360
rect 233884 355308 233936 355360
rect 118608 354628 118660 354680
rect 133972 354628 134024 354680
rect 121644 353948 121696 354000
rect 324412 353948 324464 354000
rect 133972 353336 134024 353388
rect 138020 353336 138072 353388
rect 56416 353200 56468 353252
rect 66996 353200 67048 353252
rect 67640 353268 67692 353320
rect 118056 353268 118108 353320
rect 133880 353268 133932 353320
rect 136824 353268 136876 353320
rect 11704 352520 11756 352572
rect 34244 352520 34296 352572
rect 41420 352520 41472 352572
rect 62764 352520 62816 352572
rect 67916 352520 67968 352572
rect 41420 351908 41472 351960
rect 42708 351908 42760 351960
rect 67640 351908 67692 351960
rect 116584 351296 116636 351348
rect 128452 351296 128504 351348
rect 118424 351228 118476 351280
rect 204904 351228 204956 351280
rect 64604 351160 64656 351212
rect 67732 351160 67784 351212
rect 118516 351160 118568 351212
rect 271236 351160 271288 351212
rect 118608 349868 118660 349920
rect 124404 349868 124456 349920
rect 126980 349868 127032 349920
rect 63316 349800 63368 349852
rect 68008 349800 68060 349852
rect 126244 349800 126296 349852
rect 314660 349800 314712 349852
rect 42064 349120 42116 349172
rect 45468 349120 45520 349172
rect 67640 349120 67692 349172
rect 61936 348372 61988 348424
rect 68836 348372 68888 348424
rect 118608 347828 118660 347880
rect 140872 347828 140924 347880
rect 117780 347760 117832 347812
rect 258724 347760 258776 347812
rect 117412 347692 117464 347744
rect 133788 347692 133840 347744
rect 140872 347692 140924 347744
rect 149244 347692 149296 347744
rect 133788 347080 133840 347132
rect 191104 347080 191156 347132
rect 3332 347012 3384 347064
rect 25504 347012 25556 347064
rect 64512 347012 64564 347064
rect 68560 347012 68612 347064
rect 149244 347012 149296 347064
rect 316132 347012 316184 347064
rect 65524 346400 65576 346452
rect 67640 346400 67692 346452
rect 22744 346332 22796 346384
rect 35716 346332 35768 346384
rect 118608 346332 118660 346384
rect 146392 346332 146444 346384
rect 146760 346332 146812 346384
rect 35716 345652 35768 345704
rect 63316 345652 63368 345704
rect 118332 345652 118384 345704
rect 122932 345652 122984 345704
rect 131304 345652 131356 345704
rect 146760 345652 146812 345704
rect 217232 345652 217284 345704
rect 63316 345040 63368 345092
rect 67732 345040 67784 345092
rect 116676 345040 116728 345092
rect 124312 345040 124364 345092
rect 66076 344972 66128 345024
rect 67640 344972 67692 345024
rect 118608 344972 118660 345024
rect 149060 344972 149112 345024
rect 149060 344292 149112 344344
rect 331864 344292 331916 344344
rect 63500 343680 63552 343732
rect 67732 343680 67784 343732
rect 45192 343612 45244 343664
rect 47860 343612 47912 343664
rect 67640 343612 67692 343664
rect 118608 343544 118660 343596
rect 150440 343544 150492 343596
rect 128728 342932 128780 342984
rect 129832 342932 129884 342984
rect 37004 342864 37056 342916
rect 41144 342864 41196 342916
rect 63500 342864 63552 342916
rect 150440 342864 150492 342916
rect 282184 342864 282236 342916
rect 115296 342320 115348 342372
rect 118792 342320 118844 342372
rect 118148 342252 118200 342304
rect 128728 342252 128780 342304
rect 118608 341504 118660 341556
rect 142344 341504 142396 341556
rect 38568 340824 38620 340876
rect 65984 340892 66036 340944
rect 67640 340892 67692 340944
rect 118056 340824 118108 340876
rect 118792 340892 118844 340944
rect 120080 340892 120132 340944
rect 140872 340892 140924 340944
rect 580264 340892 580316 340944
rect 117780 340756 117832 340808
rect 150532 340824 150584 340876
rect 151544 340824 151596 340876
rect 151544 340144 151596 340196
rect 352564 340144 352616 340196
rect 113916 339600 113968 339652
rect 115112 339600 115164 339652
rect 143632 339600 143684 339652
rect 61660 339532 61712 339584
rect 73252 339532 73304 339584
rect 113824 339532 113876 339584
rect 140780 339532 140832 339584
rect 48044 339464 48096 339516
rect 71964 339464 72016 339516
rect 48964 339396 49016 339448
rect 76656 339396 76708 339448
rect 77116 339396 77168 339448
rect 87420 339396 87472 339448
rect 87604 339396 87656 339448
rect 580356 339396 580408 339448
rect 56324 339328 56376 339380
rect 73896 339328 73948 339380
rect 74448 339328 74500 339380
rect 124864 339328 124916 339380
rect 58900 339260 58952 339312
rect 93216 339260 93268 339312
rect 113180 339260 113232 339312
rect 114008 339260 114060 339312
rect 144920 339260 144972 339312
rect 54944 339192 54996 339244
rect 57244 339192 57296 339244
rect 82268 339192 82320 339244
rect 100300 339192 100352 339244
rect 125600 339192 125652 339244
rect 125876 339192 125928 339244
rect 102232 339056 102284 339108
rect 103336 339056 103388 339108
rect 127164 339124 127216 339176
rect 66076 338784 66128 338836
rect 80704 338784 80756 338836
rect 62856 338716 62908 338768
rect 97264 338716 97316 338768
rect 104164 338716 104216 338768
rect 120724 338716 120776 338768
rect 91008 338104 91060 338156
rect 91928 338104 91980 338156
rect 70032 338036 70084 338088
rect 72976 338036 73028 338088
rect 75828 338036 75880 338088
rect 79968 338036 80020 338088
rect 108028 338036 108080 338088
rect 143816 338036 143868 338088
rect 47952 337968 48004 338020
rect 83556 337968 83608 338020
rect 115756 337968 115808 338020
rect 141056 337968 141108 338020
rect 141332 337968 141384 338020
rect 61384 337900 61436 337952
rect 84200 337900 84252 337952
rect 97724 337900 97776 337952
rect 128452 337900 128504 337952
rect 57612 337832 57664 337884
rect 76472 337832 76524 337884
rect 95792 337832 95844 337884
rect 125784 337832 125836 337884
rect 126888 337832 126940 337884
rect 86776 337764 86828 337816
rect 120448 337764 120500 337816
rect 57888 337696 57940 337748
rect 60372 337696 60424 337748
rect 98368 337696 98420 337748
rect 105544 337696 105596 337748
rect 108028 337696 108080 337748
rect 80980 337628 81032 337680
rect 81440 337628 81492 337680
rect 141332 337424 141384 337476
rect 196624 337424 196676 337476
rect 66996 337356 67048 337408
rect 77300 337356 77352 337408
rect 99656 337356 99708 337408
rect 103428 337356 103480 337408
rect 123116 337356 123168 337408
rect 126888 337356 126940 337408
rect 276664 337356 276716 337408
rect 102876 337220 102928 337272
rect 104900 337220 104952 337272
rect 103520 337016 103572 337068
rect 109132 337016 109184 337068
rect 92572 336812 92624 336864
rect 95240 336812 95292 336864
rect 71964 336744 72016 336796
rect 75184 336744 75236 336796
rect 81624 336744 81676 336796
rect 100024 336744 100076 336796
rect 112444 336744 112496 336796
rect 113824 336744 113876 336796
rect 128452 336744 128504 336796
rect 180064 336744 180116 336796
rect 41328 336676 41380 336728
rect 74540 336676 74592 336728
rect 75276 336676 75328 336728
rect 91284 336676 91336 336728
rect 92388 336676 92440 336728
rect 46756 336608 46808 336660
rect 78680 336608 78732 336660
rect 107568 336676 107620 336728
rect 139584 336676 139636 336728
rect 116676 336608 116728 336660
rect 126980 336608 127032 336660
rect 128544 336608 128596 336660
rect 59084 336540 59136 336592
rect 88984 336540 89036 336592
rect 109868 336540 109920 336592
rect 134064 336540 134116 336592
rect 53564 336472 53616 336524
rect 79324 336472 79376 336524
rect 56416 336404 56468 336456
rect 60556 336404 60608 336456
rect 84752 336404 84804 336456
rect 109132 335996 109184 336048
rect 126980 335996 127032 336048
rect 45284 335248 45336 335300
rect 81624 335248 81676 335300
rect 108304 335248 108356 335300
rect 136732 335248 136784 335300
rect 42616 335180 42668 335232
rect 70400 335180 70452 335232
rect 104808 335180 104860 335232
rect 128360 335180 128412 335232
rect 60556 335112 60608 335164
rect 87604 335112 87656 335164
rect 112536 335112 112588 335164
rect 113088 335112 113140 335164
rect 131212 335112 131264 335164
rect 57612 334636 57664 334688
rect 104808 334636 104860 334688
rect 62028 334568 62080 334620
rect 109868 334568 109920 334620
rect 70400 333956 70452 334008
rect 71044 333956 71096 334008
rect 46572 333888 46624 333940
rect 81440 333888 81492 333940
rect 95148 333888 95200 333940
rect 127256 333888 127308 333940
rect 52184 333820 52236 333872
rect 86224 333820 86276 333872
rect 104900 333820 104952 333872
rect 135444 333820 135496 333872
rect 107660 333276 107712 333328
rect 128636 333276 128688 333328
rect 61752 333208 61804 333260
rect 115204 333208 115256 333260
rect 135444 333208 135496 333260
rect 293960 333208 294012 333260
rect 81440 332596 81492 332648
rect 82084 332596 82136 332648
rect 94596 332596 94648 332648
rect 95148 332596 95200 332648
rect 57704 332528 57756 332580
rect 90364 332528 90416 332580
rect 94504 332528 94556 332580
rect 125784 332528 125836 332580
rect 128452 332528 128504 332580
rect 63316 331916 63368 331968
rect 98000 331916 98052 331968
rect 106280 331916 106332 331968
rect 118700 331916 118752 331968
rect 67456 331848 67508 331900
rect 338120 331848 338172 331900
rect 105452 331168 105504 331220
rect 136916 331168 136968 331220
rect 137192 331168 137244 331220
rect 137192 330488 137244 330540
rect 336004 330488 336056 330540
rect 110604 329740 110656 329792
rect 133144 329740 133196 329792
rect 133788 329740 133840 329792
rect 79968 329060 80020 329112
rect 342260 329060 342312 329112
rect 97080 328380 97132 328432
rect 129832 328380 129884 328432
rect 130568 328380 130620 328432
rect 49608 327768 49660 327820
rect 105544 327768 105596 327820
rect 106096 327768 106148 327820
rect 114468 327768 114520 327820
rect 138112 327768 138164 327820
rect 68836 327700 68888 327752
rect 251180 327700 251232 327752
rect 3424 327088 3476 327140
rect 49608 327088 49660 327140
rect 130568 327088 130620 327140
rect 333980 327088 334032 327140
rect 68652 326476 68704 326528
rect 115388 326476 115440 326528
rect 106188 326408 106240 326460
rect 116124 326408 116176 326460
rect 68928 326340 68980 326392
rect 309784 326340 309836 326392
rect 72424 324980 72476 325032
rect 108304 324980 108356 325032
rect 73344 324912 73396 324964
rect 116032 324912 116084 324964
rect 91008 324232 91060 324284
rect 124312 324232 124364 324284
rect 128544 324232 128596 324284
rect 86316 323552 86368 323604
rect 113916 323552 113968 323604
rect 66904 322192 66956 322244
rect 309140 322192 309192 322244
rect 93952 320832 94004 320884
rect 125692 320832 125744 320884
rect 118056 320492 118108 320544
rect 120264 320492 120316 320544
rect 100944 320084 100996 320136
rect 135352 320084 135404 320136
rect 136548 320084 136600 320136
rect 111248 320016 111300 320068
rect 138204 320016 138256 320068
rect 138664 320016 138716 320068
rect 94044 319472 94096 319524
rect 112444 319472 112496 319524
rect 136548 319472 136600 319524
rect 267004 319472 267056 319524
rect 75276 319404 75328 319456
rect 114560 319404 114612 319456
rect 138664 319404 138716 319456
rect 339500 319404 339552 319456
rect 101404 318248 101456 318300
rect 127072 318248 127124 318300
rect 67548 318180 67600 318232
rect 115296 318180 115348 318232
rect 75184 318112 75236 318164
rect 311900 318112 311952 318164
rect 84844 318044 84896 318096
rect 345020 318044 345072 318096
rect 93216 316752 93268 316804
rect 113824 316752 113876 316804
rect 71136 316684 71188 316736
rect 320180 316684 320232 316736
rect 152004 315936 152056 315988
rect 580356 315936 580408 315988
rect 120724 315256 120776 315308
rect 152004 315256 152056 315308
rect 57704 313964 57756 314016
rect 118792 313964 118844 314016
rect 88984 313896 89036 313948
rect 216036 313896 216088 313948
rect 91100 313284 91152 313336
rect 121644 313284 121696 313336
rect 582564 313284 582616 313336
rect 80060 312604 80112 312656
rect 91100 312604 91152 312656
rect 97264 312604 97316 312656
rect 125784 312604 125836 312656
rect 126888 312604 126940 312656
rect 89076 312536 89128 312588
rect 209044 312536 209096 312588
rect 126888 311856 126940 311908
rect 579988 311856 580040 311908
rect 3516 311788 3568 311840
rect 50712 311788 50764 311840
rect 50712 311108 50764 311160
rect 115940 311108 115992 311160
rect 74448 309816 74500 309868
rect 119712 309816 119764 309868
rect 83464 309748 83516 309800
rect 322204 309748 322256 309800
rect 88340 309136 88392 309188
rect 280804 309136 280856 309188
rect 113088 308388 113140 308440
rect 253940 308388 253992 308440
rect 74632 307912 74684 307964
rect 145564 307912 145616 307964
rect 81440 307844 81492 307896
rect 155224 307844 155276 307896
rect 78772 307776 78824 307828
rect 226984 307776 227036 307828
rect 79324 307164 79376 307216
rect 120080 307164 120132 307216
rect 65616 307096 65668 307148
rect 213184 307096 213236 307148
rect 103336 307028 103388 307080
rect 266360 307028 266412 307080
rect 3516 306280 3568 306332
rect 11704 306280 11756 306332
rect 71044 305668 71096 305720
rect 186964 305668 187016 305720
rect 100024 305600 100076 305652
rect 321560 305600 321612 305652
rect 89720 304988 89772 305040
rect 171784 304988 171836 305040
rect 80704 304308 80756 304360
rect 129832 304308 129884 304360
rect 48136 304240 48188 304292
rect 71780 304240 71832 304292
rect 109684 304240 109736 304292
rect 119344 304240 119396 304292
rect 582840 304240 582892 304292
rect 75920 303764 75972 303816
rect 163504 303764 163556 303816
rect 66168 303696 66220 303748
rect 169024 303696 169076 303748
rect 85580 303628 85632 303680
rect 278044 303628 278096 303680
rect 65984 302880 66036 302932
rect 131120 302880 131172 302932
rect 87512 302404 87564 302456
rect 222844 302404 222896 302456
rect 85672 302336 85724 302388
rect 231124 302336 231176 302388
rect 112444 302268 112496 302320
rect 272524 302268 272576 302320
rect 71872 302200 71924 302252
rect 309232 302200 309284 302252
rect 90364 301520 90416 301572
rect 195244 301520 195296 301572
rect 71044 301452 71096 301504
rect 134156 301452 134208 301504
rect 582656 301452 582708 301504
rect 84200 301044 84252 301096
rect 180156 301044 180208 301096
rect 106924 300976 106976 301028
rect 203524 300976 203576 301028
rect 74540 300908 74592 300960
rect 240416 300908 240468 300960
rect 110972 300840 111024 300892
rect 302332 300840 302384 300892
rect 93124 300296 93176 300348
rect 125876 300296 125928 300348
rect 86224 300228 86276 300280
rect 124312 300228 124364 300280
rect 61936 300160 61988 300212
rect 116584 300160 116636 300212
rect 42708 300092 42760 300144
rect 123116 300092 123168 300144
rect 81900 299548 81952 299600
rect 198188 299548 198240 299600
rect 102140 299480 102192 299532
rect 224224 299480 224276 299532
rect 61844 298732 61896 298784
rect 127164 298732 127216 298784
rect 73252 298392 73304 298444
rect 157984 298392 158036 298444
rect 82912 298324 82964 298376
rect 178776 298324 178828 298376
rect 75184 298256 75236 298308
rect 227076 298256 227128 298308
rect 102876 298188 102928 298240
rect 262220 298188 262272 298240
rect 103428 298120 103480 298172
rect 104808 298120 104860 298172
rect 106188 298120 106240 298172
rect 582380 298120 582432 298172
rect 48044 297508 48096 297560
rect 77760 297508 77812 297560
rect 60464 297440 60516 297492
rect 124404 297440 124456 297492
rect 41236 297372 41288 297424
rect 117228 297372 117280 297424
rect 117964 296964 118016 297016
rect 123024 296964 123076 297016
rect 88708 296896 88760 296948
rect 151084 296896 151136 296948
rect 100944 296828 100996 296880
rect 182824 296828 182876 296880
rect 93216 296760 93268 296812
rect 202236 296760 202288 296812
rect 110604 296692 110656 296744
rect 225604 296692 225656 296744
rect 29644 295740 29696 295792
rect 118056 295740 118108 295792
rect 91928 295672 91980 295724
rect 141424 295672 141476 295724
rect 117688 295604 117740 295656
rect 199384 295604 199436 295656
rect 83556 295536 83608 295588
rect 181444 295536 181496 295588
rect 99656 295468 99708 295520
rect 256700 295468 256752 295520
rect 68836 295400 68888 295452
rect 234620 295400 234672 295452
rect 17224 295332 17276 295384
rect 92572 295332 92624 295384
rect 92940 295332 92992 295384
rect 111892 295332 111944 295384
rect 307852 295332 307904 295384
rect 87420 294788 87472 294840
rect 106924 294788 106976 294840
rect 25504 294584 25556 294636
rect 53656 294584 53708 294636
rect 79048 294720 79100 294772
rect 84844 294720 84896 294772
rect 104164 294720 104216 294772
rect 57796 294652 57848 294704
rect 91284 294652 91336 294704
rect 70676 294584 70728 294636
rect 115848 294584 115900 294636
rect 106740 294380 106792 294432
rect 112444 294380 112496 294432
rect 71780 294312 71832 294364
rect 72332 294312 72384 294364
rect 85488 294312 85540 294364
rect 86316 294312 86368 294364
rect 93952 294312 94004 294364
rect 94780 294312 94832 294364
rect 108028 294312 108080 294364
rect 117136 294312 117188 294364
rect 71320 294244 71372 294296
rect 72424 294244 72476 294296
rect 85580 294244 85632 294296
rect 86500 294244 86552 294296
rect 105452 294244 105504 294296
rect 125508 294244 125560 294296
rect 113824 294176 113876 294228
rect 152464 294176 152516 294228
rect 112536 294108 112588 294160
rect 255320 294108 255372 294160
rect 80980 294040 81032 294092
rect 239036 294040 239088 294092
rect 47584 293972 47636 294024
rect 101404 293972 101456 294024
rect 101588 293972 101640 294024
rect 104164 293972 104216 294024
rect 110420 293972 110472 294024
rect 117228 293972 117280 294024
rect 119620 293972 119672 294024
rect 119344 293904 119396 293956
rect 303712 293972 303764 294024
rect 125508 293904 125560 293956
rect 130016 293904 130068 293956
rect 115204 293292 115256 293344
rect 125692 293292 125744 293344
rect 53104 293224 53156 293276
rect 54484 293224 54536 293276
rect 97080 293224 97132 293276
rect 110420 293224 110472 293276
rect 278136 293224 278188 293276
rect 93860 292748 93912 292800
rect 133144 292748 133196 292800
rect 77116 292680 77168 292732
rect 125232 292680 125284 292732
rect 125508 292680 125560 292732
rect 103520 292612 103572 292664
rect 271144 292612 271196 292664
rect 55128 292544 55180 292596
rect 96436 292544 96488 292596
rect 97724 292544 97776 292596
rect 273904 292544 273956 292596
rect 121644 292476 121696 292528
rect 147864 292476 147916 292528
rect 125508 292408 125560 292460
rect 142436 292408 142488 292460
rect 117136 291932 117188 291984
rect 109592 291864 109644 291916
rect 117320 291864 117372 291916
rect 166356 291864 166408 291916
rect 307944 291796 307996 291848
rect 290464 291184 290516 291236
rect 32404 290436 32456 290488
rect 67640 290436 67692 290488
rect 121644 289824 121696 289876
rect 234712 289824 234764 289876
rect 66168 289756 66220 289808
rect 68192 289756 68244 289808
rect 121736 288396 121788 288448
rect 287336 288396 287388 288448
rect 49516 288328 49568 288380
rect 67640 288328 67692 288380
rect 121644 288328 121696 288380
rect 140964 288328 141016 288380
rect 141608 288328 141660 288380
rect 141608 287648 141660 287700
rect 467104 287648 467156 287700
rect 121828 287036 121880 287088
rect 224316 287036 224368 287088
rect 121736 286900 121788 286952
rect 125876 286900 125928 286952
rect 121644 286832 121696 286884
rect 132684 286832 132736 286884
rect 121552 286628 121604 286680
rect 123116 286628 123168 286680
rect 125876 286288 125928 286340
rect 468484 286288 468536 286340
rect 46756 284316 46808 284368
rect 67640 284316 67692 284368
rect 121644 284316 121696 284368
rect 214656 284316 214708 284368
rect 56508 284248 56560 284300
rect 67732 284248 67784 284300
rect 121552 284248 121604 284300
rect 143724 284248 143776 284300
rect 121552 282888 121604 282940
rect 282920 282888 282972 282940
rect 43996 282820 44048 282872
rect 67640 282820 67692 282872
rect 222936 282140 222988 282192
rect 336740 282140 336792 282192
rect 121644 281596 121696 281648
rect 221464 281596 221516 281648
rect 121552 281528 121604 281580
rect 227168 281528 227220 281580
rect 50804 280168 50856 280220
rect 67640 280168 67692 280220
rect 121552 280168 121604 280220
rect 284576 280168 284628 280220
rect 33140 280100 33192 280152
rect 34152 280100 34204 280152
rect 67732 280100 67784 280152
rect 55036 280032 55088 280084
rect 67640 280032 67692 280084
rect 4804 279420 4856 279472
rect 33140 279420 33192 279472
rect 271236 279420 271288 279472
rect 346400 279420 346452 279472
rect 121552 278808 121604 278860
rect 204996 278808 205048 278860
rect 121644 278740 121696 278792
rect 269856 278740 269908 278792
rect 273996 277992 274048 278044
rect 347780 277992 347832 278044
rect 55036 277448 55088 277500
rect 67640 277448 67692 277500
rect 121552 277448 121604 277500
rect 192484 277448 192536 277500
rect 52092 277380 52144 277432
rect 67732 277380 67784 277432
rect 121644 277380 121696 277432
rect 302240 277380 302292 277432
rect 121552 276632 121604 276684
rect 129924 276632 129976 276684
rect 53564 276020 53616 276072
rect 67640 276020 67692 276072
rect 129924 276020 129976 276072
rect 130384 276020 130436 276072
rect 61844 274728 61896 274780
rect 67640 274728 67692 274780
rect 52184 274660 52236 274712
rect 67824 274660 67876 274712
rect 121552 274660 121604 274712
rect 211804 274660 211856 274712
rect 39764 274592 39816 274644
rect 67732 274592 67784 274644
rect 121644 274592 121696 274644
rect 125784 274592 125836 274644
rect 121736 273912 121788 273964
rect 287152 273912 287204 273964
rect 56508 273232 56560 273284
rect 67640 273232 67692 273284
rect 121552 273232 121604 273284
rect 210424 273232 210476 273284
rect 121644 273164 121696 273216
rect 126980 273164 127032 273216
rect 66076 271872 66128 271924
rect 67640 271872 67692 271924
rect 121552 271872 121604 271924
rect 173900 271872 173952 271924
rect 54852 271804 54904 271856
rect 67732 271804 67784 271856
rect 49516 270512 49568 270564
rect 67640 270512 67692 270564
rect 121552 270512 121604 270564
rect 213276 270512 213328 270564
rect 121828 269764 121880 269816
rect 471244 269764 471296 269816
rect 57520 269152 57572 269204
rect 67732 269152 67784 269204
rect 121552 269152 121604 269204
rect 237380 269152 237432 269204
rect 50896 269084 50948 269136
rect 67640 269084 67692 269136
rect 121644 269084 121696 269136
rect 248420 269084 248472 269136
rect 121552 269016 121604 269068
rect 146300 269016 146352 269068
rect 52276 268336 52328 268388
rect 67640 268336 67692 268388
rect 51724 268200 51776 268252
rect 52276 268200 52328 268252
rect 121552 267724 121604 267776
rect 295340 267724 295392 267776
rect 41144 267656 41196 267708
rect 67640 267656 67692 267708
rect 46848 267588 46900 267640
rect 67732 267588 67784 267640
rect 121460 266432 121512 266484
rect 280160 266432 280212 266484
rect 3056 266364 3108 266416
rect 14464 266364 14516 266416
rect 121736 266364 121788 266416
rect 309324 266364 309376 266416
rect 57612 266296 57664 266348
rect 67640 266296 67692 266348
rect 121460 265004 121512 265056
rect 216128 265004 216180 265056
rect 121552 264936 121604 264988
rect 310704 264936 310756 264988
rect 50712 264868 50764 264920
rect 67640 264868 67692 264920
rect 121460 264868 121512 264920
rect 133972 264868 134024 264920
rect 22744 264188 22796 264240
rect 50712 264188 50764 264240
rect 48136 263576 48188 263628
rect 67732 263576 67784 263628
rect 121552 263576 121604 263628
rect 233240 263576 233292 263628
rect 61936 263508 61988 263560
rect 67640 263508 67692 263560
rect 121460 263508 121512 263560
rect 125600 263508 125652 263560
rect 56324 262216 56376 262268
rect 67640 262216 67692 262268
rect 121460 262216 121512 262268
rect 285680 262216 285732 262268
rect 121552 262148 121604 262200
rect 132592 262148 132644 262200
rect 276664 261468 276716 261520
rect 350540 261468 350592 261520
rect 61936 260924 61988 260976
rect 67640 260924 67692 260976
rect 60280 260856 60332 260908
rect 67732 260856 67784 260908
rect 121736 260856 121788 260908
rect 291844 260856 291896 260908
rect 60464 260788 60516 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 131672 260788 131724 260840
rect 131672 260108 131724 260160
rect 353944 260108 353996 260160
rect 53656 259428 53708 259480
rect 67640 259428 67692 259480
rect 121460 259428 121512 259480
rect 207664 259428 207716 259480
rect 125416 259360 125468 259412
rect 579804 259360 579856 259412
rect 121460 259292 121512 259344
rect 127164 259292 127216 259344
rect 65984 258136 66036 258188
rect 67640 258136 67692 258188
rect 58992 258068 59044 258120
rect 67732 258068 67784 258120
rect 121552 258068 121604 258120
rect 288716 258068 288768 258120
rect 34520 258000 34572 258052
rect 35808 258000 35860 258052
rect 67640 258000 67692 258052
rect 15844 257320 15896 257372
rect 34520 257320 34572 257372
rect 233884 257320 233936 257372
rect 296720 257320 296772 257372
rect 63224 256708 63276 256760
rect 67640 256708 67692 256760
rect 121552 256708 121604 256760
rect 242900 256708 242952 256760
rect 121460 256640 121512 256692
rect 128544 256640 128596 256692
rect 54852 255280 54904 255332
rect 67732 255280 67784 255332
rect 59268 255212 59320 255264
rect 67640 255212 67692 255264
rect 125508 254532 125560 254584
rect 580448 254532 580500 254584
rect 121552 254192 121604 254244
rect 123484 254192 123536 254244
rect 3424 253920 3476 253972
rect 17316 253920 17368 253972
rect 60924 253920 60976 253972
rect 67732 253920 67784 253972
rect 121460 253920 121512 253972
rect 236000 253920 236052 253972
rect 42800 253852 42852 253904
rect 43812 253852 43864 253904
rect 67640 253852 67692 253904
rect 35164 253172 35216 253224
rect 42800 253172 42852 253224
rect 63316 252560 63368 252612
rect 67640 252560 67692 252612
rect 121460 252560 121512 252612
rect 282276 252560 282328 252612
rect 121552 251812 121604 251864
rect 231860 251812 231912 251864
rect 121460 251200 121512 251252
rect 276664 251200 276716 251252
rect 57796 249772 57848 249824
rect 67732 249772 67784 249824
rect 121552 249772 121604 249824
rect 206468 249772 206520 249824
rect 39856 249704 39908 249756
rect 67640 249704 67692 249756
rect 121460 249704 121512 249756
rect 131120 249704 131172 249756
rect 67456 248888 67508 248940
rect 68836 248888 68888 248940
rect 121460 248412 121512 248464
rect 310612 248412 310664 248464
rect 130384 247664 130436 247716
rect 580540 247664 580592 247716
rect 65892 247120 65944 247172
rect 67640 247120 67692 247172
rect 59084 247052 59136 247104
rect 67732 247052 67784 247104
rect 121460 247052 121512 247104
rect 218704 247052 218756 247104
rect 54944 246984 54996 247036
rect 67640 246984 67692 247036
rect 121460 245624 121512 245676
rect 237472 245624 237524 245676
rect 57704 245556 57756 245608
rect 67640 245556 67692 245608
rect 64788 244944 64840 244996
rect 68376 244944 68428 244996
rect 61660 244604 61712 244656
rect 66904 244604 66956 244656
rect 67364 244332 67416 244384
rect 68284 244332 68336 244384
rect 63132 244264 63184 244316
rect 67640 244264 67692 244316
rect 121552 244264 121604 244316
rect 306472 244264 306524 244316
rect 321652 244264 321704 244316
rect 580172 244264 580224 244316
rect 49608 244196 49660 244248
rect 67732 244196 67784 244248
rect 121460 244196 121512 244248
rect 125692 244196 125744 244248
rect 66168 242904 66220 242956
rect 67824 242904 67876 242956
rect 121552 242904 121604 242956
rect 275284 242904 275336 242956
rect 62028 242836 62080 242888
rect 67640 242836 67692 242888
rect 121460 242836 121512 242888
rect 142160 242836 142212 242888
rect 321652 242836 321704 242888
rect 121552 242768 121604 242820
rect 129740 242768 129792 242820
rect 122104 241544 122156 241596
rect 209136 241544 209188 241596
rect 60372 241476 60424 241528
rect 67640 241476 67692 241528
rect 121460 241476 121512 241528
rect 232044 241476 232096 241528
rect 3424 240116 3476 240168
rect 61752 240116 61804 240168
rect 67640 240116 67692 240168
rect 119896 240116 119948 240168
rect 288532 240116 288584 240168
rect 37096 240048 37148 240100
rect 118976 239912 119028 239964
rect 119988 239912 120040 239964
rect 70400 239776 70452 239828
rect 71308 239776 71360 239828
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 78680 239776 78732 239828
rect 79680 239776 79732 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 89720 239776 89772 239828
rect 90628 239776 90680 239828
rect 93952 239776 94004 239828
rect 95136 239776 95188 239828
rect 99380 239776 99432 239828
rect 100288 239776 100340 239828
rect 100760 239776 100812 239828
rect 101576 239776 101628 239828
rect 104900 239776 104952 239828
rect 106084 239776 106136 239828
rect 107660 239776 107712 239828
rect 108660 239776 108712 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 65984 239504 66036 239556
rect 254032 239504 254084 239556
rect 63316 239436 63368 239488
rect 272616 239436 272668 239488
rect 63224 239368 63276 239420
rect 299480 239368 299532 239420
rect 84292 239300 84344 239352
rect 85488 239300 85540 239352
rect 50988 238824 51040 238876
rect 82268 238824 82320 238876
rect 103520 238824 103572 238876
rect 115112 238824 115164 238876
rect 132500 238824 132552 238876
rect 37096 238756 37148 238808
rect 106740 238756 106792 238808
rect 139400 238756 139452 238808
rect 52368 238688 52420 238740
rect 98368 238688 98420 238740
rect 118332 238688 118384 238740
rect 123024 238688 123076 238740
rect 59176 238620 59228 238672
rect 91928 238620 91980 238672
rect 53748 238552 53800 238604
rect 95792 238552 95844 238604
rect 113824 238552 113876 238604
rect 128728 238552 128780 238604
rect 60556 238484 60608 238536
rect 72608 238484 72660 238536
rect 99012 238484 99064 238536
rect 124220 238484 124272 238536
rect 89352 238416 89404 238468
rect 133880 238416 133932 238468
rect 105452 238076 105504 238128
rect 184204 238076 184256 238128
rect 96436 238008 96488 238060
rect 276756 238008 276808 238060
rect 102876 237396 102928 237448
rect 105544 237396 105596 237448
rect 48228 237328 48280 237380
rect 107384 237328 107436 237380
rect 110604 237328 110656 237380
rect 136640 237328 136692 237380
rect 14464 237260 14516 237312
rect 117044 237260 117096 237312
rect 127072 237260 127124 237312
rect 57888 237192 57940 237244
rect 86776 237192 86828 237244
rect 60648 237124 60700 237176
rect 117688 237124 117740 237176
rect 110604 236784 110656 236836
rect 111064 236784 111116 236836
rect 69296 236716 69348 236768
rect 230480 236716 230532 236768
rect 282184 236716 282236 236768
rect 331220 236716 331272 236768
rect 64788 236648 64840 236700
rect 306564 236648 306616 236700
rect 17316 235900 17368 235952
rect 34336 235900 34388 235952
rect 112536 235900 112588 235952
rect 114468 235900 114520 235952
rect 124312 235900 124364 235952
rect 91284 235832 91336 235884
rect 140872 235832 140924 235884
rect 117688 235220 117740 235272
rect 177396 235220 177448 235272
rect 45468 234540 45520 234592
rect 109040 234540 109092 234592
rect 81624 234472 81676 234524
rect 135260 234472 135312 234524
rect 109040 234132 109092 234184
rect 109960 234132 110012 234184
rect 74540 233928 74592 233980
rect 75184 233928 75236 233980
rect 122380 233928 122432 233980
rect 313372 233928 313424 233980
rect 66168 233860 66220 233912
rect 276848 233860 276900 233912
rect 83464 233180 83516 233232
rect 143540 233180 143592 233232
rect 92572 232500 92624 232552
rect 238852 232500 238904 232552
rect 84108 231820 84160 231872
rect 84844 231820 84896 231872
rect 94044 231072 94096 231124
rect 271236 231072 271288 231124
rect 76012 230392 76064 230444
rect 128360 230392 128412 230444
rect 128360 229780 128412 229832
rect 187056 229780 187108 229832
rect 97632 229712 97684 229764
rect 303804 229712 303856 229764
rect 78772 226992 78824 227044
rect 231952 226992 232004 227044
rect 82820 226244 82872 226296
rect 133880 226244 133932 226296
rect 135168 226244 135220 226296
rect 135168 224952 135220 225004
rect 358084 224952 358136 225004
rect 71872 224204 71924 224256
rect 268384 224204 268436 224256
rect 61844 222844 61896 222896
rect 244280 222844 244332 222896
rect 53564 220124 53616 220176
rect 142804 220124 142856 220176
rect 103612 220056 103664 220108
rect 287244 220056 287296 220108
rect 60372 218696 60424 218748
rect 247040 218696 247092 218748
rect 74632 217336 74684 217388
rect 265624 217336 265676 217388
rect 57520 217268 57572 217320
rect 252560 217268 252612 217320
rect 231124 216044 231176 216096
rect 245660 216044 245712 216096
rect 88340 215976 88392 216028
rect 285956 215976 286008 216028
rect 73252 215908 73304 215960
rect 273996 215908 274048 215960
rect 3332 215228 3384 215280
rect 22744 215228 22796 215280
rect 50896 214548 50948 214600
rect 295432 214548 295484 214600
rect 61752 213256 61804 213308
rect 261484 213256 261536 213308
rect 48136 213188 48188 213240
rect 305092 213188 305144 213240
rect 123484 211828 123536 211880
rect 255964 211828 256016 211880
rect 77392 211760 77444 211812
rect 233332 211760 233384 211812
rect 46756 210400 46808 210452
rect 302424 210400 302476 210452
rect 89812 209040 89864 209092
rect 233424 209040 233476 209092
rect 55036 207748 55088 207800
rect 213368 207748 213420 207800
rect 104900 207680 104952 207732
rect 284392 207680 284444 207732
rect 56324 207612 56376 207664
rect 241520 207612 241572 207664
rect 100852 206388 100904 206440
rect 232136 206388 232188 206440
rect 69112 206320 69164 206372
rect 230572 206320 230624 206372
rect 102140 206252 102192 206304
rect 289912 206252 289964 206304
rect 163504 205028 163556 205080
rect 264336 205028 264388 205080
rect 105544 204960 105596 205012
rect 220176 204960 220228 205012
rect 52092 204892 52144 204944
rect 269948 204892 270000 204944
rect 93952 203600 94004 203652
rect 258816 203600 258868 203652
rect 14464 203532 14516 203584
rect 83464 203532 83516 203584
rect 113180 203532 113232 203584
rect 306656 203532 306708 203584
rect 3424 202784 3476 202836
rect 120080 202784 120132 202836
rect 100760 202172 100812 202224
rect 234804 202172 234856 202224
rect 151084 202104 151136 202156
rect 305184 202104 305236 202156
rect 133144 200812 133196 200864
rect 240232 200812 240284 200864
rect 152464 200744 152516 200796
rect 303896 200744 303948 200796
rect 96620 199656 96672 199708
rect 218796 199656 218848 199708
rect 166356 199588 166408 199640
rect 291200 199588 291252 199640
rect 93860 199520 93912 199572
rect 234896 199520 234948 199572
rect 280804 199520 280856 199572
rect 300952 199520 301004 199572
rect 107752 199452 107804 199504
rect 299664 199452 299716 199504
rect 52184 199384 52236 199436
rect 296904 199384 296956 199436
rect 157984 198024 158036 198076
rect 294052 198024 294104 198076
rect 73160 197956 73212 198008
rect 275376 197956 275428 198008
rect 67548 196732 67600 196784
rect 230664 196732 230716 196784
rect 92480 196664 92532 196716
rect 285864 196664 285916 196716
rect 86224 196596 86276 196648
rect 582564 196596 582616 196648
rect 84292 195372 84344 195424
rect 233516 195372 233568 195424
rect 107660 195304 107712 195356
rect 285772 195304 285824 195356
rect 70492 195236 70544 195288
rect 276940 195236 276992 195288
rect 145564 194080 145616 194132
rect 196716 194080 196768 194132
rect 110420 194012 110472 194064
rect 236092 194012 236144 194064
rect 50804 193944 50856 193996
rect 244372 193944 244424 193996
rect 56508 193876 56560 193928
rect 260840 193876 260892 193928
rect 54852 193808 54904 193860
rect 296996 193808 297048 193860
rect 352564 193128 352616 193180
rect 580172 193128 580224 193180
rect 142804 192516 142856 192568
rect 242992 192516 243044 192568
rect 61936 192448 61988 192500
rect 294144 192448 294196 192500
rect 103520 191292 103572 191344
rect 180248 191292 180300 191344
rect 111800 191224 111852 191276
rect 251364 191224 251416 191276
rect 114560 191156 114612 191208
rect 280252 191156 280304 191208
rect 70400 191088 70452 191140
rect 247132 191088 247184 191140
rect 214656 189728 214708 189780
rect 292764 189728 292816 189780
rect 105544 189048 105596 189100
rect 214748 189048 214800 189100
rect 3424 188980 3476 189032
rect 17224 188980 17276 189032
rect 192484 188436 192536 188488
rect 302516 188436 302568 188488
rect 89720 188368 89772 188420
rect 241612 188368 241664 188420
rect 99380 188300 99432 188352
rect 252652 188300 252704 188352
rect 101956 187756 102008 187808
rect 171876 187756 171928 187808
rect 104808 187688 104860 187740
rect 184296 187688 184348 187740
rect 224316 187008 224368 187060
rect 298284 187008 298336 187060
rect 155224 186940 155276 186992
rect 295524 186940 295576 186992
rect 128268 186396 128320 186448
rect 171968 186396 172020 186448
rect 99288 186328 99340 186380
rect 214656 186328 214708 186380
rect 40684 185784 40736 185836
rect 109040 185784 109092 185836
rect 61660 185716 61712 185768
rect 244556 185716 244608 185768
rect 58992 185648 59044 185700
rect 249800 185648 249852 185700
rect 282276 185648 282328 185700
rect 308036 185648 308088 185700
rect 84200 185580 84252 185632
rect 283012 185580 283064 185632
rect 119988 184968 120040 185020
rect 170496 184968 170548 185020
rect 114468 184900 114520 184952
rect 213460 184900 213512 184952
rect 115940 184288 115992 184340
rect 248604 184288 248656 184340
rect 271236 184288 271288 184340
rect 299572 184288 299624 184340
rect 80152 184220 80204 184272
rect 284484 184220 284536 184272
rect 69020 184152 69072 184204
rect 281540 184152 281592 184204
rect 100668 183540 100720 183592
rect 167644 183540 167696 183592
rect 159364 183064 159416 183116
rect 198096 183064 198148 183116
rect 180156 182996 180208 183048
rect 227720 182996 227772 183048
rect 65892 182928 65944 182980
rect 251272 182928 251324 182980
rect 59084 182860 59136 182912
rect 245844 182860 245896 182912
rect 80060 182792 80112 182844
rect 280436 182792 280488 182844
rect 264336 182724 264388 182776
rect 269120 182724 269172 182776
rect 118424 182248 118476 182300
rect 166356 182248 166408 182300
rect 97724 182180 97776 182232
rect 169116 182180 169168 182232
rect 278136 181772 278188 181824
rect 301044 181772 301096 181824
rect 213276 181704 213328 181756
rect 240140 181704 240192 181756
rect 261484 181704 261536 181756
rect 292580 181704 292632 181756
rect 198188 181636 198240 181688
rect 256792 181636 256844 181688
rect 269764 181636 269816 181688
rect 307760 181636 307812 181688
rect 86960 181568 87012 181620
rect 236184 181568 236236 181620
rect 264244 181568 264296 181620
rect 335360 181568 335412 181620
rect 53656 181500 53708 181552
rect 291476 181500 291528 181552
rect 60280 181432 60332 181484
rect 301136 181432 301188 181484
rect 129464 180956 129516 181008
rect 166448 180956 166500 181008
rect 122656 180888 122708 180940
rect 167920 180888 167972 180940
rect 114100 180820 114152 180872
rect 169208 180820 169260 180872
rect 226984 180412 227036 180464
rect 248512 180412 248564 180464
rect 213368 180344 213420 180396
rect 241704 180344 241756 180396
rect 166264 180276 166316 180328
rect 199476 180276 199528 180328
rect 204996 180276 205048 180328
rect 238760 180276 238812 180328
rect 273904 180276 273956 180328
rect 288440 180276 288492 180328
rect 162124 180208 162176 180260
rect 206376 180208 206428 180260
rect 207664 180208 207716 180260
rect 258080 180208 258132 180260
rect 271144 180208 271196 180260
rect 299756 180208 299808 180260
rect 182824 180140 182876 180192
rect 244464 180140 244516 180192
rect 258816 180140 258868 180192
rect 296812 180140 296864 180192
rect 69204 180072 69256 180124
rect 280344 180072 280396 180124
rect 133144 179460 133196 179512
rect 165068 179460 165120 179512
rect 126796 179392 126848 179444
rect 166540 179392 166592 179444
rect 272524 179324 272576 179376
rect 279332 179324 279384 179376
rect 211804 178984 211856 179036
rect 245752 178984 245804 179036
rect 203524 178916 203576 178968
rect 243084 178916 243136 178968
rect 178776 178848 178828 178900
rect 238944 178848 238996 178900
rect 169024 178780 169076 178832
rect 240324 178780 240376 178832
rect 269856 178780 269908 178832
rect 278780 178780 278832 178832
rect 220084 178712 220136 178764
rect 299388 178712 299440 178764
rect 214564 178644 214616 178696
rect 340972 178644 341024 178696
rect 134800 178372 134852 178424
rect 165528 178372 165580 178424
rect 132408 178304 132460 178356
rect 165436 178304 165488 178356
rect 123760 178236 123812 178288
rect 169300 178236 169352 178288
rect 115848 178168 115900 178220
rect 167828 178168 167880 178220
rect 148232 178100 148284 178152
rect 210516 178100 210568 178152
rect 130752 178032 130804 178084
rect 214104 178032 214156 178084
rect 298744 178032 298796 178084
rect 299480 178032 299532 178084
rect 222844 177964 222896 178016
rect 229376 177964 229428 178016
rect 102048 177828 102100 177880
rect 105544 177828 105596 177880
rect 276756 177624 276808 177676
rect 287060 177624 287112 177676
rect 276940 177556 276992 177608
rect 288624 177556 288676 177608
rect 221464 177488 221516 177540
rect 229100 177488 229152 177540
rect 272616 177488 272668 177540
rect 284300 177488 284352 177540
rect 220176 177420 220228 177472
rect 237656 177420 237708 177472
rect 276664 177420 276716 177472
rect 291384 177420 291436 177472
rect 218796 177352 218848 177404
rect 237564 177352 237616 177404
rect 268384 177352 268436 177404
rect 292672 177352 292724 177404
rect 227168 177284 227220 177336
rect 247224 177284 247276 177336
rect 255964 177284 256016 177336
rect 290096 177284 290148 177336
rect 291844 177148 291896 177200
rect 295616 177148 295668 177200
rect 128176 177012 128228 177064
rect 169760 177012 169812 177064
rect 107016 176944 107068 176996
rect 164424 176944 164476 176996
rect 105728 176876 105780 176928
rect 169024 176876 169076 176928
rect 103336 176808 103388 176860
rect 167736 176808 167788 176860
rect 136088 176740 136140 176792
rect 213828 176740 213880 176792
rect 108120 176672 108172 176724
rect 188436 176672 188488 176724
rect 158904 176264 158956 176316
rect 166264 176264 166316 176316
rect 164424 176196 164476 176248
rect 214564 176196 214616 176248
rect 110696 176128 110748 176180
rect 170588 176128 170640 176180
rect 210424 176128 210476 176180
rect 229192 176128 229244 176180
rect 275376 176128 275428 176180
rect 281632 176128 281684 176180
rect 124496 176060 124548 176112
rect 211804 176060 211856 176112
rect 218704 176060 218756 176112
rect 229284 176060 229336 176112
rect 276848 176060 276900 176112
rect 289820 176060 289872 176112
rect 120816 175992 120868 176044
rect 210608 175992 210660 176044
rect 225604 175992 225656 176044
rect 243176 175992 243228 176044
rect 273996 175992 274048 176044
rect 290004 175992 290056 176044
rect 290464 175992 290516 176044
rect 292856 175992 292908 176044
rect 11704 175924 11756 175976
rect 111064 175924 111116 175976
rect 116952 175924 117004 175976
rect 213276 175924 213328 175976
rect 224224 175924 224276 175976
rect 251456 175924 251508 175976
rect 275284 175924 275336 175976
rect 294236 175924 294288 175976
rect 165068 175176 165120 175228
rect 214012 175176 214064 175228
rect 236644 175176 236696 175228
rect 237380 175176 237432 175228
rect 165528 175108 165580 175160
rect 213920 175108 213972 175160
rect 254584 173952 254636 174004
rect 265808 173952 265860 174004
rect 242532 173884 242584 173936
rect 264428 173884 264480 173936
rect 165436 173816 165488 173868
rect 213920 173816 213972 173868
rect 231768 173816 231820 173868
rect 242992 173816 243044 173868
rect 231124 173748 231176 173800
rect 240232 173748 240284 173800
rect 231492 173680 231544 173732
rect 238760 173680 238812 173732
rect 243728 173136 243780 173188
rect 265716 173136 265768 173188
rect 262864 172592 262916 172644
rect 265532 172592 265584 172644
rect 238116 172524 238168 172576
rect 265900 172524 265952 172576
rect 166448 172456 166500 172508
rect 213920 172456 213972 172508
rect 231768 172456 231820 172508
rect 240140 172456 240192 172508
rect 169760 172388 169812 172440
rect 214012 172388 214064 172440
rect 282092 171776 282144 171828
rect 287060 171776 287112 171828
rect 167552 171300 167604 171352
rect 170680 171300 170732 171352
rect 257344 171232 257396 171284
rect 265624 171232 265676 171284
rect 246396 171164 246448 171216
rect 265808 171164 265860 171216
rect 241152 171096 241204 171148
rect 265900 171096 265952 171148
rect 166540 171028 166592 171080
rect 214012 171028 214064 171080
rect 231768 171028 231820 171080
rect 245660 171028 245712 171080
rect 171968 170960 172020 171012
rect 215116 170960 215168 171012
rect 231124 170960 231176 171012
rect 245844 170960 245896 171012
rect 231492 170892 231544 170944
rect 244280 170892 244332 170944
rect 229744 170416 229796 170468
rect 239036 170416 239088 170468
rect 229836 170348 229888 170400
rect 241612 170348 241664 170400
rect 258908 169872 258960 169924
rect 265256 169872 265308 169924
rect 282276 169872 282328 169924
rect 288440 169872 288492 169924
rect 244924 169804 244976 169856
rect 265440 169804 265492 169856
rect 239680 169736 239732 169788
rect 265624 169736 265676 169788
rect 281724 169736 281776 169788
rect 284300 169736 284352 169788
rect 169300 169668 169352 169720
rect 213920 169668 213972 169720
rect 231492 169668 231544 169720
rect 237564 169668 237616 169720
rect 282828 169668 282880 169720
rect 301136 169668 301188 169720
rect 211804 169600 211856 169652
rect 214012 169600 214064 169652
rect 230756 169532 230808 169584
rect 237656 169532 237708 169584
rect 256240 168512 256292 168564
rect 265348 168512 265400 168564
rect 242440 168444 242492 168496
rect 265808 168444 265860 168496
rect 239772 168376 239824 168428
rect 265624 168376 265676 168428
rect 167920 168308 167972 168360
rect 213920 168308 213972 168360
rect 231768 168308 231820 168360
rect 238944 168308 238996 168360
rect 282460 168308 282512 168360
rect 289820 168308 289872 168360
rect 210608 168240 210660 168292
rect 214012 168240 214064 168292
rect 232504 167628 232556 167680
rect 243084 167628 243136 167680
rect 250536 167084 250588 167136
rect 265348 167084 265400 167136
rect 243636 167016 243688 167068
rect 264428 167016 264480 167068
rect 231676 166948 231728 167000
rect 241520 166948 241572 167000
rect 282092 166948 282144 167000
rect 295432 166948 295484 167000
rect 353944 166948 353996 167000
rect 580172 166948 580224 167000
rect 170496 166880 170548 166932
rect 213920 166880 213972 166932
rect 231768 166880 231820 166932
rect 238852 166880 238904 166932
rect 166356 166812 166408 166864
rect 214012 166812 214064 166864
rect 282644 166268 282696 166320
rect 294144 166268 294196 166320
rect 253480 165724 253532 165776
rect 265808 165724 265860 165776
rect 246304 165656 246356 165708
rect 265716 165656 265768 165708
rect 238300 165588 238352 165640
rect 265348 165588 265400 165640
rect 167828 165520 167880 165572
rect 213920 165520 213972 165572
rect 231124 165520 231176 165572
rect 233424 165520 233476 165572
rect 282092 165520 282144 165572
rect 289912 165520 289964 165572
rect 231676 165452 231728 165504
rect 241704 165452 241756 165504
rect 231768 165384 231820 165436
rect 243176 165384 243228 165436
rect 249064 164840 249116 164892
rect 265256 164840 265308 164892
rect 255964 164296 256016 164348
rect 265164 164296 265216 164348
rect 240784 164228 240836 164280
rect 265348 164228 265400 164280
rect 3240 164160 3292 164212
rect 25504 164160 25556 164212
rect 169208 164160 169260 164212
rect 213920 164160 213972 164212
rect 231124 164160 231176 164212
rect 233240 164160 233292 164212
rect 282828 164160 282880 164212
rect 291476 164160 291528 164212
rect 231768 164092 231820 164144
rect 240416 164092 240468 164144
rect 231676 164024 231728 164076
rect 244556 164024 244608 164076
rect 242164 163480 242216 163532
rect 265164 163480 265216 163532
rect 234068 163004 234120 163056
rect 265808 163004 265860 163056
rect 258724 162868 258776 162920
rect 265532 162868 265584 162920
rect 282736 162868 282788 162920
rect 288624 162868 288676 162920
rect 170588 162800 170640 162852
rect 213920 162800 213972 162852
rect 231032 162800 231084 162852
rect 233332 162800 233384 162852
rect 282552 162800 282604 162852
rect 294236 162800 294288 162852
rect 282828 162732 282880 162784
rect 292856 162732 292908 162784
rect 231676 162664 231728 162716
rect 244372 162664 244424 162716
rect 231768 162460 231820 162512
rect 236644 162460 236696 162512
rect 233884 162120 233936 162172
rect 247132 162120 247184 162172
rect 253388 161576 253440 161628
rect 264428 161576 264480 161628
rect 247684 161508 247736 161560
rect 265532 161508 265584 161560
rect 241060 161440 241112 161492
rect 264520 161440 264572 161492
rect 188436 161372 188488 161424
rect 213920 161372 213972 161424
rect 231676 161372 231728 161424
rect 248604 161372 248656 161424
rect 282828 161372 282880 161424
rect 302332 161372 302384 161424
rect 231768 161304 231820 161356
rect 238760 161304 238812 161356
rect 282368 161304 282420 161356
rect 292764 161304 292816 161356
rect 167736 160692 167788 160744
rect 214104 160692 214156 160744
rect 247868 160216 247920 160268
rect 265900 160216 265952 160268
rect 245016 160148 245068 160200
rect 265808 160148 265860 160200
rect 242348 160080 242400 160132
rect 265992 160080 266044 160132
rect 169024 160012 169076 160064
rect 213920 160012 213972 160064
rect 231768 160012 231820 160064
rect 247224 160012 247276 160064
rect 184296 159944 184348 159996
rect 214012 159944 214064 159996
rect 231676 159944 231728 159996
rect 240324 159944 240376 159996
rect 231676 159468 231728 159520
rect 234712 159468 234764 159520
rect 261760 158788 261812 158840
rect 265440 158788 265492 158840
rect 246580 158720 246632 158772
rect 265532 158720 265584 158772
rect 282276 158652 282328 158704
rect 299756 158652 299808 158704
rect 170680 157972 170732 158024
rect 214932 157972 214984 158024
rect 256148 157972 256200 158024
rect 265808 157972 265860 158024
rect 245108 157428 245160 157480
rect 265808 157428 265860 157480
rect 237380 157360 237432 157412
rect 265992 157360 266044 157412
rect 167644 157292 167696 157344
rect 214012 157292 214064 157344
rect 231676 157292 231728 157344
rect 258080 157292 258132 157344
rect 282828 157292 282880 157344
rect 301044 157292 301096 157344
rect 171876 157224 171928 157276
rect 213920 157224 213972 157276
rect 231768 157224 231820 157276
rect 244464 157224 244516 157276
rect 239588 156612 239640 156664
rect 265072 156612 265124 156664
rect 232780 156136 232832 156188
rect 237472 156136 237524 156188
rect 250444 156000 250496 156052
rect 265900 156000 265952 156052
rect 238024 155932 238076 155984
rect 265808 155932 265860 155984
rect 169116 155864 169168 155916
rect 213920 155864 213972 155916
rect 230940 155864 230992 155916
rect 233516 155864 233568 155916
rect 282828 155864 282880 155916
rect 302516 155864 302568 155916
rect 230572 155796 230624 155848
rect 232136 155796 232188 155848
rect 263140 154708 263192 154760
rect 265808 154708 265860 154760
rect 240968 154640 241020 154692
rect 265992 154640 266044 154692
rect 233976 154572 234028 154624
rect 265716 154572 265768 154624
rect 231400 154504 231452 154556
rect 252560 154504 252612 154556
rect 231768 154300 231820 154352
rect 236184 154300 236236 154352
rect 281908 154164 281960 154216
rect 285956 154164 286008 154216
rect 231124 154096 231176 154148
rect 237380 154096 237432 154148
rect 239404 153824 239456 153876
rect 265900 153824 265952 153876
rect 231308 153348 231360 153400
rect 233884 153348 233936 153400
rect 196808 153280 196860 153332
rect 213920 153280 213972 153332
rect 258816 153280 258868 153332
rect 265808 153280 265860 153332
rect 281724 153280 281776 153332
rect 284484 153280 284536 153332
rect 167644 153212 167696 153264
rect 214012 153212 214064 153264
rect 238208 153212 238260 153264
rect 265348 153212 265400 153264
rect 230756 153144 230808 153196
rect 255320 153144 255372 153196
rect 282184 153144 282236 153196
rect 308036 153144 308088 153196
rect 468484 153144 468536 153196
rect 579804 153144 579856 153196
rect 231768 153076 231820 153128
rect 245752 153076 245804 153128
rect 231676 152668 231728 152720
rect 234620 152668 234672 152720
rect 211804 152396 211856 152448
rect 213920 152396 213972 152448
rect 235448 151920 235500 151972
rect 265256 151920 265308 151972
rect 253204 151852 253256 151904
rect 265808 151852 265860 151904
rect 171784 151784 171836 151836
rect 213920 151784 213972 151836
rect 231676 151716 231728 151768
rect 252652 151716 252704 151768
rect 282828 151716 282880 151768
rect 299664 151716 299716 151768
rect 231768 151648 231820 151700
rect 251364 151648 251416 151700
rect 282000 151648 282052 151700
rect 290004 151648 290056 151700
rect 260472 150560 260524 150612
rect 265716 150560 265768 150612
rect 245200 150492 245252 150544
rect 265808 150492 265860 150544
rect 173348 150424 173400 150476
rect 213920 150424 213972 150476
rect 236828 150424 236880 150476
rect 265440 150424 265492 150476
rect 3424 150356 3476 150408
rect 32404 150356 32456 150408
rect 210516 150356 210568 150408
rect 214012 150356 214064 150408
rect 230940 150356 230992 150408
rect 256792 150356 256844 150408
rect 282828 150356 282880 150408
rect 296904 150356 296956 150408
rect 231032 150288 231084 150340
rect 234896 150288 234948 150340
rect 282184 150288 282236 150340
rect 291384 150288 291436 150340
rect 231216 149744 231268 149796
rect 250444 149744 250496 149796
rect 236920 149676 236972 149728
rect 265900 149676 265952 149728
rect 231308 149472 231360 149524
rect 236000 149472 236052 149524
rect 259092 149132 259144 149184
rect 265348 149132 265400 149184
rect 250720 149064 250772 149116
rect 265808 149064 265860 149116
rect 166264 148996 166316 149048
rect 213920 148996 213972 149048
rect 231768 148996 231820 149048
rect 251456 148996 251508 149048
rect 282092 148928 282144 148980
rect 309324 148928 309376 148980
rect 257528 148316 257580 148368
rect 265440 148316 265492 148368
rect 235540 147704 235592 147756
rect 265716 147704 265768 147756
rect 187148 147636 187200 147688
rect 213920 147636 213972 147688
rect 233884 147636 233936 147688
rect 265532 147636 265584 147688
rect 230940 147568 230992 147620
rect 234804 147568 234856 147620
rect 281724 147568 281776 147620
rect 305184 147568 305236 147620
rect 230756 147500 230808 147552
rect 232504 147500 232556 147552
rect 231400 146956 231452 147008
rect 242532 146956 242584 147008
rect 242256 146888 242308 146940
rect 265072 146888 265124 146940
rect 261576 146344 261628 146396
rect 265900 146344 265952 146396
rect 171876 146276 171928 146328
rect 213920 146276 213972 146328
rect 235632 146276 235684 146328
rect 265532 146276 265584 146328
rect 231768 146208 231820 146260
rect 249800 146208 249852 146260
rect 282828 146208 282880 146260
rect 307944 146208 307996 146260
rect 231676 146140 231728 146192
rect 247040 146140 247092 146192
rect 282736 146140 282788 146192
rect 296996 146140 297048 146192
rect 254768 145052 254820 145104
rect 265900 145052 265952 145104
rect 243820 144984 243872 145036
rect 265716 144984 265768 145036
rect 189816 144916 189868 144968
rect 213920 144916 213972 144968
rect 234160 144916 234212 144968
rect 265808 144916 265860 144968
rect 231768 144848 231820 144900
rect 248420 144848 248472 144900
rect 282828 144848 282880 144900
rect 298192 144848 298244 144900
rect 174636 144168 174688 144220
rect 214656 144168 214708 144220
rect 230756 144168 230808 144220
rect 232688 144168 232740 144220
rect 232596 144100 232648 144152
rect 265992 144168 266044 144220
rect 282828 143692 282880 143744
rect 287152 143692 287204 143744
rect 182824 143556 182876 143608
rect 213920 143556 213972 143608
rect 262956 143556 263008 143608
rect 265532 143556 265584 143608
rect 231768 143488 231820 143540
rect 242900 143488 242952 143540
rect 282092 143488 282144 143540
rect 306564 143488 306616 143540
rect 230480 143420 230532 143472
rect 232780 143420 232832 143472
rect 282276 143420 282328 143472
rect 298284 143420 298336 143472
rect 282184 142944 282236 142996
rect 285680 142944 285732 142996
rect 167736 142808 167788 142860
rect 214012 142808 214064 142860
rect 232688 142808 232740 142860
rect 265808 142808 265860 142860
rect 195428 142196 195480 142248
rect 213920 142196 213972 142248
rect 184296 142128 184348 142180
rect 214012 142128 214064 142180
rect 252100 142128 252152 142180
rect 265348 142128 265400 142180
rect 282828 142060 282880 142112
rect 310704 142060 310756 142112
rect 282736 141992 282788 142044
rect 295524 141992 295576 142044
rect 176016 140836 176068 140888
rect 213920 140836 213972 140888
rect 250812 140836 250864 140888
rect 265532 140836 265584 140888
rect 169024 140768 169076 140820
rect 214012 140768 214064 140820
rect 232780 140768 232832 140820
rect 264428 140768 264480 140820
rect 231492 140700 231544 140752
rect 262220 140700 262272 140752
rect 282828 140700 282880 140752
rect 287336 140700 287388 140752
rect 231768 140632 231820 140684
rect 260840 140632 260892 140684
rect 230940 140564 230992 140616
rect 248512 140564 248564 140616
rect 169116 140020 169168 140072
rect 214472 140020 214524 140072
rect 253572 140020 253624 140072
rect 265808 140020 265860 140072
rect 236736 139476 236788 139528
rect 265808 139476 265860 139528
rect 170588 139408 170640 139460
rect 213920 139408 213972 139460
rect 230020 139408 230072 139460
rect 265716 139408 265768 139460
rect 231768 139340 231820 139392
rect 251272 139340 251324 139392
rect 282828 139340 282880 139392
rect 307852 139340 307904 139392
rect 282736 139272 282788 139324
rect 305276 139272 305328 139324
rect 231676 139204 231728 139256
rect 236092 139204 236144 139256
rect 181444 138660 181496 138712
rect 214012 138660 214064 138712
rect 231032 138660 231084 138712
rect 241152 138660 241204 138712
rect 251916 138048 251968 138100
rect 265164 138048 265216 138100
rect 170496 137980 170548 138032
rect 213920 137980 213972 138032
rect 240876 137980 240928 138032
rect 265808 137980 265860 138032
rect 3240 137912 3292 137964
rect 15844 137912 15896 137964
rect 231492 137912 231544 137964
rect 259460 137912 259512 137964
rect 282828 137912 282880 137964
rect 295616 137912 295668 137964
rect 231768 137844 231820 137896
rect 256700 137844 256752 137896
rect 249340 137232 249392 137284
rect 265256 137232 265308 137284
rect 236644 136688 236696 136740
rect 265716 136688 265768 136740
rect 192576 136620 192628 136672
rect 213920 136620 213972 136672
rect 229928 136620 229980 136672
rect 265808 136620 265860 136672
rect 231768 136552 231820 136604
rect 254032 136552 254084 136604
rect 282736 136552 282788 136604
rect 309232 136552 309284 136604
rect 231676 136484 231728 136536
rect 243728 136484 243780 136536
rect 282828 136484 282880 136536
rect 292672 136484 292724 136536
rect 260196 135396 260248 135448
rect 265164 135396 265216 135448
rect 203616 135328 203668 135380
rect 214012 135328 214064 135380
rect 243544 135328 243596 135380
rect 265808 135328 265860 135380
rect 185676 135260 185728 135312
rect 213920 135260 213972 135312
rect 229744 135260 229796 135312
rect 265992 135260 266044 135312
rect 231768 135192 231820 135244
rect 261484 135192 261536 135244
rect 282736 135192 282788 135244
rect 310520 135192 310572 135244
rect 231676 135124 231728 135176
rect 254584 135124 254636 135176
rect 282828 135124 282880 135176
rect 294052 135124 294104 135176
rect 230756 134172 230808 134224
rect 238116 134172 238168 134224
rect 261668 134036 261720 134088
rect 265808 134036 265860 134088
rect 177488 133968 177540 134020
rect 214012 133968 214064 134020
rect 262956 133968 263008 134020
rect 265256 133968 265308 134020
rect 173164 133900 173216 133952
rect 213920 133900 213972 133952
rect 254676 133900 254728 133952
rect 264428 133900 264480 133952
rect 231768 133832 231820 133884
rect 262864 133832 262916 133884
rect 281908 133832 281960 133884
rect 313372 133832 313424 133884
rect 231676 133764 231728 133816
rect 261760 133764 261812 133816
rect 263048 132608 263100 132660
rect 265624 132608 265676 132660
rect 230756 132404 230808 132456
rect 257344 132404 257396 132456
rect 231492 132336 231544 132388
rect 246396 132336 246448 132388
rect 282828 132336 282880 132388
rect 303896 132336 303948 132388
rect 231768 132268 231820 132320
rect 244924 132268 244976 132320
rect 246672 131724 246724 131776
rect 265532 131724 265584 131776
rect 191196 131180 191248 131232
rect 214012 131180 214064 131232
rect 175924 131112 175976 131164
rect 213920 131112 213972 131164
rect 246488 131112 246540 131164
rect 265716 131112 265768 131164
rect 231768 131044 231820 131096
rect 258908 131044 258960 131096
rect 231400 130976 231452 131028
rect 242440 130976 242492 131028
rect 231492 130908 231544 130960
rect 239680 130908 239732 130960
rect 282276 130432 282328 130484
rect 288716 130432 288768 130484
rect 281724 130092 281776 130144
rect 285864 130092 285916 130144
rect 257436 129820 257488 129872
rect 261300 129820 261352 129872
rect 174544 129752 174596 129804
rect 213920 129752 213972 129804
rect 239496 129752 239548 129804
rect 264428 129752 264480 129804
rect 231768 129684 231820 129736
rect 256240 129684 256292 129736
rect 231676 129616 231728 129668
rect 239772 129616 239824 129668
rect 282828 129208 282880 129260
rect 288532 129208 288584 129260
rect 256056 128460 256108 128512
rect 264428 128460 264480 128512
rect 247776 128392 247828 128444
rect 265808 128392 265860 128444
rect 171968 128324 172020 128376
rect 213920 128324 213972 128376
rect 235356 128324 235408 128376
rect 265348 128324 265400 128376
rect 230756 128256 230808 128308
rect 250536 128256 250588 128308
rect 231768 128188 231820 128240
rect 249064 128188 249116 128240
rect 231676 128120 231728 128172
rect 243636 128120 243688 128172
rect 281908 127916 281960 127968
rect 285772 127916 285824 127968
rect 250444 127032 250496 127084
rect 265348 127032 265400 127084
rect 192484 126964 192536 127016
rect 213920 126964 213972 127016
rect 249156 126964 249208 127016
rect 264428 126964 264480 127016
rect 231768 126896 231820 126948
rect 246304 126896 246356 126948
rect 282828 126896 282880 126948
rect 302240 126896 302292 126948
rect 467104 126896 467156 126948
rect 580172 126896 580224 126948
rect 231584 125808 231636 125860
rect 234068 125808 234120 125860
rect 256240 125740 256292 125792
rect 265716 125740 265768 125792
rect 180340 125672 180392 125724
rect 214012 125672 214064 125724
rect 253296 125672 253348 125724
rect 265808 125672 265860 125724
rect 166264 125604 166316 125656
rect 213920 125604 213972 125656
rect 238116 125604 238168 125656
rect 265624 125604 265676 125656
rect 231492 125536 231544 125588
rect 255964 125536 256016 125588
rect 282736 125536 282788 125588
rect 303712 125536 303764 125588
rect 231768 125468 231820 125520
rect 240784 125468 240836 125520
rect 282828 125468 282880 125520
rect 290096 125468 290148 125520
rect 230664 124856 230716 124908
rect 246580 124856 246632 124908
rect 261484 124312 261536 124364
rect 265532 124312 265584 124364
rect 200764 124244 200816 124296
rect 213920 124244 213972 124296
rect 251824 124244 251876 124296
rect 265808 124244 265860 124296
rect 60648 124176 60700 124228
rect 65524 124176 65576 124228
rect 170680 124176 170732 124228
rect 214012 124176 214064 124228
rect 244924 124176 244976 124228
rect 265900 124176 265952 124228
rect 231768 124108 231820 124160
rect 242164 124108 242216 124160
rect 282000 123972 282052 124024
rect 284576 123972 284628 124024
rect 170404 123428 170456 123480
rect 202236 123428 202288 123480
rect 231400 123428 231452 123480
rect 263140 123428 263192 123480
rect 260104 122952 260156 123004
rect 264428 122952 264480 123004
rect 173256 122884 173308 122936
rect 214012 122884 214064 122936
rect 262864 122884 262916 122936
rect 265808 122884 265860 122936
rect 62028 122816 62080 122868
rect 66076 122816 66128 122868
rect 167828 122816 167880 122868
rect 213920 122816 213972 122868
rect 232504 122816 232556 122868
rect 265900 122816 265952 122868
rect 230940 122748 230992 122800
rect 258724 122748 258776 122800
rect 282092 122748 282144 122800
rect 305000 122748 305052 122800
rect 231768 122680 231820 122732
rect 246672 122680 246724 122732
rect 282828 122680 282880 122732
rect 291292 122680 291344 122732
rect 231492 122612 231544 122664
rect 241060 122612 241112 122664
rect 258908 121592 258960 121644
rect 264428 121592 264480 121644
rect 184388 121524 184440 121576
rect 214012 121524 214064 121576
rect 257344 121524 257396 121576
rect 265900 121524 265952 121576
rect 177580 121456 177632 121508
rect 213920 121456 213972 121508
rect 240784 121456 240836 121508
rect 265808 121456 265860 121508
rect 231768 121388 231820 121440
rect 253388 121388 253440 121440
rect 282736 121388 282788 121440
rect 300952 121388 301004 121440
rect 231308 121320 231360 121372
rect 247684 121320 247736 121372
rect 282828 121320 282880 121372
rect 299572 121320 299624 121372
rect 231492 121252 231544 121304
rect 242348 121252 242400 121304
rect 254584 120232 254636 120284
rect 265808 120232 265860 120284
rect 178776 120164 178828 120216
rect 214012 120164 214064 120216
rect 249064 120164 249116 120216
rect 265900 120164 265952 120216
rect 173440 120096 173492 120148
rect 213920 120096 213972 120148
rect 242440 120096 242492 120148
rect 265992 120096 266044 120148
rect 231768 120028 231820 120080
rect 247868 120028 247920 120080
rect 282828 120028 282880 120080
rect 306472 120028 306524 120080
rect 231308 119960 231360 120012
rect 245016 119960 245068 120012
rect 177304 119348 177356 119400
rect 195336 119348 195388 119400
rect 238392 119348 238444 119400
rect 265532 119348 265584 119400
rect 177672 118804 177724 118856
rect 213920 118804 213972 118856
rect 246304 118804 246356 118856
rect 265532 118804 265584 118856
rect 209228 118736 209280 118788
rect 214012 118736 214064 118788
rect 247684 118736 247736 118788
rect 265624 118736 265676 118788
rect 231400 118600 231452 118652
rect 256148 118600 256200 118652
rect 282828 118600 282880 118652
rect 296812 118600 296864 118652
rect 281908 118532 281960 118584
rect 284392 118532 284444 118584
rect 231400 117784 231452 117836
rect 235632 117784 235684 117836
rect 255964 117444 256016 117496
rect 265992 117444 266044 117496
rect 210424 117376 210476 117428
rect 214012 117376 214064 117428
rect 246396 117376 246448 117428
rect 265900 117376 265952 117428
rect 207664 117308 207716 117360
rect 213920 117308 213972 117360
rect 235264 117308 235316 117360
rect 265164 117308 265216 117360
rect 230664 117240 230716 117292
rect 245108 117240 245160 117292
rect 282184 117240 282236 117292
rect 306656 117240 306708 117292
rect 231492 117172 231544 117224
rect 239588 117172 239640 117224
rect 282828 117172 282880 117224
rect 305092 117172 305144 117224
rect 231124 117104 231176 117156
rect 233976 117104 234028 117156
rect 169668 116560 169720 116612
rect 203524 116560 203576 116612
rect 259000 116084 259052 116136
rect 265532 116084 265584 116136
rect 181536 116016 181588 116068
rect 214012 116016 214064 116068
rect 245016 116016 245068 116068
rect 265624 116016 265676 116068
rect 169300 115948 169352 116000
rect 213920 115948 213972 116000
rect 234068 115948 234120 116000
rect 264428 115948 264480 116000
rect 281724 115880 281776 115932
rect 302424 115880 302476 115932
rect 282092 115812 282144 115864
rect 298744 115812 298796 115864
rect 231216 115472 231268 115524
rect 238024 115472 238076 115524
rect 230572 115200 230624 115252
rect 259092 115200 259144 115252
rect 260288 114588 260340 114640
rect 265440 114588 265492 114640
rect 172060 114520 172112 114572
rect 213920 114520 213972 114572
rect 243636 114520 243688 114572
rect 265624 114520 265676 114572
rect 231768 114452 231820 114504
rect 240968 114452 241020 114504
rect 282276 114452 282328 114504
rect 303804 114452 303856 114504
rect 231492 114384 231544 114436
rect 239404 114384 239456 114436
rect 282644 114384 282696 114436
rect 292580 114384 292632 114436
rect 168196 113636 168248 113688
rect 173348 113636 173400 113688
rect 250628 113296 250680 113348
rect 265532 113296 265584 113348
rect 188528 113228 188580 113280
rect 213920 113228 213972 113280
rect 242348 113228 242400 113280
rect 265440 113228 265492 113280
rect 174820 113160 174872 113212
rect 214012 113160 214064 113212
rect 229836 113160 229888 113212
rect 265900 113160 265952 113212
rect 231768 113092 231820 113144
rect 258816 113092 258868 113144
rect 282092 113092 282144 113144
rect 295340 113092 295392 113144
rect 231676 112820 231728 112872
rect 238208 112820 238260 112872
rect 231124 112412 231176 112464
rect 243820 112412 243872 112464
rect 258724 111936 258776 111988
rect 265624 111936 265676 111988
rect 169208 111868 169260 111920
rect 214012 111868 214064 111920
rect 253388 111868 253440 111920
rect 265900 111868 265952 111920
rect 166356 111800 166408 111852
rect 213920 111800 213972 111852
rect 239404 111800 239456 111852
rect 265532 111800 265584 111852
rect 3424 111732 3476 111784
rect 11704 111732 11756 111784
rect 168288 111732 168340 111784
rect 169116 111732 169168 111784
rect 231768 111732 231820 111784
rect 264336 111732 264388 111784
rect 282828 111732 282880 111784
rect 298100 111732 298152 111784
rect 231676 111664 231728 111716
rect 236920 111664 236972 111716
rect 230940 111120 230992 111172
rect 235448 111120 235500 111172
rect 238208 110576 238260 110628
rect 265900 110576 265952 110628
rect 191288 110508 191340 110560
rect 214012 110508 214064 110560
rect 256148 110508 256200 110560
rect 265164 110508 265216 110560
rect 178868 110440 178920 110492
rect 213920 110440 213972 110492
rect 231676 110372 231728 110424
rect 260472 110372 260524 110424
rect 282828 110372 282880 110424
rect 291200 110372 291252 110424
rect 231768 110304 231820 110356
rect 253204 110304 253256 110356
rect 231676 109692 231728 109744
rect 236828 109692 236880 109744
rect 260380 109148 260432 109200
rect 265992 109148 266044 109200
rect 188436 109080 188488 109132
rect 213920 109080 213972 109132
rect 257620 109080 257672 109132
rect 265900 109080 265952 109132
rect 169116 109012 169168 109064
rect 214012 109012 214064 109064
rect 243728 109012 243780 109064
rect 265532 109012 265584 109064
rect 167920 108944 167972 108996
rect 174636 108944 174688 108996
rect 231676 108944 231728 108996
rect 250720 108944 250772 108996
rect 282828 108944 282880 108996
rect 310612 108944 310664 108996
rect 231768 108876 231820 108928
rect 245200 108876 245252 108928
rect 231584 108400 231636 108452
rect 234160 108400 234212 108452
rect 238300 107856 238352 107908
rect 265900 107856 265952 107908
rect 250536 107788 250588 107840
rect 265992 107788 266044 107840
rect 178960 107720 179012 107772
rect 214012 107720 214064 107772
rect 245108 107720 245160 107772
rect 264520 107720 264572 107772
rect 174728 107652 174780 107704
rect 213920 107652 213972 107704
rect 261760 107652 261812 107704
rect 265348 107652 265400 107704
rect 231768 107584 231820 107636
rect 257528 107584 257580 107636
rect 231492 107108 231544 107160
rect 233884 107108 233936 107160
rect 230756 106632 230808 106684
rect 235540 106632 235592 106684
rect 240968 106428 241020 106480
rect 265900 106428 265952 106480
rect 170404 106360 170456 106412
rect 214012 106360 214064 106412
rect 249248 106360 249300 106412
rect 265992 106360 266044 106412
rect 167920 106292 167972 106344
rect 213920 106292 213972 106344
rect 231492 106224 231544 106276
rect 261576 106224 261628 106276
rect 231768 106156 231820 106208
rect 242256 106156 242308 106208
rect 282828 105068 282880 105120
rect 287244 105068 287296 105120
rect 263140 105000 263192 105052
rect 265256 105000 265308 105052
rect 210608 104932 210660 104984
rect 214012 104932 214064 104984
rect 253480 104932 253532 104984
rect 265900 104932 265952 104984
rect 176108 104864 176160 104916
rect 213920 104864 213972 104916
rect 242164 104864 242216 104916
rect 265624 104864 265676 104916
rect 230572 104796 230624 104848
rect 232596 104796 232648 104848
rect 230480 104116 230532 104168
rect 254768 104116 254820 104168
rect 258816 103980 258868 104032
rect 265624 103980 265676 104032
rect 247868 103572 247920 103624
rect 265992 103572 266044 103624
rect 206468 103504 206520 103556
rect 213920 103504 213972 103556
rect 233976 103504 234028 103556
rect 265900 103504 265952 103556
rect 231584 102756 231636 102808
rect 250812 102756 250864 102808
rect 257528 102280 257580 102332
rect 265348 102280 265400 102332
rect 232596 102212 232648 102264
rect 211896 102144 211948 102196
rect 213920 102144 213972 102196
rect 230940 102144 230992 102196
rect 232780 102144 232832 102196
rect 236920 102212 236972 102264
rect 265532 102212 265584 102264
rect 265624 102144 265676 102196
rect 230572 102076 230624 102128
rect 264612 102076 264664 102128
rect 230756 101940 230808 101992
rect 232688 101940 232740 101992
rect 231676 101396 231728 101448
rect 252100 101396 252152 101448
rect 250720 100852 250772 100904
rect 265900 100852 265952 100904
rect 210516 100784 210568 100836
rect 214012 100784 214064 100836
rect 252008 100784 252060 100836
rect 265992 100784 266044 100836
rect 200856 100716 200908 100768
rect 213920 100716 213972 100768
rect 231492 100648 231544 100700
rect 253572 100648 253624 100700
rect 471244 100648 471296 100700
rect 580172 100648 580224 100700
rect 231768 100580 231820 100632
rect 249340 100580 249392 100632
rect 254768 99492 254820 99544
rect 265900 99492 265952 99544
rect 253204 99424 253256 99476
rect 265624 99424 265676 99476
rect 166540 99356 166592 99408
rect 213920 99356 213972 99408
rect 246580 99356 246632 99408
rect 265164 99356 265216 99408
rect 231768 99288 231820 99340
rect 267096 99288 267148 99340
rect 231492 98608 231544 98660
rect 238392 98608 238444 98660
rect 166448 98064 166500 98116
rect 214012 98064 214064 98116
rect 242256 98064 242308 98116
rect 261208 98064 261260 98116
rect 164884 97996 164936 98048
rect 213920 97996 213972 98048
rect 238024 97996 238076 98048
rect 264612 97996 264664 98048
rect 3424 97928 3476 97980
rect 14464 97928 14516 97980
rect 236828 96704 236880 96756
rect 265992 96704 266044 96756
rect 231124 96636 231176 96688
rect 265348 96636 265400 96688
rect 209136 96568 209188 96620
rect 229100 96568 229152 96620
rect 230572 96568 230624 96620
rect 189724 96364 189776 96416
rect 281632 96364 281684 96416
rect 231768 95888 231820 95940
rect 268016 95888 268068 95940
rect 228364 95208 228416 95260
rect 265532 95208 265584 95260
rect 184204 95140 184256 95192
rect 281540 95140 281592 95192
rect 199384 95072 199436 95124
rect 281724 95072 281776 95124
rect 216128 95004 216180 95056
rect 279424 95004 279476 95056
rect 222844 94460 222896 94512
rect 267188 94460 267240 94512
rect 133144 94120 133196 94172
rect 171876 94120 171928 94172
rect 120632 94052 120684 94104
rect 167828 94052 167880 94104
rect 104348 93984 104400 94036
rect 174820 93984 174872 94036
rect 116676 93916 116728 93968
rect 192576 93916 192628 93968
rect 94964 93848 95016 93900
rect 178960 93848 179012 93900
rect 230572 93848 230624 93900
rect 234160 93848 234212 93900
rect 268016 93780 268068 93832
rect 276940 93780 276992 93832
rect 234160 93712 234212 93764
rect 270960 93712 271012 93764
rect 151728 93440 151780 93492
rect 167644 93440 167696 93492
rect 122104 93372 122156 93424
rect 170588 93372 170640 93424
rect 115848 93304 115900 93356
rect 173440 93304 173492 93356
rect 107752 93236 107804 93288
rect 169300 93236 169352 93288
rect 85672 93168 85724 93220
rect 164884 93168 164936 93220
rect 129740 93100 129792 93152
rect 214564 93100 214616 93152
rect 217232 93100 217284 93152
rect 277400 93100 277452 93152
rect 230480 92488 230532 92540
rect 233884 92488 233936 92540
rect 114468 92420 114520 92472
rect 203616 92420 203668 92472
rect 105728 92352 105780 92404
rect 191196 92352 191248 92404
rect 120264 92284 120316 92336
rect 181444 92284 181496 92336
rect 123208 92216 123260 92268
rect 176016 92216 176068 92268
rect 106832 92148 106884 92200
rect 129740 92148 129792 92200
rect 134432 92148 134484 92200
rect 167736 92148 167788 92200
rect 152096 92080 152148 92132
rect 171784 92080 171836 92132
rect 188344 91740 188396 91792
rect 276020 91740 276072 91792
rect 99288 91264 99340 91316
rect 106924 91264 106976 91316
rect 100024 91196 100076 91248
rect 123484 91196 123536 91248
rect 88064 91128 88116 91180
rect 120080 91128 120132 91180
rect 85120 91060 85172 91112
rect 133144 91060 133196 91112
rect 67548 90992 67600 91044
rect 214656 90992 214708 91044
rect 180248 90924 180300 90976
rect 280252 90924 280304 90976
rect 120080 90856 120132 90908
rect 214840 90856 214892 90908
rect 124128 90788 124180 90840
rect 170680 90788 170732 90840
rect 125416 90720 125468 90772
rect 166264 90720 166316 90772
rect 109684 90652 109736 90704
rect 181536 90652 181588 90704
rect 67364 89632 67416 89684
rect 210516 89632 210568 89684
rect 126888 89564 126940 89616
rect 195428 89564 195480 89616
rect 101864 89496 101916 89548
rect 169208 89496 169260 89548
rect 112720 89428 112772 89480
rect 177672 89428 177724 89480
rect 119528 89360 119580 89412
rect 170496 89360 170548 89412
rect 136272 89292 136324 89344
rect 187148 89292 187200 89344
rect 196716 88952 196768 89004
rect 265808 88952 265860 89004
rect 89076 88272 89128 88324
rect 166540 88272 166592 88324
rect 122840 88204 122892 88256
rect 200764 88204 200816 88256
rect 107108 88136 107160 88188
rect 172060 88136 172112 88188
rect 151544 88068 151596 88120
rect 211804 88068 211856 88120
rect 118240 88000 118292 88052
rect 177580 88000 177632 88052
rect 129464 87932 129516 87984
rect 182824 87932 182876 87984
rect 105728 86912 105780 86964
rect 213460 86912 213512 86964
rect 90640 86844 90692 86896
rect 176108 86844 176160 86896
rect 119712 86776 119764 86828
rect 184388 86776 184440 86828
rect 151728 86708 151780 86760
rect 196808 86708 196860 86760
rect 3148 85484 3200 85536
rect 35164 85484 35216 85536
rect 67640 85484 67692 85536
rect 216220 85484 216272 85536
rect 67732 85416 67784 85468
rect 214748 85416 214800 85468
rect 91928 85348 91980 85400
rect 167920 85348 167972 85400
rect 111064 85280 111116 85332
rect 177488 85280 177540 85332
rect 130752 85212 130804 85264
rect 189816 85212 189868 85264
rect 122288 85144 122340 85196
rect 173256 85144 173308 85196
rect 75828 84124 75880 84176
rect 216680 84124 216732 84176
rect 103336 84056 103388 84108
rect 188528 84056 188580 84108
rect 117228 83988 117280 84040
rect 178776 83988 178828 84040
rect 126796 83920 126848 83972
rect 180340 83920 180392 83972
rect 180156 83444 180208 83496
rect 265900 83444 265952 83496
rect 110236 82764 110288 82816
rect 210424 82764 210476 82816
rect 114468 82696 114520 82748
rect 213368 82696 213420 82748
rect 97908 82628 97960 82680
rect 169116 82628 169168 82680
rect 103428 82560 103480 82612
rect 174544 82560 174596 82612
rect 125508 82492 125560 82544
rect 169024 82492 169076 82544
rect 111708 81336 111760 81388
rect 207664 81336 207716 81388
rect 93768 81268 93820 81320
rect 170404 81268 170456 81320
rect 104808 81200 104860 81252
rect 175924 81200 175976 81252
rect 100576 81132 100628 81184
rect 166356 81132 166408 81184
rect 126704 81064 126756 81116
rect 184296 81064 184348 81116
rect 180064 80656 180116 80708
rect 287060 80656 287112 80708
rect 115756 79976 115808 80028
rect 209228 79976 209280 80028
rect 86868 79908 86920 79960
rect 166448 79908 166500 79960
rect 95148 79840 95200 79892
rect 174728 79840 174780 79892
rect 99196 79772 99248 79824
rect 171968 79772 172020 79824
rect 113088 79704 113140 79756
rect 185676 79704 185728 79756
rect 96528 78616 96580 78668
rect 188436 78616 188488 78668
rect 128268 78548 128320 78600
rect 213276 78548 213328 78600
rect 123484 78480 123536 78532
rect 191288 78480 191340 78532
rect 110328 78412 110380 78464
rect 173164 78412 173216 78464
rect 133144 77188 133196 77240
rect 200856 77188 200908 77240
rect 118700 76576 118752 76628
rect 256240 76576 256292 76628
rect 4160 76508 4212 76560
rect 228364 76508 228416 76560
rect 106924 75828 106976 75880
rect 192484 75828 192536 75880
rect 99104 75760 99156 75812
rect 178868 75760 178920 75812
rect 67640 75216 67692 75268
rect 263048 75216 263100 75268
rect 64696 75148 64748 75200
rect 281540 75148 281592 75200
rect 124220 73856 124272 73908
rect 230020 73856 230072 73908
rect 64604 73788 64656 73840
rect 269120 73788 269172 73840
rect 80060 72428 80112 72480
rect 242440 72428 242492 72480
rect 3424 71680 3476 71732
rect 47584 71680 47636 71732
rect 74540 71068 74592 71120
rect 261668 71068 261720 71120
rect 64420 71000 64472 71052
rect 273260 71000 273312 71052
rect 77300 69640 77352 69692
rect 254676 69640 254728 69692
rect 81440 68348 81492 68400
rect 262956 68348 263008 68400
rect 46940 68280 46992 68332
rect 236920 68280 236972 68332
rect 85580 66920 85632 66972
rect 260196 66920 260248 66972
rect 53840 66852 53892 66904
rect 247868 66852 247920 66904
rect 88340 65560 88392 65612
rect 243544 65560 243596 65612
rect 64880 65492 64932 65544
rect 253480 65492 253532 65544
rect 69020 64132 69072 64184
rect 263140 64132 263192 64184
rect 75920 62772 75972 62824
rect 249248 62772 249300 62824
rect 60740 61412 60792 61464
rect 246488 61412 246540 61464
rect 78680 61344 78732 61396
rect 264520 61344 264572 61396
rect 358084 60664 358136 60716
rect 580172 60664 580224 60716
rect 82820 60052 82872 60104
rect 238300 60052 238352 60104
rect 49700 59984 49752 60036
rect 257436 59984 257488 60036
rect 3056 59304 3108 59356
rect 53104 59304 53156 59356
rect 85672 58692 85724 58744
rect 245108 58692 245160 58744
rect 52460 58624 52512 58676
rect 265716 58624 265768 58676
rect 89720 57264 89772 57316
rect 261760 57264 261812 57316
rect 9680 57196 9732 57248
rect 253296 57196 253348 57248
rect 96620 55904 96672 55956
rect 257620 55904 257672 55956
rect 41420 55836 41472 55888
rect 234068 55836 234120 55888
rect 100760 54544 100812 54596
rect 260380 54544 260432 54596
rect 34520 54476 34572 54528
rect 243636 54476 243688 54528
rect 103520 53116 103572 53168
rect 243728 53116 243780 53168
rect 30380 53048 30432 53100
rect 260288 53048 260340 53100
rect 107660 51688 107712 51740
rect 238208 51688 238260 51740
rect 106280 50396 106332 50448
rect 229928 50396 229980 50448
rect 16580 50328 16632 50380
rect 246580 50328 246632 50380
rect 118792 49036 118844 49088
rect 253388 49036 253440 49088
rect 17960 48968 18012 49020
rect 242348 48968 242400 49020
rect 110420 47608 110472 47660
rect 256148 47608 256200 47660
rect 22100 47540 22152 47592
rect 250628 47540 250680 47592
rect 177396 46860 177448 46912
rect 580172 46860 580224 46912
rect 122840 46248 122892 46300
rect 238116 46248 238168 46300
rect 86960 46180 87012 46232
rect 258908 46180 258960 46232
rect 3424 45500 3476 45552
rect 40684 45500 40736 45552
rect 113180 44888 113232 44940
rect 240876 44888 240928 44940
rect 48320 44820 48372 44872
rect 259000 44820 259052 44872
rect 20720 43392 20772 43444
rect 254768 43392 254820 43444
rect 35900 42100 35952 42152
rect 235356 42100 235408 42152
rect 26240 42032 26292 42084
rect 250720 42032 250772 42084
rect 29000 40672 29052 40724
rect 252008 40672 252060 40724
rect 45560 39380 45612 39432
rect 239496 39380 239548 39432
rect 35992 39312 36044 39364
rect 257528 39312 257580 39364
rect 40040 37952 40092 38004
rect 261576 37952 261628 38004
rect 31760 37884 31812 37936
rect 256056 37884 256108 37936
rect 2780 36592 2832 36644
rect 236828 36592 236880 36644
rect 37188 36524 37240 36576
rect 280160 36524 280212 36576
rect 44180 35232 44232 35284
rect 232596 35232 232648 35284
rect 27712 35164 27764 35216
rect 247776 35164 247828 35216
rect 93860 33804 93912 33856
rect 250536 33804 250588 33856
rect 44272 33736 44324 33788
rect 245016 33736 245068 33788
rect 3516 33056 3568 33108
rect 51724 33056 51776 33108
rect 187056 33056 187108 33108
rect 580172 33056 580224 33108
rect 109040 32444 109092 32496
rect 261484 32444 261536 32496
rect 51080 32376 51132 32428
rect 233976 32376 234028 32428
rect 114560 31016 114612 31068
rect 264428 31016 264480 31068
rect 71780 29656 71832 29708
rect 240968 29656 241020 29708
rect 19340 29588 19392 29640
rect 249156 29588 249208 29640
rect 57980 28296 58032 28348
rect 258816 28296 258868 28348
rect 23480 28228 23532 28280
rect 250444 28228 250496 28280
rect 110512 26936 110564 26988
rect 251916 26936 251968 26988
rect 6920 26868 6972 26920
rect 242256 26868 242308 26920
rect 120080 25508 120132 25560
rect 236736 25508 236788 25560
rect 102140 22856 102192 22908
rect 236644 22856 236696 22908
rect 63408 22788 63460 22840
rect 284392 22788 284444 22840
rect 20 22720 72 22772
rect 230480 22720 230532 22772
rect 52552 21428 52604 21480
rect 246396 21428 246448 21480
rect 11060 21360 11112 21412
rect 253204 21360 253256 21412
rect 3424 20612 3476 20664
rect 29644 20612 29696 20664
rect 195336 20000 195388 20052
rect 271880 20000 271932 20052
rect 98000 19932 98052 19984
rect 260104 19932 260156 19984
rect 206376 18708 206428 18760
rect 285680 18708 285732 18760
rect 104900 18640 104952 18692
rect 222844 18640 222896 18692
rect 8300 18572 8352 18624
rect 239404 18572 239456 18624
rect 196624 17348 196676 17400
rect 241520 17348 241572 17400
rect 77392 17280 77444 17332
rect 249064 17280 249116 17332
rect 55220 17212 55272 17264
rect 255964 17212 256016 17264
rect 204904 15988 204956 16040
rect 276112 15988 276164 16040
rect 122288 15920 122340 15972
rect 258724 15920 258776 15972
rect 69848 15852 69900 15904
rect 247684 15852 247736 15904
rect 202144 14560 202196 14612
rect 268384 14560 268436 14612
rect 102232 14492 102284 14544
rect 232504 14492 232556 14544
rect 33600 14424 33652 14476
rect 264336 14424 264388 14476
rect 198004 13200 198056 13252
rect 261760 13200 261812 13252
rect 63224 13132 63276 13184
rect 246304 13132 246356 13184
rect 13544 13064 13596 13116
rect 229836 13064 229888 13116
rect 199476 11772 199528 11824
rect 292580 11772 292632 11824
rect 15936 11704 15988 11756
rect 265624 11704 265676 11756
rect 91560 10344 91612 10396
rect 257344 10344 257396 10396
rect 25320 10276 25372 10328
rect 238024 10276 238076 10328
rect 198096 9120 198148 9172
rect 262956 9120 263008 9172
rect 39672 9052 39724 9104
rect 132960 9052 133012 9104
rect 203524 9052 203576 9104
rect 271236 9052 271288 9104
rect 95148 8984 95200 9036
rect 262864 8984 262916 9036
rect 11152 8916 11204 8968
rect 231124 8916 231176 8968
rect 34428 7692 34480 7744
rect 136456 7692 136508 7744
rect 191104 7692 191156 7744
rect 239312 7692 239364 7744
rect 112812 7624 112864 7676
rect 244924 7624 244976 7676
rect 66720 7556 66772 7608
rect 264244 7556 264296 7608
rect 2964 6604 3016 6656
rect 4804 6604 4856 6656
rect 204996 6332 205048 6384
rect 260656 6332 260708 6384
rect 44088 6264 44140 6316
rect 129372 6264 129424 6316
rect 206284 6264 206336 6316
rect 283104 6264 283156 6316
rect 59636 6196 59688 6248
rect 235264 6196 235316 6248
rect 73804 6128 73856 6180
rect 254584 6128 254636 6180
rect 193864 4972 193916 5024
rect 244096 4972 244148 5024
rect 213184 4904 213236 4956
rect 264152 4904 264204 4956
rect 96252 4836 96304 4888
rect 229744 4836 229796 4888
rect 62028 4768 62080 4820
rect 242164 4768 242216 4820
rect 216036 3680 216088 3732
rect 242900 3680 242952 3732
rect 209044 3612 209096 3664
rect 247592 3612 247644 3664
rect 267004 3612 267056 3664
rect 285404 3612 285456 3664
rect 332692 3612 332744 3664
rect 333888 3612 333940 3664
rect 52460 3544 52512 3596
rect 53380 3544 53432 3596
rect 77300 3544 77352 3596
rect 78220 3544 78272 3596
rect 99840 3544 99892 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 6460 3476 6512 3528
rect 98644 3476 98696 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 110420 3544 110472 3596
rect 111616 3544 111668 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 125876 3544 125928 3596
rect 173900 3544 173952 3596
rect 202236 3544 202288 3596
rect 267740 3544 267792 3596
rect 276020 3544 276072 3596
rect 276756 3544 276808 3596
rect 316132 3544 316184 3596
rect 317328 3544 317380 3596
rect 336004 3544 336056 3596
rect 196716 3476 196768 3528
rect 215944 3476 215996 3528
rect 290188 3476 290240 3528
rect 324412 3476 324464 3528
rect 325608 3476 325660 3528
rect 331864 3476 331916 3528
rect 332692 3476 332744 3528
rect 38384 3408 38436 3460
rect 180156 3408 180208 3460
rect 195244 3408 195296 3460
rect 274824 3408 274876 3460
rect 340972 3476 341024 3528
rect 342168 3476 342220 3528
rect 349252 3476 349304 3528
rect 350448 3476 350500 3528
rect 233884 3340 233936 3392
rect 235816 3340 235868 3392
rect 309876 3340 309928 3392
rect 311440 3340 311492 3392
rect 349252 3340 349304 3392
rect 322204 3000 322256 3052
rect 324412 3000 324464 3052
rect 186964 2184 187016 2236
rect 265348 2184 265400 2236
rect 116400 2116 116452 2168
rect 251824 2116 251876 2168
rect 84476 2048 84528 2100
rect 240784 2048 240836 2100
rect 307760 824 307812 876
rect 309048 824 309100 876
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3436 587178 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3516 658144
rect 3568 658135 3570 658144
rect 7564 658164 7616 658170
rect 3516 658106 3568 658112
rect 7564 658106 7616 658112
rect 4804 632120 4856 632126
rect 4804 632062 4856 632068
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 587172 3476 587178
rect 3424 587114 3476 587120
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3252 579766 3280 579935
rect 3240 579760 3292 579766
rect 3240 579702 3292 579708
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3148 554736 3200 554742
rect 3148 554678 3200 554684
rect 3160 553897 3188 554678
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 4816 539578 4844 632062
rect 7576 588606 7604 658106
rect 35164 605872 35216 605878
rect 35164 605814 35216 605820
rect 7564 588600 7616 588606
rect 7564 588542 7616 588548
rect 34244 585268 34296 585274
rect 34244 585210 34296 585216
rect 11704 582752 11756 582758
rect 11704 582694 11756 582700
rect 7564 579760 7616 579766
rect 7564 579702 7616 579708
rect 4804 539572 4856 539578
rect 4804 539514 4856 539520
rect 7576 538218 7604 579702
rect 11716 554742 11744 582694
rect 22744 565888 22796 565894
rect 22744 565830 22796 565836
rect 11704 554736 11756 554742
rect 11704 554678 11756 554684
rect 22756 544406 22784 565830
rect 22744 544400 22796 544406
rect 22744 544342 22796 544348
rect 33140 544400 33192 544406
rect 33140 544342 33192 544348
rect 33152 543794 33180 544342
rect 33140 543788 33192 543794
rect 33140 543730 33192 543736
rect 7564 538212 7616 538218
rect 7564 538154 7616 538160
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 4804 514820 4856 514826
rect 2780 514762 2832 514768
rect 4804 514762 4856 514768
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3528 494766 3556 501735
rect 4816 497486 4844 514762
rect 4804 497480 4856 497486
rect 4804 497422 4856 497428
rect 3516 494760 3568 494766
rect 3516 494702 3568 494708
rect 34256 485790 34284 585210
rect 34428 575544 34480 575550
rect 34428 575486 34480 575492
rect 34336 543788 34388 543794
rect 34336 543730 34388 543736
rect 34244 485784 34296 485790
rect 34244 485726 34296 485732
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 7564 474768 7616 474774
rect 7564 474710 7616 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 7576 439210 7604 474710
rect 33046 474056 33102 474065
rect 33046 473991 33102 474000
rect 30288 470620 30340 470626
rect 30288 470562 30340 470568
rect 22744 462392 22796 462398
rect 22744 462334 22796 462340
rect 7564 439204 7616 439210
rect 7564 439146 7616 439152
rect 22756 438870 22784 462334
rect 22744 438864 22796 438870
rect 22744 438806 22796 438812
rect 3424 429888 3476 429894
rect 3424 429830 3476 429836
rect 3436 410553 3464 429830
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 25504 387932 25556 387938
rect 25504 387874 25556 387880
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 22744 357468 22796 357474
rect 22744 357410 22796 357416
rect 11704 352572 11756 352578
rect 11704 352514 11756 352520
rect 3332 347064 3384 347070
rect 3332 347006 3384 347012
rect 3344 345409 3372 347006
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3424 327140 3476 327146
rect 3424 327082 3476 327088
rect 3436 293185 3464 327082
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3528 311846 3556 319223
rect 3516 311840 3568 311846
rect 3516 311782 3568 311788
rect 11716 306338 11744 352514
rect 22756 346390 22784 357410
rect 25516 347070 25544 387874
rect 30300 376009 30328 470562
rect 33060 378826 33088 473991
rect 34152 458856 34204 458862
rect 34152 458798 34204 458804
rect 33048 378820 33100 378826
rect 33048 378762 33100 378768
rect 30286 376000 30342 376009
rect 30286 375935 30342 375944
rect 34164 362234 34192 458798
rect 34244 452668 34296 452674
rect 34244 452610 34296 452616
rect 34152 362228 34204 362234
rect 34152 362170 34204 362176
rect 34152 356108 34204 356114
rect 34152 356050 34204 356056
rect 25504 347064 25556 347070
rect 25504 347006 25556 347012
rect 22744 346384 22796 346390
rect 22744 346326 22796 346332
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 11704 306332 11756 306338
rect 11704 306274 11756 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 29644 295792 29696 295798
rect 29644 295734 29696 295740
rect 17224 295384 17276 295390
rect 17224 295326 17276 295332
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 4804 279472 4856 279478
rect 4804 279414 4856 279420
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240174 3464 241023
rect 3424 240168 3476 240174
rect 3424 240110 3476 240116
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 4160 76560 4212 76566
rect 4160 76502 4212 76508
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2780 36644 2832 36650
rect 2780 36586 2832 36592
rect 1398 24168 1454 24177
rect 1398 24103 1454 24112
rect 20 22772 72 22778
rect 20 22714 72 22720
rect 32 16574 60 22714
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 24103
rect 2792 3534 2820 36586
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2870 25528 2926 25537
rect 2870 25463 2926 25472
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 25463
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 76502
rect 4172 16546 4752 16574
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6497 3004 6598
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 4724 3482 4752 16546
rect 4816 6662 4844 279414
rect 14464 266416 14516 266422
rect 14464 266358 14516 266364
rect 14476 237318 14504 266358
rect 15844 257372 15896 257378
rect 15844 257314 15896 257320
rect 14464 237312 14516 237318
rect 14464 237254 14516 237260
rect 14464 203584 14516 203590
rect 14464 203526 14516 203532
rect 11704 175976 11756 175982
rect 11704 175918 11756 175924
rect 11716 111790 11744 175918
rect 11704 111784 11756 111790
rect 11704 111726 11756 111732
rect 14476 97986 14504 203526
rect 15856 137970 15884 257314
rect 17236 189038 17264 295326
rect 25504 294636 25556 294642
rect 25504 294578 25556 294584
rect 22744 264240 22796 264246
rect 22744 264182 22796 264188
rect 17316 253972 17368 253978
rect 17316 253914 17368 253920
rect 17328 235958 17356 253914
rect 17316 235952 17368 235958
rect 17316 235894 17368 235900
rect 22756 215286 22784 264182
rect 22744 215280 22796 215286
rect 22744 215222 22796 215228
rect 17224 189032 17276 189038
rect 17224 188974 17276 188980
rect 25516 164218 25544 294578
rect 25504 164212 25556 164218
rect 25504 164154 25556 164160
rect 15844 137964 15896 137970
rect 15844 137906 15896 137912
rect 14464 97980 14516 97986
rect 14464 97922 14516 97928
rect 13818 62792 13874 62801
rect 13818 62727 13874 62736
rect 9680 57248 9732 57254
rect 9680 57190 9732 57196
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6932 16574 6960 26862
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 16574 8340 18566
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 6460 3528 6512 3534
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 4724 3454 5304 3482
rect 6460 3470 6512 3476
rect 5276 480 5304 3454
rect 6472 480 6500 3470
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 57190
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11072 16574 11100 21354
rect 13832 16574 13860 62727
rect 27618 51776 27674 51785
rect 27618 51711 27674 51720
rect 16580 50380 16632 50386
rect 16580 50322 16632 50328
rect 16592 16574 16620 50322
rect 17960 49020 18012 49026
rect 17960 48962 18012 48968
rect 11072 16546 11928 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 480 11192 8910
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13544 13116 13596 13122
rect 13544 13058 13596 13064
rect 13556 480 13584 13058
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 480 15976 11698
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 48962
rect 22100 47592 22152 47598
rect 22100 47534 22152 47540
rect 20720 43444 20772 43450
rect 20720 43386 20772 43392
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19352 6914 19380 29582
rect 19430 19952 19486 19961
rect 19430 19887 19486 19896
rect 19444 16574 19472 19887
rect 20732 16574 20760 43386
rect 22112 16574 22140 47534
rect 26240 42084 26292 42090
rect 26240 42026 26292 42032
rect 23480 28280 23532 28286
rect 23480 28222 23532 28228
rect 23492 16574 23520 28222
rect 19444 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 19352 6886 19472 6914
rect 19444 480 19472 6886
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25320 10328 25372 10334
rect 25320 10270 25372 10276
rect 25332 480 25360 10270
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 42026
rect 27632 6914 27660 51711
rect 29000 40724 29052 40730
rect 29000 40666 29052 40672
rect 27712 35216 27764 35222
rect 27712 35158 27764 35164
rect 27724 16574 27752 35158
rect 29012 16574 29040 40666
rect 29656 20670 29684 295734
rect 32404 290488 32456 290494
rect 32404 290430 32456 290436
rect 32416 150414 32444 290430
rect 34164 280158 34192 356050
rect 34256 352578 34284 452610
rect 34348 443086 34376 543730
rect 34336 443080 34388 443086
rect 34336 443022 34388 443028
rect 34336 383716 34388 383722
rect 34336 383658 34388 383664
rect 34244 352572 34296 352578
rect 34244 352514 34296 352520
rect 33140 280152 33192 280158
rect 33140 280094 33192 280100
rect 34152 280152 34204 280158
rect 34152 280094 34204 280100
rect 33152 279478 33180 280094
rect 33140 279472 33192 279478
rect 33140 279414 33192 279420
rect 34348 235958 34376 383658
rect 34336 235952 34388 235958
rect 34336 235894 34388 235900
rect 32404 150408 32456 150414
rect 32404 150350 32456 150356
rect 30380 53100 30432 53106
rect 30380 53042 30432 53048
rect 29644 20664 29696 20670
rect 29644 20606 29696 20612
rect 30392 16574 30420 53042
rect 31760 37936 31812 37942
rect 31760 37878 31812 37884
rect 31772 16574 31800 37878
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 33612 480 33640 14418
rect 34440 7750 34468 575486
rect 35176 536790 35204 605814
rect 40052 591326 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 76564 703044 76616 703050
rect 76564 702986 76616 702992
rect 68928 702500 68980 702506
rect 68928 702442 68980 702448
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 57888 697604 57940 697610
rect 57888 697546 57940 697552
rect 40040 591320 40092 591326
rect 40040 591262 40092 591268
rect 55864 591320 55916 591326
rect 55864 591262 55916 591268
rect 53840 587172 53892 587178
rect 53840 587114 53892 587120
rect 46848 586628 46900 586634
rect 46848 586570 46900 586576
rect 41236 586560 41288 586566
rect 41236 586502 41288 586508
rect 37004 584112 37056 584118
rect 37004 584054 37056 584060
rect 35624 581052 35676 581058
rect 35624 580994 35676 581000
rect 35164 536784 35216 536790
rect 35164 536726 35216 536732
rect 35164 485784 35216 485790
rect 35164 485726 35216 485732
rect 35176 399498 35204 485726
rect 35636 483002 35664 580994
rect 35716 554804 35768 554810
rect 35716 554746 35768 554752
rect 35624 482996 35676 483002
rect 35624 482938 35676 482944
rect 35728 455394 35756 554746
rect 37016 490618 37044 584054
rect 39948 580304 40000 580310
rect 39948 580246 40000 580252
rect 39304 569968 39356 569974
rect 39304 569910 39356 569916
rect 37188 545760 37240 545766
rect 37188 545702 37240 545708
rect 37096 539640 37148 539646
rect 37096 539582 37148 539588
rect 35808 490612 35860 490618
rect 35808 490554 35860 490560
rect 37004 490612 37056 490618
rect 37004 490554 37056 490560
rect 35716 455388 35768 455394
rect 35716 455330 35768 455336
rect 35716 443012 35768 443018
rect 35716 442954 35768 442960
rect 35164 399492 35216 399498
rect 35164 399434 35216 399440
rect 35728 346390 35756 442954
rect 35820 387870 35848 490554
rect 36912 458244 36964 458250
rect 36912 458186 36964 458192
rect 35808 387864 35860 387870
rect 35808 387806 35860 387812
rect 35716 346384 35768 346390
rect 35716 346326 35768 346332
rect 35728 345710 35756 346326
rect 35716 345704 35768 345710
rect 35716 345646 35768 345652
rect 35820 258058 35848 387806
rect 36924 363662 36952 458186
rect 37004 443080 37056 443086
rect 37004 443022 37056 443028
rect 36912 363656 36964 363662
rect 36912 363598 36964 363604
rect 36924 362982 36952 363598
rect 36912 362976 36964 362982
rect 36912 362918 36964 362924
rect 37016 342922 37044 443022
rect 37108 439521 37136 539582
rect 37200 445738 37228 545702
rect 38568 543856 38620 543862
rect 38568 543798 38620 543804
rect 38476 536104 38528 536110
rect 38476 536046 38528 536052
rect 37188 445732 37240 445738
rect 37188 445674 37240 445680
rect 37094 439512 37150 439521
rect 37094 439447 37150 439456
rect 38488 434722 38516 536046
rect 38580 445058 38608 543798
rect 39316 470558 39344 569910
rect 39764 525836 39816 525842
rect 39764 525778 39816 525784
rect 39672 476128 39724 476134
rect 39672 476070 39724 476076
rect 39304 470552 39356 470558
rect 39304 470494 39356 470500
rect 38568 445052 38620 445058
rect 38568 444994 38620 445000
rect 38580 443018 38608 444994
rect 38568 443012 38620 443018
rect 38568 442954 38620 442960
rect 38568 442332 38620 442338
rect 38568 442274 38620 442280
rect 38476 434716 38528 434722
rect 38476 434658 38528 434664
rect 37188 367124 37240 367130
rect 37188 367066 37240 367072
rect 37096 362976 37148 362982
rect 37096 362918 37148 362924
rect 37004 342916 37056 342922
rect 37004 342858 37056 342864
rect 34520 258052 34572 258058
rect 34520 257994 34572 258000
rect 35808 258052 35860 258058
rect 35808 257994 35860 258000
rect 34532 257378 34560 257994
rect 34520 257372 34572 257378
rect 34520 257314 34572 257320
rect 35164 253224 35216 253230
rect 35164 253166 35216 253172
rect 35176 85542 35204 253166
rect 37108 240106 37136 362918
rect 37096 240100 37148 240106
rect 37096 240042 37148 240048
rect 37108 238814 37136 240042
rect 37096 238808 37148 238814
rect 37096 238750 37148 238756
rect 35164 85536 35216 85542
rect 35164 85478 35216 85484
rect 34520 54528 34572 54534
rect 34520 54470 34572 54476
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 54470
rect 35900 42152 35952 42158
rect 35900 42094 35952 42100
rect 35912 6914 35940 42094
rect 35992 39364 36044 39370
rect 35992 39306 36044 39312
rect 36004 16574 36032 39306
rect 37200 36582 37228 367066
rect 38488 338065 38516 434658
rect 38580 340882 38608 442274
rect 38568 340876 38620 340882
rect 38568 340818 38620 340824
rect 38474 338056 38530 338065
rect 38474 337991 38530 338000
rect 38658 40624 38714 40633
rect 38658 40559 38714 40568
rect 37188 36576 37240 36582
rect 37188 36518 37240 36524
rect 38672 16574 38700 40559
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38396 480 38424 3402
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39684 9110 39712 476070
rect 39776 442950 39804 525778
rect 39960 489914 39988 580246
rect 41144 547936 41196 547942
rect 41144 547878 41196 547884
rect 39868 489886 39988 489914
rect 39868 480214 39896 489886
rect 39856 480208 39908 480214
rect 39856 480150 39908 480156
rect 39764 442944 39816 442950
rect 39764 442886 39816 442892
rect 39776 442338 39804 442886
rect 39764 442332 39816 442338
rect 39764 442274 39816 442280
rect 39764 394936 39816 394942
rect 39764 394878 39816 394884
rect 39776 274650 39804 394878
rect 39868 389230 39896 480150
rect 40684 455388 40736 455394
rect 40684 455330 40736 455336
rect 39856 389224 39908 389230
rect 39856 389166 39908 389172
rect 39764 274644 39816 274650
rect 39764 274586 39816 274592
rect 39868 249762 39896 389166
rect 40696 357406 40724 455330
rect 41156 449206 41184 547878
rect 41248 494086 41276 586502
rect 46756 585200 46808 585206
rect 46756 585142 46808 585148
rect 43812 581324 43864 581330
rect 43812 581266 43864 581272
rect 42708 550656 42760 550662
rect 42708 550598 42760 550604
rect 41328 539708 41380 539714
rect 41328 539650 41380 539656
rect 41236 494080 41288 494086
rect 41236 494022 41288 494028
rect 41144 449200 41196 449206
rect 41144 449142 41196 449148
rect 41156 447982 41184 449142
rect 41144 447976 41196 447982
rect 41144 447918 41196 447924
rect 41248 391270 41276 494022
rect 41340 439006 41368 539650
rect 42616 534880 42668 534886
rect 42616 534822 42668 534828
rect 42524 469872 42576 469878
rect 42524 469814 42576 469820
rect 42064 447976 42116 447982
rect 42064 447918 42116 447924
rect 41328 439000 41380 439006
rect 41328 438942 41380 438948
rect 41236 391264 41288 391270
rect 41236 391206 41288 391212
rect 41236 387932 41288 387938
rect 41236 387874 41288 387880
rect 40684 357400 40736 357406
rect 40684 357342 40736 357348
rect 41144 342916 41196 342922
rect 41144 342858 41196 342864
rect 41156 267714 41184 342858
rect 41248 297430 41276 387874
rect 41340 336734 41368 438942
rect 41420 352572 41472 352578
rect 41420 352514 41472 352520
rect 41432 351966 41460 352514
rect 41420 351960 41472 351966
rect 41420 351902 41472 351908
rect 42076 349178 42104 447918
rect 42536 373998 42564 469814
rect 42628 437374 42656 534822
rect 42720 451926 42748 550598
rect 43824 482934 43852 581266
rect 45468 558952 45520 558958
rect 45468 558894 45520 558900
rect 43904 556232 43956 556238
rect 43904 556174 43956 556180
rect 43812 482928 43864 482934
rect 43812 482870 43864 482876
rect 43916 457502 43944 556174
rect 44088 549296 44140 549302
rect 44088 549238 44140 549244
rect 43996 493332 44048 493338
rect 43996 493274 44048 493280
rect 43904 457496 43956 457502
rect 43904 457438 43956 457444
rect 42708 451920 42760 451926
rect 42708 451862 42760 451868
rect 42616 437368 42668 437374
rect 42616 437310 42668 437316
rect 42614 383208 42670 383217
rect 42614 383143 42670 383152
rect 42524 373992 42576 373998
rect 42524 373934 42576 373940
rect 42064 349172 42116 349178
rect 42064 349114 42116 349120
rect 41328 336728 41380 336734
rect 41328 336670 41380 336676
rect 42628 335238 42656 383143
rect 43812 361616 43864 361622
rect 43812 361558 43864 361564
rect 42708 351960 42760 351966
rect 42708 351902 42760 351908
rect 42616 335232 42668 335238
rect 42616 335174 42668 335180
rect 42720 300150 42748 351902
rect 42708 300144 42760 300150
rect 42708 300086 42760 300092
rect 41236 297424 41288 297430
rect 41236 297366 41288 297372
rect 41144 267708 41196 267714
rect 41144 267650 41196 267656
rect 43824 253910 43852 361558
rect 43916 360874 43944 457438
rect 44008 393990 44036 493274
rect 44100 449886 44128 549238
rect 45284 534744 45336 534750
rect 45284 534686 45336 534692
rect 44456 460216 44508 460222
rect 44456 460158 44508 460164
rect 44468 458250 44496 460158
rect 44456 458244 44508 458250
rect 44456 458186 44508 458192
rect 44088 449880 44140 449886
rect 44088 449822 44140 449828
rect 45192 443692 45244 443698
rect 45192 443634 45244 443640
rect 43996 393984 44048 393990
rect 43996 393926 44048 393932
rect 43996 393508 44048 393514
rect 43996 393450 44048 393456
rect 43904 360868 43956 360874
rect 43904 360810 43956 360816
rect 44008 282878 44036 393450
rect 44088 382288 44140 382294
rect 44088 382230 44140 382236
rect 43996 282872 44048 282878
rect 43996 282814 44048 282820
rect 42800 253904 42852 253910
rect 42800 253846 42852 253852
rect 43812 253904 43864 253910
rect 43812 253846 43864 253852
rect 42812 253230 42840 253846
rect 42800 253224 42852 253230
rect 42800 253166 42852 253172
rect 39856 249756 39908 249762
rect 39856 249698 39908 249704
rect 40684 185836 40736 185842
rect 40684 185778 40736 185784
rect 40696 45558 40724 185778
rect 41420 55888 41472 55894
rect 41420 55830 41472 55836
rect 40684 45552 40736 45558
rect 40684 45494 40736 45500
rect 40040 38004 40092 38010
rect 40040 37946 40092 37952
rect 40052 16574 40080 37946
rect 41432 16574 41460 55830
rect 42798 30968 42854 30977
rect 42798 30903 42854 30912
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39672 9104 39724 9110
rect 39672 9046 39724 9052
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 30903
rect 44100 6322 44128 382230
rect 45204 343670 45232 443634
rect 45296 438802 45324 534686
rect 45376 497548 45428 497554
rect 45376 497490 45428 497496
rect 45388 440910 45416 497490
rect 45480 460222 45508 558894
rect 46572 529236 46624 529242
rect 46572 529178 46624 529184
rect 45468 460216 45520 460222
rect 45468 460158 45520 460164
rect 45468 459604 45520 459610
rect 45468 459546 45520 459552
rect 45376 440904 45428 440910
rect 45376 440846 45428 440852
rect 45284 438796 45336 438802
rect 45284 438738 45336 438744
rect 45284 392624 45336 392630
rect 45284 392566 45336 392572
rect 45192 343664 45244 343670
rect 45192 343606 45244 343612
rect 45296 335306 45324 392566
rect 45480 360194 45508 459546
rect 46204 448588 46256 448594
rect 46204 448530 46256 448536
rect 46216 438598 46244 448530
rect 46584 438734 46612 529178
rect 46664 492516 46716 492522
rect 46664 492458 46716 492464
rect 46572 438728 46624 438734
rect 46572 438670 46624 438676
rect 46204 438592 46256 438598
rect 46204 438534 46256 438540
rect 46584 437510 46612 438670
rect 46572 437504 46624 437510
rect 46572 437446 46624 437452
rect 46572 396908 46624 396914
rect 46572 396850 46624 396856
rect 45468 360188 45520 360194
rect 45468 360130 45520 360136
rect 45468 349172 45520 349178
rect 45468 349114 45520 349120
rect 45284 335300 45336 335306
rect 45284 335242 45336 335248
rect 45480 234598 45508 349114
rect 46584 333946 46612 396850
rect 46676 396778 46704 492458
rect 46768 491366 46796 585142
rect 46860 492658 46888 586570
rect 52184 585336 52236 585342
rect 52184 585278 52236 585284
rect 48042 583808 48098 583817
rect 48042 583743 48098 583752
rect 46848 492652 46900 492658
rect 46848 492594 46900 492600
rect 48056 492522 48084 583743
rect 52092 582548 52144 582554
rect 52092 582490 52144 582496
rect 50804 581120 50856 581126
rect 50804 581062 50856 581068
rect 49608 564460 49660 564466
rect 49608 564402 49660 564408
rect 48136 563100 48188 563106
rect 48136 563042 48188 563048
rect 48044 492516 48096 492522
rect 48044 492458 48096 492464
rect 48056 491978 48084 492458
rect 48044 491972 48096 491978
rect 48044 491914 48096 491920
rect 46756 491360 46808 491366
rect 46756 491302 46808 491308
rect 46768 489914 46796 491302
rect 47952 490680 48004 490686
rect 47952 490622 48004 490628
rect 46768 489886 46888 489914
rect 46756 437504 46808 437510
rect 46756 437446 46808 437452
rect 46664 396772 46716 396778
rect 46664 396714 46716 396720
rect 46768 336666 46796 437446
rect 46860 392086 46888 489886
rect 47860 464772 47912 464778
rect 47860 464714 47912 464720
rect 47872 464370 47900 464714
rect 47860 464364 47912 464370
rect 47860 464306 47912 464312
rect 47872 394194 47900 464306
rect 47964 436082 47992 490622
rect 48044 465044 48096 465050
rect 48044 464986 48096 464992
rect 47952 436076 48004 436082
rect 47952 436018 48004 436024
rect 47860 394188 47912 394194
rect 47860 394130 47912 394136
rect 47952 394052 48004 394058
rect 47952 393994 48004 394000
rect 46848 392080 46900 392086
rect 46848 392022 46900 392028
rect 46756 336660 46808 336666
rect 46756 336602 46808 336608
rect 46572 333940 46624 333946
rect 46572 333882 46624 333888
rect 46756 284368 46808 284374
rect 46756 284310 46808 284316
rect 45468 234592 45520 234598
rect 45468 234534 45520 234540
rect 46768 210458 46796 284310
rect 46860 267646 46888 392022
rect 47860 378820 47912 378826
rect 47860 378762 47912 378768
rect 47872 378214 47900 378762
rect 47860 378208 47912 378214
rect 47860 378150 47912 378156
rect 47860 343664 47912 343670
rect 47860 343606 47912 343612
rect 47872 335354 47900 343606
rect 47964 338026 47992 393994
rect 48056 370569 48084 464986
rect 48148 464778 48176 563042
rect 48228 555484 48280 555490
rect 48228 555426 48280 555432
rect 48136 464772 48188 464778
rect 48136 464714 48188 464720
rect 48240 454102 48268 555426
rect 49424 542428 49476 542434
rect 49424 542370 49476 542376
rect 49332 529304 49384 529310
rect 49332 529246 49384 529252
rect 48228 454096 48280 454102
rect 48228 454038 48280 454044
rect 48964 434036 49016 434042
rect 48964 433978 49016 433984
rect 48976 433265 49004 433978
rect 48962 433256 49018 433265
rect 48962 433191 49018 433200
rect 48136 422340 48188 422346
rect 48136 422282 48188 422288
rect 48042 370560 48098 370569
rect 48042 370495 48098 370504
rect 48042 340776 48098 340785
rect 48042 340711 48098 340720
rect 48056 339522 48084 340711
rect 48044 339516 48096 339522
rect 48044 339458 48096 339464
rect 47952 338020 48004 338026
rect 47952 337962 48004 337968
rect 47872 335326 48084 335354
rect 48056 297566 48084 335326
rect 48148 304298 48176 422282
rect 48228 378208 48280 378214
rect 48228 378150 48280 378156
rect 48136 304292 48188 304298
rect 48136 304234 48188 304240
rect 48044 297560 48096 297566
rect 48044 297502 48096 297508
rect 47584 294024 47636 294030
rect 47584 293966 47636 293972
rect 46848 267640 46900 267646
rect 46848 267582 46900 267588
rect 46756 210452 46808 210458
rect 46756 210394 46808 210400
rect 47596 71738 47624 293966
rect 48136 263628 48188 263634
rect 48136 263570 48188 263576
rect 48148 213246 48176 263570
rect 48240 237386 48268 378150
rect 48976 339454 49004 433191
rect 49344 431905 49372 529246
rect 49436 444378 49464 542370
rect 49516 494828 49568 494834
rect 49516 494770 49568 494776
rect 49424 444372 49476 444378
rect 49424 444314 49476 444320
rect 49436 443698 49464 444314
rect 49424 443692 49476 443698
rect 49424 443634 49476 443640
rect 49330 431896 49386 431905
rect 49330 431831 49386 431840
rect 49344 430681 49372 431831
rect 49330 430672 49386 430681
rect 49330 430607 49386 430616
rect 49528 395350 49556 494770
rect 49620 465730 49648 564402
rect 50712 534812 50764 534818
rect 50712 534754 50764 534760
rect 49608 465724 49660 465730
rect 49608 465666 49660 465672
rect 49620 465050 49648 465666
rect 49608 465044 49660 465050
rect 49608 464986 49660 464992
rect 49608 454708 49660 454714
rect 49608 454650 49660 454656
rect 49516 395344 49568 395350
rect 49516 395286 49568 395292
rect 49056 389836 49108 389842
rect 49056 389778 49108 389784
rect 49068 372570 49096 389778
rect 49516 376032 49568 376038
rect 49516 375974 49568 375980
rect 49056 372564 49108 372570
rect 49056 372506 49108 372512
rect 48964 339448 49016 339454
rect 48964 339390 49016 339396
rect 49528 288386 49556 375974
rect 49620 355337 49648 454650
rect 50724 438870 50752 534754
rect 50816 493338 50844 581062
rect 50988 560312 51040 560318
rect 50988 560254 51040 560260
rect 50896 552084 50948 552090
rect 50896 552026 50948 552032
rect 50804 493332 50856 493338
rect 50804 493274 50856 493280
rect 50804 459672 50856 459678
rect 50804 459614 50856 459620
rect 50712 438864 50764 438870
rect 50712 438806 50764 438812
rect 50724 438190 50752 438806
rect 50712 438184 50764 438190
rect 50712 438126 50764 438132
rect 50712 380724 50764 380730
rect 50712 380666 50764 380672
rect 50620 362976 50672 362982
rect 50620 362918 50672 362924
rect 49606 355328 49662 355337
rect 49606 355263 49662 355272
rect 49608 327820 49660 327826
rect 49608 327762 49660 327768
rect 49620 327146 49648 327762
rect 49608 327140 49660 327146
rect 49608 327082 49660 327088
rect 49516 288380 49568 288386
rect 49516 288322 49568 288328
rect 49516 270564 49568 270570
rect 49516 270506 49568 270512
rect 48228 237380 48280 237386
rect 48228 237322 48280 237328
rect 49528 222873 49556 270506
rect 49620 244254 49648 327082
rect 50632 287054 50660 362918
rect 50724 311846 50752 380666
rect 50816 363730 50844 459614
rect 50908 453354 50936 552026
rect 51000 460290 51028 560254
rect 52104 494902 52132 582490
rect 52092 494896 52144 494902
rect 52090 494864 52092 494873
rect 52144 494864 52146 494873
rect 52090 494799 52146 494808
rect 52092 492856 52144 492862
rect 52092 492798 52144 492804
rect 52104 492697 52132 492798
rect 52090 492688 52146 492697
rect 52090 492623 52146 492632
rect 52196 491502 52224 585278
rect 53564 583976 53616 583982
rect 53852 583953 53880 587114
rect 54484 585404 54536 585410
rect 54484 585346 54536 585352
rect 53564 583918 53616 583924
rect 53838 583944 53894 583953
rect 52276 562352 52328 562358
rect 52276 562294 52328 562300
rect 52184 491496 52236 491502
rect 52184 491438 52236 491444
rect 52196 489914 52224 491438
rect 52104 489886 52224 489914
rect 52000 463684 52052 463690
rect 52000 463626 52052 463632
rect 52012 463010 52040 463626
rect 52000 463004 52052 463010
rect 52000 462946 52052 462952
rect 50988 460284 51040 460290
rect 50988 460226 51040 460232
rect 51000 459678 51028 460226
rect 50988 459672 51040 459678
rect 50988 459614 51040 459620
rect 50896 453348 50948 453354
rect 50896 453290 50948 453296
rect 50804 363724 50856 363730
rect 50804 363666 50856 363672
rect 50816 362982 50844 363666
rect 50804 362976 50856 362982
rect 50804 362918 50856 362924
rect 50908 356726 50936 453290
rect 50988 398132 51040 398138
rect 50988 398074 51040 398080
rect 51000 397526 51028 398074
rect 50988 397520 51040 397526
rect 50988 397462 51040 397468
rect 50896 356720 50948 356726
rect 50896 356662 50948 356668
rect 50712 311840 50764 311846
rect 50712 311782 50764 311788
rect 50724 311166 50752 311782
rect 50712 311160 50764 311166
rect 50712 311102 50764 311108
rect 50632 287026 50752 287054
rect 50724 264926 50752 287026
rect 50804 280220 50856 280226
rect 50804 280162 50856 280168
rect 50712 264920 50764 264926
rect 50712 264862 50764 264868
rect 50724 264246 50752 264862
rect 50712 264240 50764 264246
rect 50712 264182 50764 264188
rect 49608 244248 49660 244254
rect 49608 244190 49660 244196
rect 49514 222864 49570 222873
rect 49514 222799 49570 222808
rect 48136 213240 48188 213246
rect 48136 213182 48188 213188
rect 50816 194002 50844 280162
rect 50896 269136 50948 269142
rect 50896 269078 50948 269084
rect 50908 214606 50936 269078
rect 51000 238882 51028 397462
rect 52012 367810 52040 462946
rect 52104 394126 52132 489886
rect 52288 463690 52316 562294
rect 52368 537600 52420 537606
rect 52368 537542 52420 537548
rect 52276 463684 52328 463690
rect 52276 463626 52328 463632
rect 52184 438184 52236 438190
rect 52184 438126 52236 438132
rect 52092 394120 52144 394126
rect 52092 394062 52144 394068
rect 52000 367804 52052 367810
rect 52000 367746 52052 367752
rect 52196 333878 52224 438126
rect 52380 437306 52408 537542
rect 53288 492108 53340 492114
rect 53288 492050 53340 492056
rect 53300 492017 53328 492050
rect 53472 492040 53524 492046
rect 53286 492008 53342 492017
rect 53472 491982 53524 491988
rect 53286 491943 53342 491952
rect 53380 475380 53432 475386
rect 53380 475322 53432 475328
rect 52368 437300 52420 437306
rect 52368 437242 52420 437248
rect 52276 392012 52328 392018
rect 52276 391954 52328 391960
rect 52184 333872 52236 333878
rect 52184 333814 52236 333820
rect 52092 277432 52144 277438
rect 52092 277374 52144 277380
rect 51724 268252 51776 268258
rect 51724 268194 51776 268200
rect 50988 238876 51040 238882
rect 50988 238818 51040 238824
rect 50896 214600 50948 214606
rect 50896 214542 50948 214548
rect 50804 193996 50856 194002
rect 50804 193938 50856 193944
rect 47584 71732 47636 71738
rect 47584 71674 47636 71680
rect 46940 68332 46992 68338
rect 46940 68274 46992 68280
rect 45560 39432 45612 39438
rect 45560 39374 45612 39380
rect 44180 35284 44232 35290
rect 44180 35226 44232 35232
rect 44192 6914 44220 35226
rect 44272 33788 44324 33794
rect 44272 33730 44324 33736
rect 44284 16574 44312 33730
rect 45572 16574 45600 39374
rect 46952 16574 46980 68274
rect 49700 60036 49752 60042
rect 49700 59978 49752 59984
rect 48320 44872 48372 44878
rect 48320 44814 48372 44820
rect 48332 16574 48360 44814
rect 49712 16574 49740 59978
rect 51736 33114 51764 268194
rect 52104 204950 52132 277374
rect 52184 274712 52236 274718
rect 52184 274654 52236 274660
rect 52092 204944 52144 204950
rect 52092 204886 52144 204892
rect 52196 199442 52224 274654
rect 52288 268394 52316 391954
rect 52368 386504 52420 386510
rect 52368 386446 52420 386452
rect 52276 268388 52328 268394
rect 52276 268330 52328 268336
rect 52288 268258 52316 268330
rect 52276 268252 52328 268258
rect 52276 268194 52328 268200
rect 52380 238746 52408 386446
rect 53392 380730 53420 475322
rect 53484 396098 53512 491982
rect 53576 487898 53604 583918
rect 53838 583879 53894 583888
rect 53748 574116 53800 574122
rect 53748 574058 53800 574064
rect 53656 556300 53708 556306
rect 53656 556242 53708 556248
rect 53564 487892 53616 487898
rect 53564 487834 53616 487840
rect 53668 458182 53696 556242
rect 53760 475386 53788 574058
rect 54496 492114 54524 585346
rect 55876 584089 55904 591262
rect 55862 584080 55918 584089
rect 55862 584015 55918 584024
rect 56506 584080 56562 584089
rect 56506 584015 56562 584024
rect 55034 583944 55090 583953
rect 55034 583879 55090 583888
rect 54760 493400 54812 493406
rect 54760 493342 54812 493348
rect 54484 492108 54536 492114
rect 54484 492050 54536 492056
rect 53748 475380 53800 475386
rect 53748 475322 53800 475328
rect 53656 458176 53708 458182
rect 53656 458118 53708 458124
rect 53564 396840 53616 396846
rect 53564 396782 53616 396788
rect 53472 396092 53524 396098
rect 53472 396034 53524 396040
rect 53470 387560 53526 387569
rect 53470 387495 53526 387504
rect 53484 386510 53512 387495
rect 53472 386504 53524 386510
rect 53472 386446 53524 386452
rect 53380 380724 53432 380730
rect 53380 380666 53432 380672
rect 53576 336530 53604 396782
rect 54484 396092 54536 396098
rect 54484 396034 54536 396040
rect 53656 389904 53708 389910
rect 53656 389846 53708 389852
rect 53564 336524 53616 336530
rect 53564 336466 53616 336472
rect 53668 294642 53696 389846
rect 53748 387524 53800 387530
rect 53748 387466 53800 387472
rect 53656 294636 53708 294642
rect 53656 294578 53708 294584
rect 53104 293276 53156 293282
rect 53104 293218 53156 293224
rect 52368 238740 52420 238746
rect 52368 238682 52420 238688
rect 52184 199436 52236 199442
rect 52184 199378 52236 199384
rect 53116 59362 53144 293218
rect 53564 276072 53616 276078
rect 53564 276014 53616 276020
rect 53576 220182 53604 276014
rect 53656 259480 53708 259486
rect 53656 259422 53708 259428
rect 53564 220176 53616 220182
rect 53564 220118 53616 220124
rect 53668 181558 53696 259422
rect 53760 238610 53788 387466
rect 54496 293282 54524 396034
rect 54772 391406 54800 493342
rect 54944 492720 54996 492726
rect 54944 492662 54996 492668
rect 54852 490748 54904 490754
rect 54852 490690 54904 490696
rect 54864 436014 54892 490690
rect 54956 454714 54984 492662
rect 55048 484362 55076 583879
rect 55128 582684 55180 582690
rect 55128 582626 55180 582632
rect 55140 492046 55168 582626
rect 56324 582616 56376 582622
rect 56324 582558 56376 582564
rect 56232 496256 56284 496262
rect 56232 496198 56284 496204
rect 55128 492040 55180 492046
rect 55128 491982 55180 491988
rect 55036 484356 55088 484362
rect 55036 484298 55088 484304
rect 55036 480276 55088 480282
rect 55036 480218 55088 480224
rect 54944 454708 54996 454714
rect 54944 454650 54996 454656
rect 54852 436008 54904 436014
rect 54852 435950 54904 435956
rect 54760 391400 54812 391406
rect 54760 391342 54812 391348
rect 55048 388142 55076 480218
rect 55128 454096 55180 454102
rect 55128 454038 55180 454044
rect 55036 388136 55088 388142
rect 55036 388078 55088 388084
rect 54852 358080 54904 358086
rect 54852 358022 54904 358028
rect 54484 293276 54536 293282
rect 54484 293218 54536 293224
rect 54864 271862 54892 358022
rect 54944 339244 54996 339250
rect 54944 339186 54996 339192
rect 54852 271856 54904 271862
rect 54852 271798 54904 271804
rect 54852 255332 54904 255338
rect 54852 255274 54904 255280
rect 53748 238604 53800 238610
rect 53748 238546 53800 238552
rect 54864 193866 54892 255274
rect 54956 247042 54984 339186
rect 55048 280090 55076 388078
rect 55140 358086 55168 454038
rect 56244 439414 56272 496198
rect 56336 496126 56364 582558
rect 56416 534948 56468 534954
rect 56416 534890 56468 534896
rect 56324 496120 56376 496126
rect 56324 496062 56376 496068
rect 56232 439408 56284 439414
rect 56232 439350 56284 439356
rect 56428 439074 56456 534890
rect 56520 487830 56548 584015
rect 57704 583908 57756 583914
rect 57704 583850 57756 583856
rect 57244 553444 57296 553450
rect 57244 553386 57296 553392
rect 57256 492658 57284 553386
rect 57520 538620 57572 538626
rect 57520 538562 57572 538568
rect 57244 492652 57296 492658
rect 57244 492594 57296 492600
rect 56508 487824 56560 487830
rect 56508 487766 56560 487772
rect 56416 439068 56468 439074
rect 56416 439010 56468 439016
rect 56416 418804 56468 418810
rect 56416 418746 56468 418752
rect 56232 394188 56284 394194
rect 56232 394130 56284 394136
rect 56244 369850 56272 394130
rect 56324 385688 56376 385694
rect 56324 385630 56376 385636
rect 56232 369844 56284 369850
rect 56232 369786 56284 369792
rect 55128 358080 55180 358086
rect 55128 358022 55180 358028
rect 56336 339386 56364 385630
rect 56428 353258 56456 418746
rect 56520 388006 56548 487766
rect 57336 484356 57388 484362
rect 57336 484298 57388 484304
rect 57244 439408 57296 439414
rect 57244 439350 57296 439356
rect 57256 439142 57284 439350
rect 57244 439136 57296 439142
rect 57244 439078 57296 439084
rect 56508 388000 56560 388006
rect 56508 387942 56560 387948
rect 56520 387530 56548 387942
rect 56508 387524 56560 387530
rect 56508 387466 56560 387472
rect 56508 385076 56560 385082
rect 56508 385018 56560 385024
rect 56416 353252 56468 353258
rect 56416 353194 56468 353200
rect 56324 339380 56376 339386
rect 56324 339322 56376 339328
rect 56416 336456 56468 336462
rect 56416 336398 56468 336404
rect 55128 292596 55180 292602
rect 55128 292538 55180 292544
rect 55036 280084 55088 280090
rect 55036 280026 55088 280032
rect 55036 277500 55088 277506
rect 55036 277442 55088 277448
rect 54944 247036 54996 247042
rect 54944 246978 54996 246984
rect 55048 207806 55076 277442
rect 55036 207800 55088 207806
rect 55036 207742 55088 207748
rect 54852 193860 54904 193866
rect 54852 193802 54904 193808
rect 53656 181552 53708 181558
rect 53656 181494 53708 181500
rect 53840 66904 53892 66910
rect 53840 66846 53892 66852
rect 53104 59356 53156 59362
rect 53104 59298 53156 59304
rect 52460 58676 52512 58682
rect 52460 58618 52512 58624
rect 51724 33108 51776 33114
rect 51724 33050 51776 33056
rect 51080 32428 51132 32434
rect 51080 32370 51132 32376
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44088 6316 44140 6322
rect 44088 6258 44140 6264
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 32370
rect 52472 3602 52500 58618
rect 52552 21480 52604 21486
rect 52552 21422 52604 21428
rect 52460 3596 52512 3602
rect 52460 3538 52512 3544
rect 52564 480 52592 21422
rect 53852 16574 53880 66846
rect 55140 24857 55168 292538
rect 56324 262268 56376 262274
rect 56324 262210 56376 262216
rect 56336 207670 56364 262210
rect 56428 253881 56456 336398
rect 56520 284306 56548 385018
rect 57256 339250 57284 439078
rect 57348 388482 57376 484298
rect 57532 437442 57560 538562
rect 57612 497616 57664 497622
rect 57612 497558 57664 497564
rect 57624 439550 57652 497558
rect 57716 492930 57744 583850
rect 57796 581188 57848 581194
rect 57796 581130 57848 581136
rect 57808 537538 57836 581130
rect 57900 556170 57928 697546
rect 57980 670744 58032 670750
rect 57980 670686 58032 670692
rect 57888 556164 57940 556170
rect 57888 556106 57940 556112
rect 57900 555490 57928 556106
rect 57888 555484 57940 555490
rect 57888 555426 57940 555432
rect 57992 539510 58020 670686
rect 59268 584044 59320 584050
rect 59268 583986 59320 583992
rect 59084 581256 59136 581262
rect 59084 581198 59136 581204
rect 57980 539504 58032 539510
rect 57980 539446 58032 539452
rect 57992 538626 58020 539446
rect 59096 538801 59124 581198
rect 59176 578332 59228 578338
rect 59176 578274 59228 578280
rect 59082 538792 59138 538801
rect 59082 538727 59138 538736
rect 57980 538620 58032 538626
rect 57980 538562 58032 538568
rect 59084 537668 59136 537674
rect 59084 537610 59136 537616
rect 57796 537532 57848 537538
rect 57796 537474 57848 537480
rect 58624 512236 58676 512242
rect 58624 512178 58676 512184
rect 57704 492924 57756 492930
rect 57704 492866 57756 492872
rect 57716 489914 57744 492866
rect 57716 489886 57928 489914
rect 57612 439544 57664 439550
rect 57612 439486 57664 439492
rect 57520 437436 57572 437442
rect 57520 437378 57572 437384
rect 57704 392692 57756 392698
rect 57704 392634 57756 392640
rect 57336 388476 57388 388482
rect 57336 388418 57388 388424
rect 57612 387184 57664 387190
rect 57612 387126 57664 387132
rect 57244 339244 57296 339250
rect 57244 339186 57296 339192
rect 57624 337890 57652 387126
rect 57612 337884 57664 337890
rect 57612 337826 57664 337832
rect 57612 334688 57664 334694
rect 57612 334630 57664 334636
rect 56508 284300 56560 284306
rect 56508 284242 56560 284248
rect 56508 273284 56560 273290
rect 56508 273226 56560 273232
rect 56414 253872 56470 253881
rect 56414 253807 56470 253816
rect 56324 207664 56376 207670
rect 56324 207606 56376 207612
rect 56520 193934 56548 273226
rect 57520 269204 57572 269210
rect 57520 269146 57572 269152
rect 57532 217326 57560 269146
rect 57624 266354 57652 334630
rect 57716 332586 57744 392634
rect 57900 386442 57928 489886
rect 58636 480282 58664 512178
rect 58624 480276 58676 480282
rect 58624 480218 58676 480224
rect 58636 480146 58664 480218
rect 58624 480140 58676 480146
rect 58624 480082 58676 480088
rect 58992 472048 59044 472054
rect 58992 471990 59044 471996
rect 58900 387116 58952 387122
rect 58900 387058 58952 387064
rect 57888 386436 57940 386442
rect 57888 386378 57940 386384
rect 57900 373994 57928 386378
rect 57808 373966 57928 373994
rect 57704 332580 57756 332586
rect 57704 332522 57756 332528
rect 57704 314016 57756 314022
rect 57704 313958 57756 313964
rect 57612 266348 57664 266354
rect 57612 266290 57664 266296
rect 57716 245614 57744 313958
rect 57808 294710 57836 373966
rect 58912 339318 58940 387058
rect 59004 377466 59032 471990
rect 59096 438666 59124 537610
rect 59188 512242 59216 578274
rect 59176 512236 59228 512242
rect 59176 512178 59228 512184
rect 59188 512038 59216 512178
rect 59176 512032 59228 512038
rect 59176 511974 59228 511980
rect 59280 493406 59308 583986
rect 61752 583840 61804 583846
rect 61752 583782 61804 583788
rect 60004 583024 60056 583030
rect 60004 582966 60056 582972
rect 60016 539714 60044 582966
rect 60740 563032 60792 563038
rect 60740 562974 60792 562980
rect 60752 562358 60780 562974
rect 60740 562352 60792 562358
rect 60740 562294 60792 562300
rect 60648 546508 60700 546514
rect 60648 546450 60700 546456
rect 60556 542496 60608 542502
rect 60556 542438 60608 542444
rect 60004 539708 60056 539714
rect 60004 539650 60056 539656
rect 60016 538150 60044 539650
rect 60004 538144 60056 538150
rect 60004 538086 60056 538092
rect 59268 493400 59320 493406
rect 59268 493342 59320 493348
rect 59268 492788 59320 492794
rect 59268 492730 59320 492736
rect 59176 487892 59228 487898
rect 59176 487834 59228 487840
rect 59188 487218 59216 487834
rect 59176 487212 59228 487218
rect 59176 487154 59228 487160
rect 59084 438660 59136 438666
rect 59084 438602 59136 438608
rect 59188 388074 59216 487154
rect 59280 389910 59308 492730
rect 60372 490816 60424 490822
rect 60372 490758 60424 490764
rect 60384 435946 60412 490758
rect 60464 465044 60516 465050
rect 60464 464986 60516 464992
rect 60372 435940 60424 435946
rect 60372 435882 60424 435888
rect 60372 391332 60424 391338
rect 60372 391274 60424 391280
rect 59268 389904 59320 389910
rect 59268 389846 59320 389852
rect 59176 388068 59228 388074
rect 59176 388010 59228 388016
rect 59084 385756 59136 385762
rect 59084 385698 59136 385704
rect 58992 377460 59044 377466
rect 58992 377402 59044 377408
rect 58900 339312 58952 339318
rect 58900 339254 58952 339260
rect 57888 337748 57940 337754
rect 57888 337690 57940 337696
rect 57796 294704 57848 294710
rect 57796 294646 57848 294652
rect 57796 249824 57848 249830
rect 57796 249766 57848 249772
rect 57704 245608 57756 245614
rect 57704 245550 57756 245556
rect 57520 217320 57572 217326
rect 57520 217262 57572 217268
rect 56508 193928 56560 193934
rect 56508 193870 56560 193876
rect 57808 186969 57836 249766
rect 57900 237250 57928 337690
rect 59096 336598 59124 385698
rect 59188 383654 59216 388010
rect 59188 383626 59308 383654
rect 59176 377460 59228 377466
rect 59176 377402 59228 377408
rect 59188 376038 59216 377402
rect 59176 376032 59228 376038
rect 59176 375974 59228 375980
rect 59176 360868 59228 360874
rect 59176 360810 59228 360816
rect 59188 359514 59216 360810
rect 59176 359508 59228 359514
rect 59176 359450 59228 359456
rect 59084 336592 59136 336598
rect 59084 336534 59136 336540
rect 58992 258120 59044 258126
rect 58992 258062 59044 258068
rect 57888 237244 57940 237250
rect 57888 237186 57940 237192
rect 57794 186960 57850 186969
rect 57794 186895 57850 186904
rect 59004 185706 59032 258062
rect 59084 247104 59136 247110
rect 59084 247046 59136 247052
rect 58992 185700 59044 185706
rect 58992 185642 59044 185648
rect 59096 182918 59124 247046
rect 59188 238678 59216 359450
rect 59280 255270 59308 383626
rect 60280 378820 60332 378826
rect 60280 378762 60332 378768
rect 60292 335354 60320 378762
rect 60384 337754 60412 391274
rect 60476 367130 60504 464986
rect 60568 442898 60596 542438
rect 60660 445942 60688 546450
rect 61764 538898 61792 583782
rect 61844 572756 61896 572762
rect 61844 572698 61896 572704
rect 61752 538892 61804 538898
rect 61752 538834 61804 538840
rect 61752 478916 61804 478922
rect 61752 478858 61804 478864
rect 61382 463584 61438 463593
rect 61382 463519 61438 463528
rect 61396 462369 61424 463519
rect 61382 462360 61438 462369
rect 61382 462295 61438 462304
rect 60648 445936 60700 445942
rect 60648 445878 60700 445884
rect 60738 442912 60794 442921
rect 60568 442870 60738 442898
rect 60738 442847 60794 442856
rect 60556 391536 60608 391542
rect 60556 391478 60608 391484
rect 60464 367124 60516 367130
rect 60464 367066 60516 367072
rect 60372 337748 60424 337754
rect 60372 337690 60424 337696
rect 60568 336462 60596 391478
rect 61396 367062 61424 462295
rect 61764 386374 61792 478858
rect 61856 474366 61884 572698
rect 61936 563168 61988 563174
rect 61936 563110 61988 563116
rect 61844 474360 61896 474366
rect 61844 474302 61896 474308
rect 61948 465050 61976 563110
rect 62040 563038 62068 700266
rect 68836 596828 68888 596834
rect 68836 596770 68888 596776
rect 68468 589960 68520 589966
rect 68468 589902 68520 589908
rect 67638 581360 67694 581369
rect 67638 581295 67640 581304
rect 67692 581295 67694 581304
rect 67640 581266 67692 581272
rect 67914 580680 67970 580689
rect 67914 580615 67970 580624
rect 67928 580310 67956 580615
rect 67916 580304 67968 580310
rect 67916 580246 67968 580252
rect 67362 579184 67418 579193
rect 67362 579119 67418 579128
rect 63224 576904 63276 576910
rect 63224 576846 63276 576852
rect 62028 563032 62080 563038
rect 62028 562974 62080 562980
rect 62764 557592 62816 557598
rect 62764 557534 62816 557540
rect 62028 541000 62080 541006
rect 62028 540942 62080 540948
rect 61936 465044 61988 465050
rect 61936 464986 61988 464992
rect 61936 448520 61988 448526
rect 61936 448462 61988 448468
rect 61752 386368 61804 386374
rect 61752 386310 61804 386316
rect 61660 385892 61712 385898
rect 61660 385834 61712 385840
rect 61476 367804 61528 367810
rect 61476 367746 61528 367752
rect 61384 367056 61436 367062
rect 61384 366998 61436 367004
rect 61488 366382 61516 367746
rect 61476 366376 61528 366382
rect 61476 366318 61528 366324
rect 60740 362228 60792 362234
rect 60740 362170 60792 362176
rect 60752 361690 60780 362170
rect 60740 361684 60792 361690
rect 60740 361626 60792 361632
rect 61488 359582 61516 366318
rect 61672 364334 61700 385834
rect 61580 364306 61700 364334
rect 61476 359576 61528 359582
rect 61476 359518 61528 359524
rect 60648 356720 60700 356726
rect 60648 356662 60700 356668
rect 60660 356182 60688 356662
rect 60648 356176 60700 356182
rect 60648 356118 60700 356124
rect 60556 336456 60608 336462
rect 60556 336398 60608 336404
rect 60292 335326 60596 335354
rect 60568 335170 60596 335326
rect 60556 335164 60608 335170
rect 60556 335106 60608 335112
rect 60464 297492 60516 297498
rect 60464 297434 60516 297440
rect 60280 260908 60332 260914
rect 60280 260850 60332 260856
rect 59268 255264 59320 255270
rect 59268 255206 59320 255212
rect 59176 238672 59228 238678
rect 59176 238614 59228 238620
rect 59084 182912 59136 182918
rect 59084 182854 59136 182860
rect 60292 181490 60320 260850
rect 60476 260846 60504 297434
rect 60464 260840 60516 260846
rect 60464 260782 60516 260788
rect 60372 241528 60424 241534
rect 60372 241470 60424 241476
rect 60384 218754 60412 241470
rect 60568 238542 60596 335106
rect 60556 238536 60608 238542
rect 60556 238478 60608 238484
rect 60660 237182 60688 356118
rect 61580 354674 61608 364306
rect 61752 361684 61804 361690
rect 61752 361626 61804 361632
rect 61580 354646 61700 354674
rect 61672 339590 61700 354646
rect 61660 339584 61712 339590
rect 61660 339526 61712 339532
rect 61384 337952 61436 337958
rect 61382 337920 61384 337929
rect 61436 337920 61438 337929
rect 61382 337855 61438 337864
rect 61764 333266 61792 361626
rect 61844 359576 61896 359582
rect 61844 359518 61896 359524
rect 61752 333260 61804 333266
rect 61752 333202 61804 333208
rect 61856 298790 61884 359518
rect 61948 348430 61976 448462
rect 62040 440366 62068 540942
rect 62776 459610 62804 557534
rect 63236 480078 63264 576846
rect 64604 574184 64656 574190
rect 64604 574126 64656 574132
rect 63408 549364 63460 549370
rect 63408 549306 63460 549312
rect 63316 546576 63368 546582
rect 63316 546518 63368 546524
rect 63224 480072 63276 480078
rect 63224 480014 63276 480020
rect 63236 478922 63264 480014
rect 63224 478916 63276 478922
rect 63224 478858 63276 478864
rect 63222 467800 63278 467809
rect 63222 467735 63278 467744
rect 62764 459604 62816 459610
rect 62764 459546 62816 459552
rect 62764 449948 62816 449954
rect 62764 449890 62816 449896
rect 62028 440360 62080 440366
rect 62028 440302 62080 440308
rect 62026 401704 62082 401713
rect 62026 401639 62082 401648
rect 62040 382226 62068 401639
rect 62028 382220 62080 382226
rect 62028 382162 62080 382168
rect 62776 352578 62804 449890
rect 63236 371278 63264 467735
rect 63328 448526 63356 546518
rect 63420 449274 63448 549306
rect 64144 482996 64196 483002
rect 64144 482938 64196 482944
rect 63408 449268 63460 449274
rect 63408 449210 63460 449216
rect 63316 448520 63368 448526
rect 63316 448462 63368 448468
rect 63314 447808 63370 447817
rect 63314 447743 63370 447752
rect 63224 371272 63276 371278
rect 63224 371214 63276 371220
rect 62856 357468 62908 357474
rect 62856 357410 62908 357416
rect 62764 352572 62816 352578
rect 62764 352514 62816 352520
rect 61936 348424 61988 348430
rect 61936 348366 61988 348372
rect 62868 338774 62896 357410
rect 63328 349858 63356 447743
rect 64156 436762 64184 482938
rect 64616 477465 64644 574126
rect 64696 572824 64748 572830
rect 64696 572766 64748 572772
rect 64602 477456 64658 477465
rect 64602 477391 64658 477400
rect 64708 475046 64736 572766
rect 66168 571600 66220 571606
rect 66168 571542 66220 571548
rect 64788 568676 64840 568682
rect 64788 568618 64840 568624
rect 64696 475040 64748 475046
rect 64696 474982 64748 474988
rect 64512 445936 64564 445942
rect 64512 445878 64564 445884
rect 64144 436756 64196 436762
rect 64144 436698 64196 436704
rect 64420 380860 64472 380866
rect 64420 380802 64472 380808
rect 63408 367124 63460 367130
rect 63408 367066 63460 367072
rect 63316 349852 63368 349858
rect 63316 349794 63368 349800
rect 63316 345704 63368 345710
rect 63316 345646 63368 345652
rect 63328 345098 63356 345646
rect 63316 345092 63368 345098
rect 63316 345034 63368 345040
rect 62856 338768 62908 338774
rect 62856 338710 62908 338716
rect 62028 334620 62080 334626
rect 62028 334562 62080 334568
rect 61936 300212 61988 300218
rect 61936 300154 61988 300160
rect 61844 298784 61896 298790
rect 61844 298726 61896 298732
rect 61844 274780 61896 274786
rect 61844 274722 61896 274728
rect 60924 253972 60976 253978
rect 60924 253914 60976 253920
rect 60936 253881 60964 253914
rect 60922 253872 60978 253881
rect 60922 253807 60978 253816
rect 61660 244656 61712 244662
rect 61660 244598 61712 244604
rect 60648 237176 60700 237182
rect 60648 237118 60700 237124
rect 60372 218748 60424 218754
rect 60372 218690 60424 218696
rect 61672 185774 61700 244598
rect 61752 240168 61804 240174
rect 61752 240110 61804 240116
rect 61764 213314 61792 240110
rect 61856 222902 61884 274722
rect 61948 263566 61976 300154
rect 61936 263560 61988 263566
rect 61936 263502 61988 263508
rect 61936 260976 61988 260982
rect 61936 260918 61988 260924
rect 61844 222896 61896 222902
rect 61844 222838 61896 222844
rect 61752 213308 61804 213314
rect 61752 213250 61804 213256
rect 61948 192506 61976 260918
rect 62040 242894 62068 334562
rect 63328 331974 63356 345034
rect 63316 331968 63368 331974
rect 63316 331910 63368 331916
rect 63224 256760 63276 256766
rect 63224 256702 63276 256708
rect 63132 244316 63184 244322
rect 63132 244258 63184 244264
rect 62028 242888 62080 242894
rect 62028 242830 62080 242836
rect 63144 196761 63172 244258
rect 63236 239426 63264 256702
rect 63316 252612 63368 252618
rect 63316 252554 63368 252560
rect 63328 239494 63356 252554
rect 63316 239488 63368 239494
rect 63316 239430 63368 239436
rect 63224 239420 63276 239426
rect 63224 239362 63276 239368
rect 63130 196752 63186 196761
rect 63130 196687 63186 196696
rect 61936 192500 61988 192506
rect 61936 192442 61988 192448
rect 61660 185768 61712 185774
rect 61660 185710 61712 185716
rect 60280 181484 60332 181490
rect 60280 181426 60332 181432
rect 60648 124228 60700 124234
rect 60648 124170 60700 124176
rect 60660 93673 60688 124170
rect 62028 122868 62080 122874
rect 62028 122810 62080 122816
rect 60646 93664 60702 93673
rect 60646 93599 60702 93608
rect 62040 89729 62068 122810
rect 62026 89720 62082 89729
rect 62026 89655 62082 89664
rect 56598 73808 56654 73817
rect 56598 73743 56654 73752
rect 53930 24848 53986 24857
rect 53930 24783 53986 24792
rect 55126 24848 55182 24857
rect 55126 24783 55182 24792
rect 53944 24177 53972 24783
rect 53930 24168 53986 24177
rect 53930 24103 53986 24112
rect 55220 17264 55272 17270
rect 55220 17206 55272 17212
rect 55232 16574 55260 17206
rect 56612 16574 56640 73743
rect 60740 61464 60792 61470
rect 60740 61406 60792 61412
rect 57980 28348 58032 28354
rect 57980 28290 58032 28296
rect 57992 16574 58020 28290
rect 60752 16574 60780 61406
rect 63420 22846 63448 367066
rect 63500 355360 63552 355366
rect 63498 355328 63500 355337
rect 63552 355328 63554 355337
rect 63498 355263 63554 355272
rect 63500 343732 63552 343738
rect 63500 343674 63552 343680
rect 63512 342922 63540 343674
rect 63500 342916 63552 342922
rect 63500 342858 63552 342864
rect 63498 72448 63554 72457
rect 63498 72383 63554 72392
rect 63408 22840 63460 22846
rect 63408 22782 63460 22788
rect 63512 16574 63540 72383
rect 64432 71058 64460 380802
rect 64524 347070 64552 445878
rect 64708 380798 64736 474982
rect 64800 470558 64828 568618
rect 66076 567248 66128 567254
rect 66076 567190 66128 567196
rect 65984 564528 66036 564534
rect 65984 564470 66036 564476
rect 65892 484628 65944 484634
rect 65892 484570 65944 484576
rect 64788 470552 64840 470558
rect 64788 470494 64840 470500
rect 64788 468172 64840 468178
rect 64788 468114 64840 468120
rect 64800 398857 64828 468114
rect 65524 445800 65576 445806
rect 65524 445742 65576 445748
rect 64786 398848 64842 398857
rect 64786 398783 64842 398792
rect 64696 380792 64748 380798
rect 64696 380734 64748 380740
rect 64696 375352 64748 375358
rect 64696 375294 64748 375300
rect 64604 351212 64656 351218
rect 64604 351154 64656 351160
rect 64512 347064 64564 347070
rect 64512 347006 64564 347012
rect 64616 73846 64644 351154
rect 64708 75206 64736 375294
rect 64800 372570 64828 398783
rect 64788 372564 64840 372570
rect 64788 372506 64840 372512
rect 65536 346458 65564 445742
rect 65904 438258 65932 484570
rect 65996 465610 66024 564470
rect 66088 468178 66116 567190
rect 66180 472054 66208 571542
rect 67178 568712 67234 568721
rect 67178 568647 67234 568656
rect 66168 472048 66220 472054
rect 66168 471990 66220 471996
rect 66904 470552 66956 470558
rect 66904 470494 66956 470500
rect 66076 468172 66128 468178
rect 66076 468114 66128 468120
rect 65996 465582 66208 465610
rect 66180 465458 66208 465582
rect 66168 465452 66220 465458
rect 66168 465394 66220 465400
rect 66074 461408 66130 461417
rect 66074 461343 66130 461352
rect 66088 461009 66116 461343
rect 66074 461000 66130 461009
rect 66074 460935 66130 460944
rect 65982 440328 66038 440337
rect 65982 440263 65984 440272
rect 66036 440263 66038 440272
rect 65984 440234 66036 440240
rect 65892 438252 65944 438258
rect 65892 438194 65944 438200
rect 66088 402974 66116 460935
rect 65996 402946 66116 402974
rect 65996 397526 66024 402946
rect 65984 397520 66036 397526
rect 65984 397462 66036 397468
rect 65996 393314 66024 397462
rect 66076 394868 66128 394874
rect 66076 394810 66128 394816
rect 66088 394194 66116 394810
rect 66076 394188 66128 394194
rect 66076 394130 66128 394136
rect 65996 393286 66116 393314
rect 66088 376718 66116 393286
rect 66076 376712 66128 376718
rect 66076 376654 66128 376660
rect 66180 369170 66208 465394
rect 66916 375358 66944 470494
rect 67192 469878 67220 568647
rect 67272 549160 67324 549166
rect 67272 549102 67324 549108
rect 67180 469872 67232 469878
rect 67180 469814 67232 469820
rect 67284 459513 67312 549102
rect 67376 480593 67404 579119
rect 67638 578504 67694 578513
rect 67638 578439 67694 578448
rect 67652 578338 67680 578439
rect 67640 578332 67692 578338
rect 67640 578274 67692 578280
rect 67638 577824 67694 577833
rect 67638 577759 67694 577768
rect 67652 576910 67680 577759
rect 67640 576904 67692 576910
rect 67640 576846 67692 576852
rect 67638 575784 67694 575793
rect 67638 575719 67694 575728
rect 67652 575550 67680 575719
rect 67640 575544 67692 575550
rect 67640 575486 67692 575492
rect 67730 575104 67786 575113
rect 67730 575039 67786 575048
rect 67638 574424 67694 574433
rect 67638 574359 67694 574368
rect 67652 574122 67680 574359
rect 67744 574190 67772 575039
rect 67732 574184 67784 574190
rect 67732 574126 67784 574132
rect 67640 574116 67692 574122
rect 67640 574058 67692 574064
rect 67730 573472 67786 573481
rect 67730 573407 67786 573416
rect 67744 572830 67772 573407
rect 67732 572824 67784 572830
rect 67638 572792 67694 572801
rect 67732 572766 67784 572772
rect 67638 572727 67640 572736
rect 67692 572727 67694 572736
rect 67640 572698 67692 572704
rect 68480 571713 68508 589902
rect 68848 586514 68876 596770
rect 68756 586486 68876 586514
rect 68756 586378 68784 586486
rect 68572 586350 68784 586378
rect 68572 580689 68600 586350
rect 68940 582570 68968 702442
rect 69020 696992 69072 696998
rect 69020 696934 69072 696940
rect 68664 582542 68968 582570
rect 68558 580680 68614 580689
rect 68558 580615 68614 580624
rect 68664 571849 68692 582542
rect 68744 582412 68796 582418
rect 68744 582354 68796 582360
rect 68650 571840 68706 571849
rect 68650 571775 68706 571784
rect 68282 571704 68338 571713
rect 68282 571639 68338 571648
rect 68466 571704 68522 571713
rect 68466 571639 68522 571648
rect 68296 571606 68324 571639
rect 68284 571600 68336 571606
rect 68284 571542 68336 571548
rect 67638 570072 67694 570081
rect 67638 570007 67694 570016
rect 67652 569974 67680 570007
rect 67640 569968 67692 569974
rect 67640 569910 67692 569916
rect 67638 568984 67694 568993
rect 67638 568919 67694 568928
rect 67652 568682 67680 568919
rect 67640 568676 67692 568682
rect 67640 568618 67692 568624
rect 67546 567624 67602 567633
rect 67546 567559 67602 567568
rect 67362 480584 67418 480593
rect 67362 480519 67418 480528
rect 67456 471980 67508 471986
rect 67456 471922 67508 471928
rect 67270 459504 67326 459513
rect 67270 459439 67326 459448
rect 67284 458862 67312 459439
rect 67272 458856 67324 458862
rect 67272 458798 67324 458804
rect 67008 451926 67036 451957
rect 66996 451920 67048 451926
rect 66994 451888 66996 451897
rect 67048 451888 67050 451897
rect 66994 451823 67050 451832
rect 67008 419490 67036 451823
rect 66996 419484 67048 419490
rect 66996 419426 67048 419432
rect 67364 419484 67416 419490
rect 67364 419426 67416 419432
rect 67376 418810 67404 419426
rect 67364 418804 67416 418810
rect 67364 418746 67416 418752
rect 67468 380866 67496 471922
rect 67560 469010 67588 567559
rect 67640 567248 67692 567254
rect 67638 567216 67640 567225
rect 67692 567216 67694 567225
rect 67638 567151 67694 567160
rect 67638 564904 67694 564913
rect 67638 564839 67694 564848
rect 67652 564466 67680 564839
rect 67732 564528 67784 564534
rect 67730 564496 67732 564505
rect 67784 564496 67786 564505
rect 67640 564460 67692 564466
rect 67730 564431 67786 564440
rect 67640 564402 67692 564408
rect 67730 564224 67786 564233
rect 67730 564159 67786 564168
rect 67638 563680 67694 563689
rect 67638 563615 67694 563624
rect 67652 563174 67680 563615
rect 67640 563168 67692 563174
rect 67640 563110 67692 563116
rect 67744 563106 67772 564159
rect 67732 563100 67784 563106
rect 67732 563042 67784 563048
rect 67640 563032 67692 563038
rect 67638 563000 67640 563009
rect 67692 563000 67694 563009
rect 67638 562935 67694 562944
rect 67638 560416 67694 560425
rect 67638 560351 67694 560360
rect 67652 560318 67680 560351
rect 67640 560312 67692 560318
rect 67640 560254 67692 560260
rect 67638 559464 67694 559473
rect 67638 559399 67694 559408
rect 67652 558958 67680 559399
rect 67640 558952 67692 558958
rect 67640 558894 67692 558900
rect 68374 558920 68430 558929
rect 68374 558855 68430 558864
rect 67640 557592 67692 557598
rect 67638 557560 67640 557569
rect 67692 557560 67694 557569
rect 67638 557495 67694 557504
rect 67730 556744 67786 556753
rect 67730 556679 67786 556688
rect 67744 556306 67772 556679
rect 67732 556300 67784 556306
rect 67732 556242 67784 556248
rect 67640 556232 67692 556238
rect 67638 556200 67640 556209
rect 67692 556200 67694 556209
rect 67638 556135 67694 556144
rect 67732 556164 67784 556170
rect 67732 556106 67784 556112
rect 67638 555384 67694 555393
rect 67638 555319 67694 555328
rect 67652 554810 67680 555319
rect 67744 554849 67772 556106
rect 67730 554840 67786 554849
rect 67640 554804 67692 554810
rect 67730 554775 67786 554784
rect 67640 554746 67692 554752
rect 67638 553480 67694 553489
rect 67638 553415 67640 553424
rect 67692 553415 67694 553424
rect 67640 553386 67692 553392
rect 67638 552120 67694 552129
rect 67638 552055 67640 552064
rect 67692 552055 67694 552064
rect 67640 552026 67692 552032
rect 67638 551304 67694 551313
rect 67638 551239 67694 551248
rect 67652 550662 67680 551239
rect 68282 550760 68338 550769
rect 68282 550695 68338 550704
rect 67640 550656 67692 550662
rect 67640 550598 67692 550604
rect 67730 549944 67786 549953
rect 67730 549879 67786 549888
rect 67638 549400 67694 549409
rect 67638 549335 67640 549344
rect 67692 549335 67694 549344
rect 67640 549306 67692 549312
rect 67744 549302 67772 549879
rect 67732 549296 67784 549302
rect 67732 549238 67784 549244
rect 67638 548584 67694 548593
rect 67638 548519 67694 548528
rect 67652 547942 67680 548519
rect 67640 547936 67692 547942
rect 67640 547878 67692 547884
rect 67730 547224 67786 547233
rect 67730 547159 67786 547168
rect 67744 546582 67772 547159
rect 67732 546576 67784 546582
rect 67638 546544 67694 546553
rect 67732 546518 67784 546524
rect 67638 546479 67640 546488
rect 67692 546479 67694 546488
rect 67640 546450 67692 546456
rect 67730 544504 67786 544513
rect 67730 544439 67786 544448
rect 67744 543862 67772 544439
rect 67732 543856 67784 543862
rect 67638 543824 67694 543833
rect 67732 543798 67784 543804
rect 67638 543759 67640 543768
rect 67692 543759 67694 543768
rect 67640 543730 67692 543736
rect 67638 542600 67694 542609
rect 67638 542535 67694 542544
rect 67652 542502 67680 542535
rect 67640 542496 67692 542502
rect 67640 542438 67692 542444
rect 67638 541240 67694 541249
rect 67638 541175 67694 541184
rect 67652 541006 67680 541175
rect 67640 541000 67692 541006
rect 67640 540942 67692 540948
rect 67638 540152 67694 540161
rect 67638 540087 67694 540096
rect 67652 539646 67680 540087
rect 67640 539640 67692 539646
rect 67640 539582 67692 539588
rect 68008 493400 68060 493406
rect 68008 493342 68060 493348
rect 68020 491706 68048 493342
rect 68008 491700 68060 491706
rect 68008 491642 68060 491648
rect 67730 488064 67786 488073
rect 67730 487999 67786 488008
rect 67638 487928 67694 487937
rect 67638 487863 67694 487872
rect 67652 487830 67680 487863
rect 67640 487824 67692 487830
rect 67640 487766 67692 487772
rect 67744 487218 67772 487999
rect 67732 487212 67784 487218
rect 67732 487154 67784 487160
rect 67638 485888 67694 485897
rect 67638 485823 67640 485832
rect 67692 485823 67694 485832
rect 67640 485794 67692 485800
rect 67638 485208 67694 485217
rect 67638 485143 67694 485152
rect 67652 484430 67680 485143
rect 67640 484424 67692 484430
rect 67640 484366 67692 484372
rect 67638 483712 67694 483721
rect 67638 483647 67694 483656
rect 67652 483070 67680 483647
rect 67640 483064 67692 483070
rect 67640 483006 67692 483012
rect 68100 482928 68152 482934
rect 68100 482870 68152 482876
rect 68112 482497 68140 482870
rect 68098 482488 68154 482497
rect 68098 482423 68154 482432
rect 67638 480176 67694 480185
rect 67638 480111 67640 480120
rect 67692 480111 67694 480120
rect 67640 480082 67692 480088
rect 67732 480072 67784 480078
rect 67732 480014 67784 480020
rect 67744 479913 67772 480014
rect 67730 479904 67786 479913
rect 67730 479839 67786 479848
rect 67730 477456 67786 477465
rect 67730 477391 67786 477400
rect 67638 476368 67694 476377
rect 67638 476303 67694 476312
rect 67652 476134 67680 476303
rect 67744 476241 67772 477391
rect 67730 476232 67786 476241
rect 67730 476167 67786 476176
rect 67640 476128 67692 476134
rect 67640 476070 67692 476076
rect 67638 475688 67694 475697
rect 67638 475623 67694 475632
rect 67652 475386 67680 475623
rect 67640 475380 67692 475386
rect 67640 475322 67692 475328
rect 67640 475040 67692 475046
rect 67638 475008 67640 475017
rect 67692 475008 67694 475017
rect 67638 474943 67694 474952
rect 67640 474360 67692 474366
rect 67638 474328 67640 474337
rect 67692 474328 67694 474337
rect 67694 474286 67772 474314
rect 67638 474263 67694 474272
rect 67638 472288 67694 472297
rect 67638 472223 67694 472232
rect 67652 472054 67680 472223
rect 67640 472048 67692 472054
rect 67640 471990 67692 471996
rect 67744 471986 67772 474286
rect 67732 471980 67784 471986
rect 67732 471922 67784 471928
rect 67638 470928 67694 470937
rect 67638 470863 67694 470872
rect 67652 470626 67680 470863
rect 67640 470620 67692 470626
rect 67640 470562 67692 470568
rect 67732 470552 67784 470558
rect 67732 470494 67784 470500
rect 67744 470393 67772 470494
rect 67730 470384 67786 470393
rect 67730 470319 67786 470328
rect 67640 469872 67692 469878
rect 67640 469814 67692 469820
rect 67652 469713 67680 469814
rect 67638 469704 67694 469713
rect 67638 469639 67694 469648
rect 67638 469024 67694 469033
rect 67560 468982 67638 469010
rect 67638 468959 67694 468968
rect 67638 468208 67694 468217
rect 67638 468143 67640 468152
rect 67692 468143 67694 468152
rect 67640 468114 67692 468120
rect 67640 465724 67692 465730
rect 67640 465666 67692 465672
rect 67652 465633 67680 465666
rect 67638 465624 67694 465633
rect 67638 465559 67694 465568
rect 67638 465488 67694 465497
rect 67638 465423 67640 465432
rect 67692 465423 67694 465432
rect 67640 465394 67692 465400
rect 67732 465044 67784 465050
rect 67732 464986 67784 464992
rect 67638 464808 67694 464817
rect 67638 464743 67694 464752
rect 67652 464370 67680 464743
rect 67640 464364 67692 464370
rect 67640 464306 67692 464312
rect 67744 464273 67772 464986
rect 67730 464264 67786 464273
rect 67730 464199 67786 464208
rect 67640 463004 67692 463010
rect 67640 462946 67692 462952
rect 67652 462913 67680 462946
rect 67638 462904 67694 462913
rect 67638 462839 67694 462848
rect 67638 460728 67694 460737
rect 67638 460663 67694 460672
rect 67652 460290 67680 460663
rect 67640 460284 67692 460290
rect 67640 460226 67692 460232
rect 67732 460216 67784 460222
rect 67730 460184 67732 460193
rect 67784 460184 67786 460193
rect 67730 460119 67786 460128
rect 67640 459536 67692 459542
rect 67640 459478 67692 459484
rect 67652 458833 67680 459478
rect 67638 458824 67694 458833
rect 67638 458759 67694 458768
rect 68100 458176 68152 458182
rect 68100 458118 68152 458124
rect 68112 458017 68140 458118
rect 68098 458008 68154 458017
rect 68098 457943 68154 457952
rect 67640 457496 67692 457502
rect 67638 457464 67640 457473
rect 67692 457464 67694 457473
rect 67638 457399 67694 457408
rect 67638 455968 67694 455977
rect 67638 455903 67694 455912
rect 67652 455462 67680 455903
rect 67640 455456 67692 455462
rect 67640 455398 67692 455404
rect 67732 454708 67784 454714
rect 67732 454650 67784 454656
rect 67638 454608 67694 454617
rect 67638 454543 67694 454552
rect 67652 454102 67680 454543
rect 67640 454096 67692 454102
rect 67640 454038 67692 454044
rect 67744 453937 67772 454650
rect 67730 453928 67786 453937
rect 67730 453863 67786 453872
rect 67640 453348 67692 453354
rect 67640 453290 67692 453296
rect 67652 453257 67680 453290
rect 67638 453248 67694 453257
rect 67638 453183 67694 453192
rect 68296 452674 68324 550695
rect 68388 549166 68416 558855
rect 68376 549160 68428 549166
rect 68376 549102 68428 549108
rect 68756 545873 68784 582354
rect 68834 576464 68890 576473
rect 68834 576399 68890 576408
rect 68742 545864 68798 545873
rect 68742 545799 68798 545808
rect 68756 545766 68784 545799
rect 68744 545760 68796 545766
rect 68744 545702 68796 545708
rect 68742 484664 68798 484673
rect 68742 484599 68744 484608
rect 68796 484599 68798 484608
rect 68744 484570 68796 484576
rect 68558 481128 68614 481137
rect 68558 481063 68614 481072
rect 68572 480282 68600 481063
rect 68560 480276 68612 480282
rect 68560 480218 68612 480224
rect 68848 477057 68876 576399
rect 68926 543280 68982 543289
rect 69032 543266 69060 696934
rect 71792 596174 71820 702986
rect 75184 702840 75236 702846
rect 75184 702782 75236 702788
rect 71792 596146 71912 596174
rect 69112 585812 69164 585818
rect 69112 585754 69164 585760
rect 69124 558929 69152 585754
rect 71778 583944 71834 583953
rect 71778 583879 71834 583888
rect 69204 583772 69256 583778
rect 69204 583714 69256 583720
rect 69110 558920 69166 558929
rect 69110 558855 69166 558864
rect 69110 554024 69166 554033
rect 69110 553959 69166 553968
rect 68982 543238 69060 543266
rect 68926 543215 68982 543224
rect 68940 542434 68968 543215
rect 68928 542428 68980 542434
rect 68928 542370 68980 542376
rect 68926 541784 68982 541793
rect 68926 541719 68982 541728
rect 68940 525774 68968 541719
rect 68928 525768 68980 525774
rect 68928 525710 68980 525716
rect 68374 477048 68430 477057
rect 68374 476983 68430 476992
rect 68834 477048 68890 477057
rect 68834 476983 68890 476992
rect 67732 452668 67784 452674
rect 67732 452610 67784 452616
rect 68284 452668 68336 452674
rect 68284 452610 68336 452616
rect 67744 451353 67772 452610
rect 67730 451344 67786 451353
rect 67730 451279 67786 451288
rect 67638 449984 67694 449993
rect 67638 449919 67640 449928
rect 67692 449919 67694 449928
rect 67640 449890 67692 449896
rect 67730 449304 67786 449313
rect 67730 449239 67732 449248
rect 67784 449239 67786 449248
rect 68282 449304 68338 449313
rect 68282 449239 68338 449248
rect 67732 449210 67784 449216
rect 67640 449200 67692 449206
rect 67638 449168 67640 449177
rect 67692 449168 67694 449177
rect 67638 449103 67694 449112
rect 67640 448520 67692 448526
rect 67640 448462 67692 448468
rect 67652 447273 67680 448462
rect 67638 447264 67694 447273
rect 67638 447199 67694 447208
rect 67638 446448 67694 446457
rect 67638 446383 67694 446392
rect 67652 445942 67680 446383
rect 67640 445936 67692 445942
rect 67640 445878 67692 445884
rect 67730 445904 67786 445913
rect 67730 445839 67786 445848
rect 67744 445806 67772 445839
rect 67732 445800 67784 445806
rect 67732 445742 67784 445748
rect 67638 445088 67694 445097
rect 67638 445023 67640 445032
rect 67692 445023 67694 445032
rect 67640 444994 67692 445000
rect 67640 444372 67692 444378
rect 67640 444314 67692 444320
rect 67652 443873 67680 444314
rect 67730 444272 67786 444281
rect 67730 444207 67786 444216
rect 67638 443864 67694 443873
rect 67638 443799 67694 443808
rect 67744 443018 67772 444207
rect 67732 443012 67784 443018
rect 67732 442954 67784 442960
rect 67640 442944 67692 442950
rect 67640 442886 67692 442892
rect 67730 442912 67786 442921
rect 67652 442513 67680 442886
rect 67730 442847 67786 442856
rect 67638 442504 67694 442513
rect 67638 442439 67694 442448
rect 67744 441697 67772 442847
rect 67730 441688 67786 441697
rect 67730 441623 67786 441632
rect 67730 441144 67786 441153
rect 67730 441079 67786 441088
rect 67744 440366 67772 441079
rect 67548 440360 67600 440366
rect 67732 440360 67784 440366
rect 67548 440302 67600 440308
rect 67638 440328 67694 440337
rect 67456 380860 67508 380866
rect 67456 380802 67508 380808
rect 67468 379953 67496 380802
rect 67454 379944 67510 379953
rect 67454 379879 67510 379888
rect 66904 375352 66956 375358
rect 66904 375294 66956 375300
rect 66904 373992 66956 373998
rect 66904 373934 66956 373940
rect 66168 369164 66220 369170
rect 66168 369106 66220 369112
rect 65616 360256 65668 360262
rect 65616 360198 65668 360204
rect 65524 346452 65576 346458
rect 65524 346394 65576 346400
rect 65628 307154 65656 360198
rect 66076 345024 66128 345030
rect 66076 344966 66128 344972
rect 65984 340944 66036 340950
rect 65984 340886 66036 340892
rect 65616 307148 65668 307154
rect 65616 307090 65668 307096
rect 65996 302938 66024 340886
rect 66088 338842 66116 344966
rect 66076 338836 66128 338842
rect 66076 338778 66128 338784
rect 66180 320793 66208 369106
rect 66916 322250 66944 373934
rect 67456 371272 67508 371278
rect 67456 371214 67508 371220
rect 66996 353252 67048 353258
rect 66996 353194 67048 353200
rect 67008 337414 67036 353194
rect 66996 337408 67048 337414
rect 66996 337350 67048 337356
rect 67468 331906 67496 371214
rect 67560 341601 67588 440302
rect 67732 440302 67784 440308
rect 67638 440263 67694 440272
rect 67652 439521 67680 440263
rect 67638 439512 67694 439521
rect 67638 439447 67694 439456
rect 67730 382528 67786 382537
rect 67730 382463 67786 382472
rect 67744 382294 67772 382463
rect 67732 382288 67784 382294
rect 67732 382230 67784 382236
rect 67640 382220 67692 382226
rect 67640 382162 67692 382168
rect 67652 382129 67680 382162
rect 67638 382120 67694 382129
rect 67638 382055 67694 382064
rect 68008 380792 68060 380798
rect 67638 380760 67694 380769
rect 68008 380734 68060 380740
rect 67638 380695 67640 380704
rect 67692 380695 67694 380704
rect 67640 380666 67692 380672
rect 68020 380361 68048 380734
rect 68006 380352 68062 380361
rect 68006 380287 68062 380296
rect 67638 378312 67694 378321
rect 67638 378247 67694 378256
rect 67652 378214 67680 378247
rect 67640 378208 67692 378214
rect 67640 378150 67692 378156
rect 67640 377460 67692 377466
rect 67640 377402 67692 377408
rect 67652 377369 67680 377402
rect 67638 377360 67694 377369
rect 67638 377295 67694 377304
rect 67640 375352 67692 375358
rect 67640 375294 67692 375300
rect 67652 375193 67680 375294
rect 67638 375184 67694 375193
rect 67638 375119 67694 375128
rect 67730 374232 67786 374241
rect 67730 374167 67786 374176
rect 67744 374066 67772 374167
rect 67732 374060 67784 374066
rect 67732 374002 67784 374008
rect 67640 372564 67692 372570
rect 67640 372506 67692 372512
rect 67652 372473 67680 372506
rect 67638 372464 67694 372473
rect 67638 372399 67694 372408
rect 67638 371512 67694 371521
rect 67638 371447 67694 371456
rect 67652 371278 67680 371447
rect 67640 371272 67692 371278
rect 67640 371214 67692 371220
rect 67640 369844 67692 369850
rect 67640 369786 67692 369792
rect 67652 369073 67680 369786
rect 67730 369200 67786 369209
rect 67730 369135 67732 369144
rect 67784 369135 67786 369144
rect 67732 369106 67784 369112
rect 67638 369064 67694 369073
rect 67638 368999 67694 369008
rect 67638 367160 67694 367169
rect 67638 367095 67640 367104
rect 67692 367095 67694 367104
rect 67640 367066 67692 367072
rect 67732 367056 67784 367062
rect 67732 366998 67784 367004
rect 67638 366480 67694 366489
rect 67638 366415 67694 366424
rect 67652 366382 67680 366415
rect 67640 366376 67692 366382
rect 67744 366353 67772 366998
rect 67640 366318 67692 366324
rect 67730 366344 67786 366353
rect 67730 366279 67786 366288
rect 67638 363760 67694 363769
rect 67638 363695 67640 363704
rect 67692 363695 67694 363704
rect 67640 363666 67692 363672
rect 67732 363656 67784 363662
rect 67730 363624 67732 363633
rect 67784 363624 67786 363633
rect 67730 363559 67786 363568
rect 67638 362128 67694 362137
rect 67638 362063 67694 362072
rect 67652 361690 67680 362063
rect 67640 361684 67692 361690
rect 67640 361626 67692 361632
rect 67638 361040 67694 361049
rect 67638 360975 67694 360984
rect 67652 360262 67680 360975
rect 67640 360256 67692 360262
rect 67640 360198 67692 360204
rect 67638 359544 67694 359553
rect 67638 359479 67640 359488
rect 67692 359479 67694 359488
rect 67640 359450 67692 359456
rect 67730 358184 67786 358193
rect 67730 358119 67786 358128
rect 67640 358080 67692 358086
rect 67638 358048 67640 358057
rect 67692 358048 67694 358057
rect 67638 357983 67694 357992
rect 67744 357474 67772 358119
rect 67732 357468 67784 357474
rect 67732 357410 67784 357416
rect 67732 356176 67784 356182
rect 67732 356118 67784 356124
rect 67638 355600 67694 355609
rect 67638 355535 67694 355544
rect 67652 355366 67680 355535
rect 67744 355473 67772 356118
rect 67730 355464 67786 355473
rect 67730 355399 67786 355408
rect 67640 355360 67692 355366
rect 67640 355302 67692 355308
rect 67638 353832 67694 353841
rect 67638 353767 67694 353776
rect 67652 353326 67680 353767
rect 67640 353320 67692 353326
rect 67640 353262 67692 353268
rect 67638 352608 67694 352617
rect 67638 352543 67694 352552
rect 67916 352572 67968 352578
rect 67652 351966 67680 352543
rect 67916 352514 67968 352520
rect 67928 352481 67956 352514
rect 67914 352472 67970 352481
rect 67914 352407 67970 352416
rect 67640 351960 67692 351966
rect 67640 351902 67692 351908
rect 68296 351529 68324 449239
rect 68388 402974 68416 476983
rect 68926 469024 68982 469033
rect 68926 468959 68982 468968
rect 68388 402946 68784 402974
rect 68756 383722 68784 402946
rect 68836 386368 68888 386374
rect 68836 386310 68888 386316
rect 68848 385801 68876 386310
rect 68834 385792 68890 385801
rect 68834 385727 68890 385736
rect 68744 383716 68796 383722
rect 68744 383658 68796 383664
rect 68756 383489 68784 383658
rect 68742 383480 68798 383489
rect 68742 383415 68798 383424
rect 68376 376712 68428 376718
rect 68376 376654 68428 376660
rect 68388 365129 68416 376654
rect 68940 372881 68968 468959
rect 69124 454073 69152 553959
rect 69216 486577 69244 583714
rect 71792 581890 71820 583879
rect 71884 583030 71912 596146
rect 75196 586514 75224 702782
rect 75104 586486 75224 586514
rect 72240 585268 72292 585274
rect 72240 585210 72292 585216
rect 71872 583024 71924 583030
rect 71872 582966 71924 582972
rect 72252 581890 72280 585210
rect 74630 584352 74686 584361
rect 74630 584287 74686 584296
rect 73344 583772 73396 583778
rect 73344 583714 73396 583720
rect 73356 581890 73384 583714
rect 74644 581890 74672 584287
rect 75104 583982 75132 586486
rect 76576 585410 76604 702986
rect 79324 702568 79376 702574
rect 79324 702510 79376 702516
rect 78036 595468 78088 595474
rect 78036 595410 78088 595416
rect 76564 585404 76616 585410
rect 76564 585346 76616 585352
rect 75460 584112 75512 584118
rect 75460 584054 75512 584060
rect 75092 583976 75144 583982
rect 75092 583918 75144 583924
rect 75104 582162 75132 583918
rect 71792 581862 71944 581890
rect 72252 581862 72588 581890
rect 73278 581862 73384 581890
rect 74566 581862 74672 581890
rect 75012 582134 75132 582162
rect 75012 581754 75040 582134
rect 75472 581890 75500 584054
rect 76576 581890 76604 585346
rect 78048 585342 78076 595410
rect 78036 585336 78088 585342
rect 78036 585278 78088 585284
rect 77852 584112 77904 584118
rect 77852 584054 77904 584060
rect 77864 581890 77892 584054
rect 75472 581862 75808 581890
rect 76498 581862 76604 581890
rect 77786 581862 77892 581890
rect 78048 581890 78076 585278
rect 79336 584118 79364 702510
rect 89180 702434 89208 703520
rect 95148 703180 95200 703186
rect 95148 703122 95200 703128
rect 88352 702406 89208 702434
rect 85580 700392 85632 700398
rect 85580 700334 85632 700340
rect 83464 670744 83516 670750
rect 83464 670686 83516 670692
rect 83476 587858 83504 670686
rect 81716 587852 81768 587858
rect 81716 587794 81768 587800
rect 83464 587852 83516 587858
rect 83464 587794 83516 587800
rect 80612 586560 80664 586566
rect 80612 586502 80664 586508
rect 79324 584112 79376 584118
rect 79324 584054 79376 584060
rect 78680 582684 78732 582690
rect 78680 582626 78732 582632
rect 78692 581890 78720 582626
rect 79324 582548 79376 582554
rect 79324 582490 79376 582496
rect 79336 581890 79364 582490
rect 80624 581890 80652 586502
rect 81728 583914 81756 587794
rect 85120 586628 85172 586634
rect 85120 586570 85172 586576
rect 83186 586392 83242 586401
rect 83186 586327 83242 586336
rect 81440 583908 81492 583914
rect 81440 583850 81492 583856
rect 81716 583908 81768 583914
rect 81716 583850 81768 583856
rect 81452 581890 81480 583850
rect 81900 582616 81952 582622
rect 81900 582558 81952 582564
rect 81912 581890 81940 582558
rect 83200 581890 83228 586327
rect 84382 583944 84438 583953
rect 84382 583879 84438 583888
rect 84396 581890 84424 583879
rect 84474 583808 84530 583817
rect 84474 583743 84530 583752
rect 78048 581862 78384 581890
rect 78692 581862 79028 581890
rect 79336 581862 79672 581890
rect 80624 581862 80960 581890
rect 81452 581862 81604 581890
rect 81912 581862 82248 581890
rect 83200 581862 83536 581890
rect 84226 581862 84424 581890
rect 84488 581890 84516 583743
rect 85132 581890 85160 586570
rect 85592 585206 85620 700334
rect 87604 618316 87656 618322
rect 87604 618258 87656 618264
rect 87328 588600 87380 588606
rect 87328 588542 87380 588548
rect 87340 585206 87368 588542
rect 87616 587926 87644 618258
rect 87604 587920 87656 587926
rect 87604 587862 87656 587868
rect 88352 587178 88380 702406
rect 88340 587172 88392 587178
rect 88340 587114 88392 587120
rect 94136 586832 94188 586838
rect 94136 586774 94188 586780
rect 91560 586764 91612 586770
rect 91560 586706 91612 586712
rect 90272 586628 90324 586634
rect 90272 586570 90324 586576
rect 85580 585200 85632 585206
rect 85580 585142 85632 585148
rect 87328 585200 87380 585206
rect 87328 585142 87380 585148
rect 87512 585200 87564 585206
rect 87512 585142 87564 585148
rect 85592 581890 85620 585142
rect 87524 581890 87552 585142
rect 88984 583908 89036 583914
rect 88984 583850 89036 583856
rect 87696 583840 87748 583846
rect 87696 583782 87748 583788
rect 84488 581862 84824 581890
rect 85132 581862 85468 581890
rect 85592 581862 86112 581890
rect 87446 581862 87552 581890
rect 87708 581890 87736 583782
rect 88996 581890 89024 583850
rect 89628 582616 89680 582622
rect 89628 582558 89680 582564
rect 89640 581890 89668 582558
rect 90284 581890 90312 586570
rect 91006 584080 91062 584089
rect 91006 584015 91062 584024
rect 91020 581890 91048 584015
rect 91572 581890 91600 586706
rect 92296 585268 92348 585274
rect 92296 585210 92348 585216
rect 92308 581890 92336 585210
rect 92846 582448 92902 582457
rect 92846 582383 92902 582392
rect 92860 581890 92888 582383
rect 94148 581890 94176 586774
rect 94872 586696 94924 586702
rect 94872 586638 94924 586644
rect 94884 581890 94912 586638
rect 95160 585342 95188 703122
rect 104808 702976 104860 702982
rect 104808 702918 104860 702924
rect 97264 700392 97316 700398
rect 97264 700334 97316 700340
rect 97276 589966 97304 700334
rect 97264 589960 97316 589966
rect 97264 589902 97316 589908
rect 95240 587920 95292 587926
rect 95240 587862 95292 587868
rect 95252 585410 95280 587862
rect 98736 586560 98788 586566
rect 98736 586502 98788 586508
rect 95240 585404 95292 585410
rect 95240 585346 95292 585352
rect 95884 585404 95936 585410
rect 95884 585346 95936 585352
rect 95148 585336 95200 585342
rect 95148 585278 95200 585284
rect 95160 582162 95188 585278
rect 87708 581862 88044 581890
rect 88734 581862 89024 581890
rect 89378 581862 89668 581890
rect 90022 581862 90312 581890
rect 90666 581862 91048 581890
rect 91310 581862 91600 581890
rect 91954 581862 92336 581890
rect 92598 581862 92888 581890
rect 93886 581862 94176 581890
rect 94530 581862 94912 581890
rect 94976 582134 95188 582162
rect 82728 581800 82780 581806
rect 70964 581738 71300 581754
rect 70400 581732 70452 581738
rect 70400 581674 70452 581680
rect 70952 581732 71300 581738
rect 71004 581726 71300 581732
rect 75012 581726 75164 581754
rect 76760 581738 77096 581754
rect 94976 581754 95004 582134
rect 95896 581890 95924 585346
rect 96528 583840 96580 583846
rect 96528 583782 96580 583788
rect 97906 583808 97962 583817
rect 96540 581890 96568 583782
rect 97448 583772 97500 583778
rect 97906 583743 97962 583752
rect 97448 583714 97500 583720
rect 97460 581890 97488 583714
rect 97920 581890 97948 583743
rect 98748 581890 98776 586502
rect 104820 584458 104848 702918
rect 105464 702434 105492 703520
rect 116584 703112 116636 703118
rect 116584 703054 116636 703060
rect 113088 702908 113140 702914
rect 113088 702850 113140 702856
rect 110328 702772 110380 702778
rect 110328 702714 110380 702720
rect 105464 702406 105584 702434
rect 105556 596174 105584 702406
rect 106280 698964 106332 698970
rect 106280 698906 106332 698912
rect 105556 596146 105676 596174
rect 103152 584452 103204 584458
rect 103152 584394 103204 584400
rect 104808 584452 104860 584458
rect 104808 584394 104860 584400
rect 101312 584044 101364 584050
rect 101312 583986 101364 583992
rect 100760 583908 100812 583914
rect 100760 583850 100812 583856
rect 100772 583030 100800 583850
rect 100760 583024 100812 583030
rect 100760 582966 100812 582972
rect 99288 582548 99340 582554
rect 99288 582490 99340 582496
rect 99300 581890 99328 582490
rect 101324 581890 101352 583986
rect 101864 583976 101916 583982
rect 101864 583918 101916 583924
rect 101876 581890 101904 583918
rect 103164 581890 103192 584394
rect 105544 583908 105596 583914
rect 105544 583850 105596 583856
rect 103888 582480 103940 582486
rect 103888 582422 103940 582428
rect 103900 581890 103928 582422
rect 105556 581890 105584 583850
rect 95818 581862 95924 581890
rect 96462 581862 96568 581890
rect 97106 581862 97488 581890
rect 97750 581862 97948 581890
rect 98394 581862 98776 581890
rect 99038 581862 99328 581890
rect 100970 581862 101352 581890
rect 101614 581862 101904 581890
rect 102902 581862 103192 581890
rect 103546 581862 103928 581890
rect 105478 581862 105584 581890
rect 104992 581800 105044 581806
rect 102598 581768 102654 581777
rect 82780 581748 82892 581754
rect 82728 581742 82892 581748
rect 76748 581732 77096 581738
rect 70952 581674 71004 581680
rect 76800 581726 77096 581732
rect 82740 581726 82892 581742
rect 94976 581726 95128 581754
rect 100326 581738 100616 581754
rect 100326 581732 100628 581738
rect 100326 581726 100576 581732
rect 76748 581674 76800 581680
rect 102258 581726 102598 581754
rect 104190 581738 104480 581754
rect 104834 581748 104992 581754
rect 104834 581742 105044 581748
rect 104190 581732 104492 581738
rect 104190 581726 104440 581732
rect 102598 581703 102654 581712
rect 100576 581674 100628 581680
rect 104834 581726 105032 581742
rect 104440 581674 104492 581680
rect 69308 581318 70058 581346
rect 69202 486568 69258 486577
rect 69202 486503 69258 486512
rect 69308 482633 69336 581318
rect 70412 581262 70440 581674
rect 70504 581318 70702 581346
rect 70400 581256 70452 581262
rect 70400 581198 70452 581204
rect 70504 581058 70532 581318
rect 70492 581052 70544 581058
rect 70492 580994 70544 581000
rect 105648 572354 105676 596146
rect 105636 572348 105688 572354
rect 105636 572290 105688 572296
rect 106292 560425 106320 698906
rect 107106 583944 107162 583953
rect 107106 583879 107162 583888
rect 106738 583808 106794 583817
rect 106738 583743 106794 583752
rect 106752 578950 106780 583743
rect 106740 578944 106792 578950
rect 107120 578921 107148 583879
rect 107660 582752 107712 582758
rect 107660 582694 107712 582700
rect 106740 578886 106792 578892
rect 107106 578912 107162 578921
rect 107106 578847 107162 578856
rect 106462 578096 106518 578105
rect 106462 578031 106518 578040
rect 106370 574696 106426 574705
rect 106370 574631 106426 574640
rect 106278 560416 106334 560425
rect 106278 560351 106334 560360
rect 106186 552120 106242 552129
rect 106186 552055 106242 552064
rect 105818 543824 105874 543833
rect 105818 543759 105874 543768
rect 69768 540110 70058 540138
rect 70412 540110 70702 540138
rect 69768 537674 69796 540110
rect 69756 537668 69808 537674
rect 69756 537610 69808 537616
rect 70412 532273 70440 540110
rect 71332 536110 71360 540138
rect 71320 536104 71372 536110
rect 71320 536046 71372 536052
rect 71044 535016 71096 535022
rect 71044 534958 71096 534964
rect 70398 532264 70454 532273
rect 70398 532199 70454 532208
rect 71056 499574 71084 534958
rect 71976 529310 72004 540138
rect 71964 529304 72016 529310
rect 71964 529246 72016 529252
rect 70872 499546 71084 499574
rect 70308 493332 70360 493338
rect 70308 493274 70360 493280
rect 70032 492108 70084 492114
rect 70032 492050 70084 492056
rect 69756 490612 69808 490618
rect 69756 490554 69808 490560
rect 69768 489977 69796 490554
rect 69754 489968 69810 489977
rect 70044 489940 70072 492050
rect 70320 491314 70348 493274
rect 70320 491286 70440 491314
rect 70412 489954 70440 491286
rect 70412 489926 70656 489954
rect 69754 489903 69810 489912
rect 70872 489870 70900 499546
rect 72620 497554 72648 540138
rect 73264 534886 73292 540138
rect 73908 538150 73936 540138
rect 73896 538144 73948 538150
rect 73896 538086 73948 538092
rect 73252 534880 73304 534886
rect 73252 534822 73304 534828
rect 74552 532001 74580 540138
rect 74724 537532 74776 537538
rect 74724 537474 74776 537480
rect 74538 531992 74594 532001
rect 74538 531927 74594 531936
rect 72608 497548 72660 497554
rect 72608 497490 72660 497496
rect 73252 494896 73304 494902
rect 73252 494838 73304 494844
rect 72240 492040 72292 492046
rect 72240 491982 72292 491988
rect 71136 491700 71188 491706
rect 71136 491642 71188 491648
rect 71148 489954 71176 491642
rect 71780 491496 71832 491502
rect 71780 491438 71832 491444
rect 71792 489954 71820 491438
rect 72252 489954 72280 491982
rect 71148 489926 71300 489954
rect 71792 489926 71944 489954
rect 72252 489926 72588 489954
rect 73264 489940 73292 494838
rect 74736 494834 74764 537474
rect 75196 534954 75224 540138
rect 76467 540110 76512 540138
rect 75184 534948 75236 534954
rect 75184 534890 75236 534896
rect 76484 532137 76512 540110
rect 76562 537568 76618 537577
rect 76562 537503 76618 537512
rect 76470 532128 76526 532137
rect 76470 532063 76526 532072
rect 76576 499574 76604 537503
rect 77128 529242 77156 540138
rect 77116 529236 77168 529242
rect 77116 529178 77168 529184
rect 76576 499546 76696 499574
rect 75828 496120 75880 496126
rect 75828 496062 75880 496068
rect 74724 494828 74776 494834
rect 74724 494770 74776 494776
rect 74540 494080 74592 494086
rect 74540 494022 74592 494028
rect 74552 489940 74580 494022
rect 75000 492924 75052 492930
rect 75000 492866 75052 492872
rect 75012 489954 75040 492866
rect 75012 489926 75164 489954
rect 75840 489940 75868 496062
rect 76104 494828 76156 494834
rect 76104 494770 76156 494776
rect 76116 489954 76144 494770
rect 76668 494086 76696 499546
rect 77772 497622 77800 540138
rect 78416 534750 78444 540138
rect 78404 534744 78456 534750
rect 78404 534686 78456 534692
rect 77760 497616 77812 497622
rect 77760 497558 77812 497564
rect 77758 495544 77814 495553
rect 77758 495479 77814 495488
rect 76656 494080 76708 494086
rect 76656 494022 76708 494028
rect 76668 489954 76696 494022
rect 76116 489926 76452 489954
rect 76668 489926 77096 489954
rect 77772 489940 77800 495479
rect 78036 491972 78088 491978
rect 78036 491914 78088 491920
rect 78048 489954 78076 491914
rect 79060 490686 79088 540138
rect 79704 535022 79732 540138
rect 80348 537470 80376 540138
rect 80336 537464 80388 537470
rect 80336 537406 80388 537412
rect 79692 535016 79744 535022
rect 79692 534958 79744 534964
rect 80992 499574 81020 540138
rect 81440 537464 81492 537470
rect 81636 537441 81664 540138
rect 82907 540110 82952 540138
rect 82924 537606 82952 540110
rect 83004 538892 83056 538898
rect 83004 538834 83056 538840
rect 82912 537600 82964 537606
rect 82912 537542 82964 537548
rect 81440 537406 81492 537412
rect 81622 537432 81678 537441
rect 80900 499546 81020 499574
rect 79324 492856 79376 492862
rect 79324 492798 79376 492804
rect 79048 490680 79100 490686
rect 79048 490622 79100 490628
rect 79336 489954 79364 492798
rect 80060 491360 80112 491366
rect 80060 491302 80112 491308
rect 80072 489954 80100 491302
rect 80900 490521 80928 499546
rect 81452 496262 81480 537406
rect 81622 537367 81678 537376
rect 81440 496256 81492 496262
rect 81440 496198 81492 496204
rect 81440 496120 81492 496126
rect 81440 496062 81492 496068
rect 81452 495514 81480 496062
rect 81440 495508 81492 495514
rect 81440 495450 81492 495456
rect 82912 494828 82964 494834
rect 82912 494770 82964 494776
rect 82820 494760 82872 494766
rect 82820 494702 82872 494708
rect 80980 494148 81032 494154
rect 80980 494090 81032 494096
rect 80886 490512 80942 490521
rect 80886 490447 80942 490456
rect 78048 489926 78384 489954
rect 79336 489926 79672 489954
rect 80072 489926 80316 489954
rect 80992 489940 81020 494090
rect 82832 494018 82860 494702
rect 82820 494012 82872 494018
rect 82820 493954 82872 493960
rect 81624 491972 81676 491978
rect 81624 491914 81676 491920
rect 81636 489940 81664 491914
rect 82268 491564 82320 491570
rect 82268 491506 82320 491512
rect 82280 489940 82308 491506
rect 82924 489940 82952 494770
rect 83016 491978 83044 538834
rect 83464 536852 83516 536858
rect 83464 536794 83516 536800
rect 83004 491972 83056 491978
rect 83004 491914 83056 491920
rect 83476 490754 83504 536794
rect 83568 534818 83596 540138
rect 83556 534812 83608 534818
rect 83556 534754 83608 534760
rect 84212 500274 84240 540138
rect 84856 536858 84884 540138
rect 85500 537674 85528 540138
rect 85488 537668 85540 537674
rect 85488 537610 85540 537616
rect 84844 536852 84896 536858
rect 84844 536794 84896 536800
rect 84200 500268 84252 500274
rect 84200 500210 84252 500216
rect 85488 494420 85540 494426
rect 85488 494362 85540 494368
rect 83556 494012 83608 494018
rect 83556 493954 83608 493960
rect 83464 490748 83516 490754
rect 83464 490690 83516 490696
rect 83568 489940 83596 493954
rect 84842 490104 84898 490113
rect 84842 490039 84898 490048
rect 84856 489940 84884 490039
rect 85500 489940 85528 494362
rect 86144 490822 86172 540138
rect 86788 497622 86816 540138
rect 87432 532098 87460 540138
rect 88076 538898 88104 540138
rect 89347 540110 89392 540138
rect 88064 538892 88116 538898
rect 88064 538834 88116 538840
rect 89364 537441 89392 540110
rect 89350 537432 89406 537441
rect 89350 537367 89406 537376
rect 90008 534886 90036 540138
rect 89996 534880 90048 534886
rect 89996 534822 90048 534828
rect 87420 532092 87472 532098
rect 87420 532034 87472 532040
rect 86776 497616 86828 497622
rect 86776 497558 86828 497564
rect 89628 496188 89680 496194
rect 89628 496130 89680 496136
rect 88064 496120 88116 496126
rect 88064 496062 88116 496068
rect 87420 492652 87472 492658
rect 87420 492594 87472 492600
rect 86408 491632 86460 491638
rect 86408 491574 86460 491580
rect 86132 490816 86184 490822
rect 86132 490758 86184 490764
rect 86420 489954 86448 491574
rect 86158 489926 86448 489954
rect 86802 489938 87000 489954
rect 87432 489940 87460 492594
rect 88076 489940 88104 496062
rect 89640 494426 89668 496130
rect 90652 494737 90680 540138
rect 91296 539510 91324 540138
rect 91284 539504 91336 539510
rect 91284 539446 91336 539452
rect 91940 499574 91968 540138
rect 92584 532030 92612 540138
rect 92572 532024 92624 532030
rect 92572 531966 92624 531972
rect 93228 499574 93256 540138
rect 93872 534750 93900 540138
rect 94516 538150 94544 540138
rect 95787 540110 95832 540138
rect 95148 538960 95200 538966
rect 95148 538902 95200 538908
rect 94504 538144 94556 538150
rect 94504 538086 94556 538092
rect 95056 534812 95108 534818
rect 95056 534754 95108 534760
rect 93860 534744 93912 534750
rect 93860 534686 93912 534692
rect 93768 532160 93820 532166
rect 93768 532102 93820 532108
rect 91940 499546 92060 499574
rect 93228 499546 93348 499574
rect 91284 497548 91336 497554
rect 91284 497490 91336 497496
rect 90638 494728 90694 494737
rect 90638 494663 90694 494672
rect 89628 494420 89680 494426
rect 89628 494362 89680 494368
rect 90272 493468 90324 493474
rect 90272 493410 90324 493416
rect 90284 492794 90312 493410
rect 90272 492788 90324 492794
rect 90272 492730 90324 492736
rect 89996 491428 90048 491434
rect 89996 491370 90048 491376
rect 88984 490680 89036 490686
rect 88984 490622 89036 490628
rect 88996 489954 89024 490622
rect 86802 489932 87012 489938
rect 86802 489926 86960 489932
rect 88734 489926 89024 489954
rect 90008 489940 90036 491370
rect 90284 489954 90312 492730
rect 90284 489926 90620 489954
rect 91296 489940 91324 497490
rect 91928 493400 91980 493406
rect 91928 493342 91980 493348
rect 91940 489940 91968 493342
rect 92032 490657 92060 499546
rect 92572 497480 92624 497486
rect 92572 497422 92624 497428
rect 92480 492788 92532 492794
rect 92480 492730 92532 492736
rect 92492 492658 92520 492730
rect 92480 492652 92532 492658
rect 92480 492594 92532 492600
rect 92018 490648 92074 490657
rect 92018 490583 92074 490592
rect 92584 489940 92612 497422
rect 93216 493332 93268 493338
rect 93216 493274 93268 493280
rect 92846 491600 92902 491609
rect 92846 491535 92902 491544
rect 92860 491434 92888 491535
rect 92848 491428 92900 491434
rect 92848 491370 92900 491376
rect 93228 489940 93256 493274
rect 93320 492182 93348 499546
rect 93780 492794 93808 532102
rect 93768 492788 93820 492794
rect 93768 492730 93820 492736
rect 93308 492176 93360 492182
rect 93308 492118 93360 492124
rect 95068 490618 95096 534754
rect 95160 493406 95188 538902
rect 95804 537742 95832 540110
rect 95792 537736 95844 537742
rect 95792 537678 95844 537684
rect 96448 497690 96476 540138
rect 97092 532234 97120 540138
rect 97080 532228 97132 532234
rect 97080 532170 97132 532176
rect 96436 497684 96488 497690
rect 96436 497626 96488 497632
rect 97736 494766 97764 540138
rect 98380 538218 98408 540138
rect 99024 539578 99052 540138
rect 99012 539572 99064 539578
rect 99012 539514 99064 539520
rect 99024 539034 99052 539514
rect 99196 539096 99248 539102
rect 99196 539038 99248 539044
rect 99012 539028 99064 539034
rect 99012 538970 99064 538976
rect 98368 538212 98420 538218
rect 99208 538214 99236 539038
rect 99668 538214 99696 540138
rect 99208 538186 99328 538214
rect 99668 538186 99788 538214
rect 98368 538154 98420 538160
rect 98380 537606 98408 538154
rect 98644 537668 98696 537674
rect 98644 537610 98696 537616
rect 98368 537600 98420 537606
rect 98368 537542 98420 537548
rect 97906 536072 97962 536081
rect 97906 536007 97962 536016
rect 97816 534948 97868 534954
rect 97816 534890 97868 534896
rect 97724 494760 97776 494766
rect 97724 494702 97776 494708
rect 95792 494692 95844 494698
rect 95792 494634 95844 494640
rect 95148 493400 95200 493406
rect 95148 493342 95200 493348
rect 94136 490612 94188 490618
rect 94136 490554 94188 490560
rect 95056 490612 95108 490618
rect 95056 490554 95108 490560
rect 94148 489954 94176 490554
rect 95146 490512 95202 490521
rect 95146 490447 95202 490456
rect 93886 489926 94176 489954
rect 95160 489940 95188 490447
rect 95804 489940 95832 494634
rect 97080 492040 97132 492046
rect 97080 491982 97132 491988
rect 96436 491836 96488 491842
rect 96436 491778 96488 491784
rect 96448 489940 96476 491778
rect 97092 489940 97120 491982
rect 97828 491473 97856 534890
rect 97920 492114 97948 536007
rect 98656 494902 98684 537610
rect 98644 494896 98696 494902
rect 98644 494838 98696 494844
rect 97908 492108 97960 492114
rect 97908 492050 97960 492056
rect 97920 491842 97948 492050
rect 97908 491836 97960 491842
rect 97908 491778 97960 491784
rect 97814 491464 97870 491473
rect 97814 491399 97870 491408
rect 97828 489954 97856 491399
rect 99300 491337 99328 538186
rect 99378 536888 99434 536897
rect 99378 536823 99434 536832
rect 99286 491328 99342 491337
rect 99286 491263 99342 491272
rect 99300 489954 99328 491263
rect 97750 489926 97856 489954
rect 99038 489926 99328 489954
rect 86960 489874 87012 489880
rect 69848 489864 69900 489870
rect 69848 489806 69900 489812
rect 70860 489864 70912 489870
rect 98736 489864 98788 489870
rect 70860 489806 70912 489812
rect 98394 489812 98736 489818
rect 98394 489806 98788 489812
rect 99288 489864 99340 489870
rect 99288 489806 99340 489812
rect 69860 489161 69888 489806
rect 98394 489790 98776 489806
rect 99300 489297 99328 489806
rect 99286 489288 99342 489297
rect 99286 489223 99342 489232
rect 69846 489152 69902 489161
rect 69846 489087 69902 489096
rect 69294 482624 69350 482633
rect 69294 482559 69350 482568
rect 69386 482488 69442 482497
rect 69386 482423 69442 482432
rect 69202 458008 69258 458017
rect 69202 457943 69258 457952
rect 69110 454064 69166 454073
rect 69110 453999 69166 454008
rect 68926 372872 68982 372881
rect 68926 372807 68982 372816
rect 68374 365120 68430 365129
rect 68374 365055 68430 365064
rect 69124 356969 69152 453999
rect 69216 361622 69244 457943
rect 69400 438394 69428 482423
rect 99392 446593 99420 536823
rect 99656 491428 99708 491434
rect 99656 491370 99708 491376
rect 99668 489940 99696 491370
rect 99470 476368 99526 476377
rect 99470 476303 99526 476312
rect 99378 446584 99434 446593
rect 99378 446519 99434 446528
rect 99286 442504 99342 442513
rect 99286 442439 99342 442448
rect 69846 441280 69902 441289
rect 69846 441215 69902 441224
rect 69860 440706 69888 441215
rect 99300 441153 99328 442439
rect 99286 441144 99342 441153
rect 99286 441079 99342 441088
rect 79322 440736 79378 440745
rect 72344 440706 73016 440722
rect 69848 440700 69900 440706
rect 69848 440642 69900 440648
rect 70400 440700 70452 440706
rect 70400 440642 70452 440648
rect 72332 440700 73016 440706
rect 72384 440694 73016 440700
rect 72332 440642 72384 440648
rect 70412 440042 70440 440642
rect 71136 440292 71188 440298
rect 71136 440234 71188 440240
rect 70412 440028 70702 440042
rect 70044 438666 70072 440028
rect 70412 440014 70716 440028
rect 70032 438660 70084 438666
rect 70032 438602 70084 438608
rect 69388 438388 69440 438394
rect 69388 438330 69440 438336
rect 70044 437918 70072 438602
rect 69296 437912 69348 437918
rect 69296 437854 69348 437860
rect 70032 437912 70084 437918
rect 70032 437854 70084 437860
rect 69308 364334 69336 437854
rect 70688 437753 70716 440014
rect 71042 438968 71098 438977
rect 71042 438903 71098 438912
rect 70674 437744 70730 437753
rect 70674 437679 70730 437688
rect 70400 395004 70452 395010
rect 70400 394946 70452 394952
rect 69756 388136 69808 388142
rect 69756 388078 69808 388084
rect 69768 385914 69796 388078
rect 70412 385914 70440 394946
rect 71056 387841 71084 438903
rect 71148 395010 71176 440234
rect 71332 434722 71360 440028
rect 71792 440014 71990 440042
rect 71320 434716 71372 434722
rect 71320 434658 71372 434664
rect 71792 431905 71820 440014
rect 72988 438938 73016 440694
rect 79322 440671 79378 440680
rect 81438 440736 81494 440745
rect 81494 440694 81650 440722
rect 87446 440706 87736 440722
rect 87446 440700 87748 440706
rect 87446 440694 87696 440700
rect 81438 440671 81494 440680
rect 73278 440014 73384 440042
rect 72976 438932 73028 438938
rect 72976 438874 73028 438880
rect 71872 438388 71924 438394
rect 71872 438330 71924 438336
rect 71778 431896 71834 431905
rect 71778 431831 71834 431840
rect 71136 395004 71188 395010
rect 71136 394946 71188 394952
rect 71148 394738 71176 394946
rect 71136 394732 71188 394738
rect 71136 394674 71188 394680
rect 71780 389224 71832 389230
rect 71780 389166 71832 389172
rect 71042 387832 71098 387841
rect 71042 387767 71098 387776
rect 71792 385914 71820 389166
rect 71884 388890 71912 438330
rect 73356 437374 73384 440014
rect 73908 439006 73936 440028
rect 73896 439000 73948 439006
rect 73896 438942 73948 438948
rect 73436 438932 73488 438938
rect 73436 438874 73488 438880
rect 73344 437368 73396 437374
rect 73344 437310 73396 437316
rect 71872 388884 71924 388890
rect 71872 388826 71924 388832
rect 72332 388884 72384 388890
rect 72332 388826 72384 388832
rect 72344 387938 72372 388826
rect 72332 387932 72384 387938
rect 72332 387874 72384 387880
rect 72344 385914 72372 387874
rect 69768 385886 70058 385914
rect 70412 385886 70702 385914
rect 71792 385886 71990 385914
rect 72344 385886 72634 385914
rect 70308 385824 70360 385830
rect 70308 385766 70360 385772
rect 73356 385778 73384 437310
rect 73448 385898 73476 438874
rect 74552 434625 74580 440028
rect 75840 439074 75868 440028
rect 76012 439544 76064 439550
rect 76012 439486 76064 439492
rect 74632 439068 74684 439074
rect 74632 439010 74684 439016
rect 75828 439068 75880 439074
rect 75828 439010 75880 439016
rect 74538 434616 74594 434625
rect 74538 434551 74594 434560
rect 74644 431954 74672 439010
rect 75184 438252 75236 438258
rect 75184 438194 75236 438200
rect 74552 431926 74672 431954
rect 73526 387832 73582 387841
rect 73526 387767 73582 387776
rect 73436 385892 73488 385898
rect 73436 385834 73488 385840
rect 70320 378826 70348 385766
rect 73356 385750 73476 385778
rect 73448 385694 73476 385750
rect 73436 385688 73488 385694
rect 73436 385630 73488 385636
rect 73540 385506 73568 387767
rect 74552 387190 74580 431926
rect 74632 400240 74684 400246
rect 74632 400182 74684 400188
rect 74540 387184 74592 387190
rect 74540 387126 74592 387132
rect 74644 385914 74672 400182
rect 75196 388142 75224 438194
rect 75276 436756 75328 436762
rect 75276 436698 75328 436704
rect 75288 400246 75316 436698
rect 75276 400240 75328 400246
rect 75276 400182 75328 400188
rect 75920 399492 75972 399498
rect 75920 399434 75972 399440
rect 75932 393378 75960 399434
rect 75920 393372 75972 393378
rect 75920 393314 75972 393320
rect 75828 388476 75880 388482
rect 75828 388418 75880 388424
rect 75184 388136 75236 388142
rect 75184 388078 75236 388084
rect 75552 388136 75604 388142
rect 75552 388078 75604 388084
rect 75564 385914 75592 388078
rect 75840 387938 75868 388418
rect 75828 387932 75880 387938
rect 75828 387874 75880 387880
rect 75840 386186 75868 387874
rect 74566 385886 74672 385914
rect 75210 385886 75592 385914
rect 75656 386158 75868 386186
rect 75656 385778 75684 386158
rect 75932 386050 75960 393314
rect 76024 387705 76052 439486
rect 76484 434042 76512 440028
rect 77128 438734 77156 440028
rect 77772 439550 77800 440028
rect 77760 439544 77812 439550
rect 77760 439486 77812 439492
rect 77942 439512 77998 439521
rect 77942 439447 77998 439456
rect 77116 438728 77168 438734
rect 77116 438670 77168 438676
rect 76472 434036 76524 434042
rect 76472 433978 76524 433984
rect 77956 394670 77984 439447
rect 78416 438802 78444 440028
rect 78404 438796 78456 438802
rect 78404 438738 78456 438744
rect 78416 437578 78444 438738
rect 78678 437608 78734 437617
rect 78404 437572 78456 437578
rect 78678 437543 78734 437552
rect 78404 437514 78456 437520
rect 77944 394664 77996 394670
rect 77944 394606 77996 394612
rect 77956 393314 77984 394606
rect 77864 393286 77984 393314
rect 76010 387696 76066 387705
rect 76010 387631 76066 387640
rect 75932 386022 76696 386050
rect 76668 385914 76696 386022
rect 77864 385914 77892 393286
rect 78692 392630 78720 437543
rect 79060 437510 79088 440028
rect 79048 437504 79100 437510
rect 79048 437446 79100 437452
rect 79336 394058 79364 440671
rect 87696 440642 87748 440648
rect 88432 440700 88484 440706
rect 88432 440642 88484 440648
rect 79704 438841 79732 440028
rect 80624 440014 81006 440042
rect 81912 440014 82294 440042
rect 80624 439142 80652 440014
rect 80612 439136 80664 439142
rect 80612 439078 80664 439084
rect 79690 438832 79746 438841
rect 79690 438767 79746 438776
rect 79704 437617 79732 438767
rect 79690 437608 79746 437617
rect 79690 437543 79746 437552
rect 80704 437572 80756 437578
rect 80704 437514 80756 437520
rect 80060 437504 80112 437510
rect 80060 437446 80112 437452
rect 80072 436082 80100 437446
rect 80060 436076 80112 436082
rect 80060 436018 80112 436024
rect 80072 396914 80100 436018
rect 80716 431254 80744 437514
rect 81912 437481 81940 440014
rect 81898 437472 81954 437481
rect 81898 437407 81954 437416
rect 81912 431954 81940 437407
rect 82924 437306 82952 440028
rect 83568 438190 83596 440028
rect 84212 438977 84240 440028
rect 84198 438968 84254 438977
rect 84198 438903 84254 438912
rect 83556 438184 83608 438190
rect 83556 438126 83608 438132
rect 84856 437510 84884 440028
rect 86158 440014 86264 440042
rect 83648 437504 83700 437510
rect 83648 437446 83700 437452
rect 84844 437504 84896 437510
rect 84844 437446 84896 437452
rect 85028 437504 85080 437510
rect 85028 437446 85080 437452
rect 82912 437300 82964 437306
rect 82912 437242 82964 437248
rect 82924 431954 82952 437242
rect 83660 436014 83688 437446
rect 83096 436008 83148 436014
rect 83096 435950 83148 435956
rect 83648 436008 83700 436014
rect 83648 435950 83700 435956
rect 81544 431926 81940 431954
rect 82832 431926 82952 431954
rect 80704 431248 80756 431254
rect 80704 431190 80756 431196
rect 80060 396908 80112 396914
rect 80060 396850 80112 396856
rect 80716 396846 80744 431190
rect 80704 396840 80756 396846
rect 80704 396782 80756 396788
rect 79324 394052 79376 394058
rect 79324 393994 79376 394000
rect 81440 393984 81492 393990
rect 81440 393926 81492 393932
rect 81452 393446 81480 393926
rect 81440 393440 81492 393446
rect 81440 393382 81492 393388
rect 78680 392624 78732 392630
rect 78680 392566 78732 392572
rect 79324 388068 79376 388074
rect 79324 388010 79376 388016
rect 78036 388000 78088 388006
rect 78036 387942 78088 387948
rect 76668 385886 77142 385914
rect 77786 385886 77892 385914
rect 78048 385914 78076 387942
rect 79336 385914 79364 388010
rect 80060 387864 80112 387870
rect 80060 387806 80112 387812
rect 80072 385914 80100 387806
rect 80612 386504 80664 386510
rect 80612 386446 80664 386452
rect 80624 385914 80652 386446
rect 81452 386050 81480 393382
rect 81544 391241 81572 431926
rect 82832 391542 82860 431926
rect 82912 394120 82964 394126
rect 82912 394062 82964 394068
rect 82820 391536 82872 391542
rect 82820 391478 82872 391484
rect 82820 391400 82872 391406
rect 82820 391342 82872 391348
rect 81530 391232 81586 391241
rect 81530 391167 81586 391176
rect 82832 390590 82860 391342
rect 82924 390658 82952 394062
rect 82912 390652 82964 390658
rect 82912 390594 82964 390600
rect 82820 390584 82872 390590
rect 82820 390526 82872 390532
rect 83004 390584 83056 390590
rect 83004 390526 83056 390532
rect 82452 388136 82504 388142
rect 82452 388078 82504 388084
rect 81452 386022 81848 386050
rect 81820 385914 81848 386022
rect 78048 385886 78430 385914
rect 79336 385886 79718 385914
rect 80072 385886 80362 385914
rect 80624 385886 81006 385914
rect 81820 385886 82294 385914
rect 75656 385750 75854 385778
rect 73278 385478 73568 385506
rect 77864 385370 77892 385886
rect 82464 385694 82492 388078
rect 83016 385914 83044 390526
rect 82938 385886 83044 385914
rect 83108 385830 83136 435950
rect 85040 435946 85068 437446
rect 86236 437374 86264 440014
rect 86788 437510 86816 440028
rect 88090 440014 88288 440042
rect 86776 437504 86828 437510
rect 86776 437446 86828 437452
rect 86224 437368 86276 437374
rect 86224 437310 86276 437316
rect 84200 435940 84252 435946
rect 84200 435882 84252 435888
rect 85028 435940 85080 435946
rect 85028 435882 85080 435888
rect 84212 399673 84240 435882
rect 86236 402974 86264 437310
rect 88260 436082 88288 440014
rect 88248 436076 88300 436082
rect 88248 436018 88300 436024
rect 86236 402946 86356 402974
rect 84198 399664 84254 399673
rect 84198 399599 84254 399608
rect 85118 399528 85174 399537
rect 85118 399463 85174 399472
rect 85132 396098 85160 399463
rect 84200 396092 84252 396098
rect 84200 396034 84252 396040
rect 85120 396092 85172 396098
rect 85120 396034 85172 396040
rect 83648 390652 83700 390658
rect 83648 390594 83700 390600
rect 83660 385914 83688 390594
rect 84212 386050 84240 396034
rect 84212 386022 84424 386050
rect 83582 385886 83688 385914
rect 84396 385914 84424 386022
rect 85132 385914 85160 396034
rect 85948 391264 86000 391270
rect 85948 391206 86000 391212
rect 85960 386481 85988 391206
rect 85946 386472 86002 386481
rect 85946 386407 86002 386416
rect 84396 385886 84870 385914
rect 85132 385886 85514 385914
rect 83096 385824 83148 385830
rect 83096 385766 83148 385772
rect 85960 385778 85988 386407
rect 85960 385750 86158 385778
rect 82452 385688 82504 385694
rect 82452 385630 82504 385636
rect 86328 385626 86356 402946
rect 88260 402286 88288 436018
rect 88248 402280 88300 402286
rect 88248 402222 88300 402228
rect 88340 395344 88392 395350
rect 88340 395286 88392 395292
rect 88352 394806 88380 395286
rect 88340 394800 88392 394806
rect 88340 394742 88392 394748
rect 87696 393984 87748 393990
rect 87696 393926 87748 393932
rect 87052 386436 87104 386442
rect 87052 386378 87104 386384
rect 87064 385914 87092 386378
rect 87708 385914 87736 393926
rect 88352 385914 88380 394742
rect 88444 392698 88472 440642
rect 97448 440224 97500 440230
rect 97106 440172 97448 440178
rect 97106 440166 97500 440172
rect 98644 440224 98696 440230
rect 98644 440166 98696 440172
rect 97106 440150 97488 440166
rect 88720 439006 88748 440028
rect 89378 440014 89668 440042
rect 90022 440014 90404 440042
rect 88708 439000 88760 439006
rect 88708 438942 88760 438948
rect 89640 435985 89668 440014
rect 90376 438705 90404 440014
rect 91296 438841 91324 440028
rect 91756 440014 91954 440042
rect 91282 438832 91338 438841
rect 91282 438767 91338 438776
rect 90362 438696 90418 438705
rect 90362 438631 90418 438640
rect 89626 435976 89682 435985
rect 89626 435911 89682 435920
rect 89640 398206 89668 435911
rect 89628 398200 89680 398206
rect 89628 398142 89680 398148
rect 88432 392692 88484 392698
rect 88432 392634 88484 392640
rect 90272 387864 90324 387870
rect 90272 387806 90324 387812
rect 90284 385914 90312 387806
rect 90376 387122 90404 438631
rect 91100 437640 91152 437646
rect 91020 437588 91100 437594
rect 91020 437582 91152 437588
rect 91020 437566 91140 437582
rect 91020 393314 91048 437566
rect 91756 437442 91784 440014
rect 92584 439113 92612 440028
rect 92570 439104 92626 439113
rect 92570 439039 92626 439048
rect 92584 437646 92612 439039
rect 93228 438666 93256 440028
rect 93872 439056 93900 440028
rect 93780 439028 93900 439056
rect 93780 438818 93808 439028
rect 93860 438932 93912 438938
rect 93860 438874 93912 438880
rect 93688 438790 93808 438818
rect 93216 438660 93268 438666
rect 93216 438602 93268 438608
rect 93688 438530 93716 438790
rect 93768 438660 93820 438666
rect 93768 438602 93820 438608
rect 93676 438524 93728 438530
rect 93676 438466 93728 438472
rect 92572 437640 92624 437646
rect 92572 437582 92624 437588
rect 91744 437436 91796 437442
rect 91744 437378 91796 437384
rect 91756 396846 91784 437378
rect 93688 404977 93716 438466
rect 93674 404968 93730 404977
rect 93674 404903 93730 404912
rect 91836 404388 91888 404394
rect 91836 404330 91888 404336
rect 91744 396840 91796 396846
rect 91744 396782 91796 396788
rect 91848 394670 91876 404330
rect 93780 399537 93808 438602
rect 93766 399528 93822 399537
rect 93766 399463 93822 399472
rect 92478 398032 92534 398041
rect 92478 397967 92534 397976
rect 92492 397594 92520 397967
rect 92480 397588 92532 397594
rect 92480 397530 92532 397536
rect 92664 397588 92716 397594
rect 92664 397530 92716 397536
rect 91928 396772 91980 396778
rect 91928 396714 91980 396720
rect 91836 394664 91888 394670
rect 91836 394606 91888 394612
rect 90928 393286 91048 393314
rect 90928 387190 90956 393286
rect 91940 390697 91968 396714
rect 91558 390688 91614 390697
rect 91558 390623 91614 390632
rect 91926 390688 91982 390697
rect 91926 390623 91982 390632
rect 91008 388000 91060 388006
rect 91008 387942 91060 387948
rect 90916 387184 90968 387190
rect 90916 387126 90968 387132
rect 90364 387116 90416 387122
rect 90364 387058 90416 387064
rect 91020 385914 91048 387942
rect 91572 385914 91600 390623
rect 87064 385886 87446 385914
rect 87708 385886 88090 385914
rect 88352 385886 88734 385914
rect 90022 385886 90312 385914
rect 90666 385886 91048 385914
rect 91310 385886 91600 385914
rect 92676 385778 92704 397530
rect 93872 396778 93900 438874
rect 94516 437442 94544 440028
rect 95160 438938 95188 440028
rect 96448 439210 96476 440028
rect 96436 439204 96488 439210
rect 96436 439146 96488 439152
rect 95148 438932 95200 438938
rect 95148 438874 95200 438880
rect 96448 438734 96476 439146
rect 97736 439074 97764 440028
rect 97724 439068 97776 439074
rect 97724 439010 97776 439016
rect 97736 438938 97764 439010
rect 96620 438932 96672 438938
rect 96620 438874 96672 438880
rect 97724 438932 97776 438938
rect 97724 438874 97776 438880
rect 96436 438728 96488 438734
rect 96436 438670 96488 438676
rect 94504 437436 94556 437442
rect 94504 437378 94556 437384
rect 93860 396772 93912 396778
rect 93860 396714 93912 396720
rect 92940 392080 92992 392086
rect 92940 392022 92992 392028
rect 92952 385914 92980 392022
rect 94516 391338 94544 437378
rect 96448 431954 96476 438670
rect 96448 431926 96568 431954
rect 96540 392766 96568 431926
rect 96632 402354 96660 438874
rect 98380 438326 98408 440028
rect 98368 438320 98420 438326
rect 98368 438262 98420 438268
rect 96620 402348 96672 402354
rect 96620 402290 96672 402296
rect 98656 399498 98684 440166
rect 99024 438802 99052 440028
rect 99012 438796 99064 438802
rect 99012 438738 99064 438744
rect 99288 438320 99340 438326
rect 99288 438262 99340 438268
rect 98644 399492 98696 399498
rect 98644 399434 98696 399440
rect 97908 395344 97960 395350
rect 97908 395286 97960 395292
rect 96528 392760 96580 392766
rect 96528 392702 96580 392708
rect 96252 392692 96304 392698
rect 96252 392634 96304 392640
rect 94504 391332 94556 391338
rect 94504 391274 94556 391280
rect 94136 391264 94188 391270
rect 94136 391206 94188 391212
rect 94148 385914 94176 391206
rect 95882 389192 95938 389201
rect 95882 389127 95938 389136
rect 94872 387116 94924 387122
rect 94872 387058 94924 387064
rect 94884 385914 94912 387058
rect 95896 385914 95924 389127
rect 92952 385886 93242 385914
rect 93886 385886 94176 385914
rect 94530 385886 94912 385914
rect 95818 385886 95924 385914
rect 92598 385750 92704 385778
rect 96264 385778 96292 392634
rect 97448 389972 97500 389978
rect 97448 389914 97500 389920
rect 96526 389872 96582 389881
rect 96526 389807 96582 389816
rect 96540 389201 96568 389807
rect 96526 389192 96582 389201
rect 96526 389127 96582 389136
rect 97460 385914 97488 389914
rect 97920 387818 97948 395286
rect 99300 392630 99328 438262
rect 99484 402974 99512 476303
rect 99760 475726 99788 538186
rect 100114 489968 100170 489977
rect 100114 489903 100170 489912
rect 100128 488345 100156 489903
rect 100114 488336 100170 488345
rect 100114 488271 100170 488280
rect 99748 475720 99800 475726
rect 99748 475662 99800 475668
rect 100024 447908 100076 447914
rect 100024 447850 100076 447856
rect 99746 443728 99802 443737
rect 99746 443663 99802 443672
rect 99668 438870 99696 440028
rect 99656 438864 99708 438870
rect 99656 438806 99708 438812
rect 99760 438598 99788 443663
rect 99748 438592 99800 438598
rect 99748 438534 99800 438540
rect 100036 437374 100064 447850
rect 100312 441153 100340 540138
rect 100956 537033 100984 540138
rect 102227 540110 102272 540138
rect 102046 537976 102102 537985
rect 102046 537911 102102 537920
rect 102060 537033 102088 537911
rect 102244 537810 102272 540110
rect 102232 537804 102284 537810
rect 102232 537746 102284 537752
rect 102888 537674 102916 540138
rect 103532 538218 103560 540138
rect 103520 538212 103572 538218
rect 103520 538154 103572 538160
rect 102876 537668 102928 537674
rect 102876 537610 102928 537616
rect 100942 537024 100998 537033
rect 100942 536959 100998 536968
rect 102046 537024 102102 537033
rect 102046 536959 102102 536968
rect 101956 535016 102008 535022
rect 101956 534958 102008 534964
rect 100668 491632 100720 491638
rect 100668 491574 100720 491580
rect 100680 491298 100708 491574
rect 100668 491292 100720 491298
rect 100668 491234 100720 491240
rect 101864 491156 101916 491162
rect 101864 491098 101916 491104
rect 101312 490680 101364 490686
rect 101312 490622 101364 490628
rect 101324 489870 101352 490622
rect 101876 489977 101904 491098
rect 101862 489968 101918 489977
rect 101862 489903 101864 489912
rect 101916 489903 101918 489912
rect 101864 489874 101916 489880
rect 101312 489864 101364 489870
rect 101876 489843 101904 489874
rect 101312 489806 101364 489812
rect 101324 485774 101352 489806
rect 101324 485746 101444 485774
rect 100668 477488 100720 477494
rect 100668 477430 100720 477436
rect 100680 476377 100708 477430
rect 100666 476368 100722 476377
rect 100666 476303 100722 476312
rect 100760 475720 100812 475726
rect 100760 475662 100812 475668
rect 100298 441144 100354 441153
rect 100298 441079 100354 441088
rect 100772 439793 100800 475662
rect 100850 451208 100906 451217
rect 100850 451143 100906 451152
rect 100864 450634 100892 451143
rect 100852 450628 100904 450634
rect 100852 450570 100904 450576
rect 100758 439784 100814 439793
rect 100758 439719 100814 439728
rect 100024 437368 100076 437374
rect 100024 437310 100076 437316
rect 100864 429894 100892 450570
rect 100852 429888 100904 429894
rect 100852 429830 100904 429836
rect 100668 422272 100720 422278
rect 100668 422214 100720 422220
rect 99392 402946 99512 402974
rect 99392 398274 99420 402946
rect 99380 398268 99432 398274
rect 99380 398210 99432 398216
rect 99392 398138 99420 398210
rect 99380 398132 99432 398138
rect 99380 398074 99432 398080
rect 99288 392624 99340 392630
rect 99194 392592 99250 392601
rect 99288 392566 99340 392572
rect 99194 392527 99250 392536
rect 98826 388376 98882 388385
rect 98826 388311 98882 388320
rect 98840 387870 98868 388311
rect 98828 387864 98880 387870
rect 97920 387790 98040 387818
rect 98828 387806 98880 387812
rect 97106 385886 97488 385914
rect 98012 385914 98040 387790
rect 99208 385914 99236 392527
rect 100680 391406 100708 422214
rect 101416 393514 101444 485746
rect 101968 478961 101996 534958
rect 101954 478952 102010 478961
rect 101954 478887 102010 478896
rect 102060 441833 102088 536959
rect 102140 494760 102192 494766
rect 102140 494702 102192 494708
rect 102152 449426 102180 494702
rect 102232 492176 102284 492182
rect 102232 492118 102284 492124
rect 102244 458402 102272 492118
rect 103336 488504 103388 488510
rect 103336 488446 103388 488452
rect 103348 487393 103376 488446
rect 103428 488436 103480 488442
rect 103428 488378 103480 488384
rect 103440 487937 103468 488378
rect 103426 487928 103482 487937
rect 103426 487863 103482 487872
rect 103520 487824 103572 487830
rect 103520 487766 103572 487772
rect 103334 487384 103390 487393
rect 103334 487319 103390 487328
rect 103426 486704 103482 486713
rect 103532 486690 103560 487766
rect 103482 486662 103560 486690
rect 103426 486639 103482 486648
rect 102322 485344 102378 485353
rect 102322 485279 102378 485288
rect 102336 485110 102364 485279
rect 102324 485104 102376 485110
rect 102324 485046 102376 485052
rect 102322 483848 102378 483857
rect 102322 483783 102378 483792
rect 102336 483682 102364 483783
rect 102324 483676 102376 483682
rect 102324 483618 102376 483624
rect 102416 482996 102468 483002
rect 102416 482938 102468 482944
rect 102324 482928 102376 482934
rect 102322 482896 102324 482905
rect 102376 482896 102378 482905
rect 102322 482831 102378 482840
rect 102428 482633 102456 482938
rect 102414 482624 102470 482633
rect 102414 482559 102470 482568
rect 102416 481636 102468 481642
rect 102416 481578 102468 481584
rect 102324 481568 102376 481574
rect 102322 481536 102324 481545
rect 102376 481536 102378 481545
rect 102322 481471 102378 481480
rect 102428 481273 102456 481578
rect 102414 481264 102470 481273
rect 102414 481199 102470 481208
rect 102324 480208 102376 480214
rect 102324 480150 102376 480156
rect 102336 479913 102364 480150
rect 102322 479904 102378 479913
rect 102322 479839 102378 479848
rect 103426 478136 103482 478145
rect 103426 478071 103482 478080
rect 102414 477864 102470 477873
rect 102414 477799 102470 477808
rect 102428 477562 102456 477799
rect 102416 477556 102468 477562
rect 102416 477498 102468 477504
rect 102506 477048 102562 477057
rect 102506 476983 102562 476992
rect 102322 476504 102378 476513
rect 102322 476439 102378 476448
rect 102336 476134 102364 476439
rect 102324 476128 102376 476134
rect 102324 476070 102376 476076
rect 102416 476060 102468 476066
rect 102416 476002 102468 476008
rect 102324 475992 102376 475998
rect 102324 475934 102376 475940
rect 102336 475697 102364 475934
rect 102322 475688 102378 475697
rect 102322 475623 102378 475632
rect 102428 475153 102456 476002
rect 102414 475144 102470 475153
rect 102414 475079 102470 475088
rect 102324 474700 102376 474706
rect 102324 474642 102376 474648
rect 102336 474337 102364 474642
rect 102322 474328 102378 474337
rect 102322 474263 102378 474272
rect 102520 474065 102548 476983
rect 102506 474056 102562 474065
rect 102506 473991 102562 474000
rect 102322 472968 102378 472977
rect 102322 472903 102378 472912
rect 102336 472802 102364 472903
rect 102324 472796 102376 472802
rect 102324 472738 102376 472744
rect 103440 472734 103468 478071
rect 103428 472728 103480 472734
rect 103428 472670 103480 472676
rect 102324 472660 102376 472666
rect 102324 472602 102376 472608
rect 102336 471753 102364 472602
rect 103440 472433 103468 472670
rect 103426 472424 103482 472433
rect 103426 472359 103482 472368
rect 102416 471980 102468 471986
rect 102416 471922 102468 471928
rect 102322 471744 102378 471753
rect 102322 471679 102378 471688
rect 102428 471073 102456 471922
rect 103426 471200 103482 471209
rect 103426 471135 103482 471144
rect 102414 471064 102470 471073
rect 102414 470999 102470 471008
rect 102784 470620 102836 470626
rect 102784 470562 102836 470568
rect 102796 469713 102824 470562
rect 103440 470257 103468 471135
rect 103426 470248 103482 470257
rect 103426 470183 103482 470192
rect 102782 469704 102838 469713
rect 102782 469639 102838 469648
rect 102324 469192 102376 469198
rect 102324 469134 102376 469140
rect 102336 468897 102364 469134
rect 102322 468888 102378 468897
rect 102322 468823 102378 468832
rect 103520 468512 103572 468518
rect 103520 468454 103572 468460
rect 102782 466984 102838 466993
rect 102782 466919 102838 466928
rect 102796 466478 102824 466919
rect 103426 466848 103482 466857
rect 103426 466783 103482 466792
rect 103440 466562 103468 466783
rect 103532 466562 103560 468454
rect 103440 466534 103560 466562
rect 102784 466472 102836 466478
rect 102784 466414 102836 466420
rect 102324 466404 102376 466410
rect 102324 466346 102376 466352
rect 102336 466177 102364 466346
rect 102322 466168 102378 466177
rect 102322 466103 102378 466112
rect 103426 465760 103482 465769
rect 103426 465695 103482 465704
rect 103440 465497 103468 465695
rect 103426 465488 103482 465497
rect 103426 465423 103482 465432
rect 102324 465044 102376 465050
rect 102324 464986 102376 464992
rect 102336 464273 102364 464986
rect 102414 464808 102470 464817
rect 102414 464743 102470 464752
rect 102322 464264 102378 464273
rect 102322 464199 102378 464208
rect 102428 463758 102456 464743
rect 102416 463752 102468 463758
rect 102416 463694 102468 463700
rect 102324 463684 102376 463690
rect 102324 463626 102376 463632
rect 102336 463457 102364 463626
rect 102322 463448 102378 463457
rect 102322 463383 102378 463392
rect 102324 462324 102376 462330
rect 102324 462266 102376 462272
rect 102336 462097 102364 462266
rect 102322 462088 102378 462097
rect 102322 462023 102378 462032
rect 102322 461408 102378 461417
rect 102322 461343 102378 461352
rect 102336 460970 102364 461343
rect 102324 460964 102376 460970
rect 102324 460906 102376 460912
rect 102324 460216 102376 460222
rect 102324 460158 102376 460164
rect 102874 460184 102930 460193
rect 102336 460057 102364 460158
rect 102874 460119 102930 460128
rect 102322 460048 102378 460057
rect 102322 459983 102378 459992
rect 102888 459610 102916 460119
rect 102876 459604 102928 459610
rect 102876 459546 102928 459552
rect 102324 459468 102376 459474
rect 102324 459410 102376 459416
rect 102336 459377 102364 459410
rect 102322 459368 102378 459377
rect 102322 459303 102378 459312
rect 102414 458688 102470 458697
rect 102414 458623 102470 458632
rect 102244 458374 102364 458402
rect 102230 456104 102286 456113
rect 102230 456039 102286 456048
rect 102244 455530 102272 456039
rect 102232 455524 102284 455530
rect 102232 455466 102284 455472
rect 102232 455388 102284 455394
rect 102232 455330 102284 455336
rect 102244 454753 102272 455330
rect 102230 454744 102286 454753
rect 102230 454679 102286 454688
rect 102232 454028 102284 454034
rect 102232 453970 102284 453976
rect 102244 453937 102272 453970
rect 102230 453928 102286 453937
rect 102230 453863 102286 453872
rect 102232 453416 102284 453422
rect 102232 453358 102284 453364
rect 102244 453257 102272 453358
rect 102230 453248 102286 453257
rect 102230 453183 102286 453192
rect 102232 452600 102284 452606
rect 102230 452568 102232 452577
rect 102284 452568 102286 452577
rect 102230 452503 102286 452512
rect 102152 449398 102272 449426
rect 102138 449304 102194 449313
rect 102138 449239 102140 449248
rect 102192 449239 102194 449248
rect 102140 449210 102192 449216
rect 102140 448520 102192 448526
rect 102138 448488 102140 448497
rect 102192 448488 102194 448497
rect 102138 448423 102194 448432
rect 102138 446312 102194 446321
rect 102138 446247 102194 446256
rect 102152 445874 102180 446247
rect 102140 445868 102192 445874
rect 102140 445810 102192 445816
rect 102046 441824 102102 441833
rect 102046 441759 102102 441768
rect 102046 440192 102102 440201
rect 102046 440127 102102 440136
rect 102060 438977 102088 440127
rect 102046 438968 102102 438977
rect 102046 438903 102102 438912
rect 101404 393508 101456 393514
rect 101404 393450 101456 393456
rect 100758 393408 100814 393417
rect 100758 393343 100814 393352
rect 100668 391400 100720 391406
rect 100668 391342 100720 391348
rect 100024 388068 100076 388074
rect 100024 388010 100076 388016
rect 100036 385914 100064 388010
rect 98012 385886 98394 385914
rect 99038 385886 99236 385914
rect 99682 385886 100064 385914
rect 100772 385914 100800 393343
rect 101416 389162 101444 393450
rect 102060 391338 102088 438903
rect 102244 438326 102272 449398
rect 102336 438530 102364 458374
rect 102428 458250 102456 458623
rect 102416 458244 102468 458250
rect 102416 458186 102468 458192
rect 102414 456648 102470 456657
rect 102414 456583 102470 456592
rect 102428 455462 102456 456583
rect 102416 455456 102468 455462
rect 102416 455398 102468 455404
rect 102416 449880 102468 449886
rect 102416 449822 102468 449828
rect 102428 449177 102456 449822
rect 102414 449168 102470 449177
rect 102414 449103 102470 449112
rect 102416 448452 102468 448458
rect 102416 448394 102468 448400
rect 102428 447953 102456 448394
rect 102414 447944 102470 447953
rect 102414 447879 102470 447888
rect 102600 445052 102652 445058
rect 102600 444994 102652 445000
rect 102612 443737 102640 444994
rect 102598 443728 102654 443737
rect 102598 443663 102654 443672
rect 102874 443048 102930 443057
rect 102874 442983 102930 442992
rect 102888 442882 102916 442983
rect 102876 442876 102928 442882
rect 102876 442818 102928 442824
rect 103334 441824 103390 441833
rect 103334 441759 103390 441768
rect 103348 441658 103376 441759
rect 103336 441652 103388 441658
rect 103336 441594 103388 441600
rect 102874 441144 102930 441153
rect 102874 441079 102930 441088
rect 102888 440298 102916 441079
rect 102876 440292 102928 440298
rect 102876 440234 102928 440240
rect 103058 439784 103114 439793
rect 103058 439719 103114 439728
rect 103072 439142 103100 439719
rect 103060 439136 103112 439142
rect 103060 439078 103112 439084
rect 102324 438524 102376 438530
rect 102324 438466 102376 438472
rect 102232 438320 102284 438326
rect 102232 438262 102284 438268
rect 103440 394097 103468 465423
rect 103520 458856 103572 458862
rect 103520 458798 103572 458804
rect 103532 458153 103560 458798
rect 103518 458144 103574 458153
rect 103518 458079 103574 458088
rect 103520 457156 103572 457162
rect 103520 457098 103572 457104
rect 103532 455433 103560 457098
rect 103518 455424 103574 455433
rect 103518 455359 103574 455368
rect 103520 451920 103572 451926
rect 103520 451862 103572 451868
rect 103532 450673 103560 451862
rect 104176 451274 104204 540138
rect 104716 538144 104768 538150
rect 104820 538121 104848 540138
rect 105478 540110 105584 540138
rect 104716 538086 104768 538092
rect 104806 538112 104862 538121
rect 104728 537849 104756 538086
rect 104806 538047 104862 538056
rect 104714 537840 104770 537849
rect 104714 537775 104770 537784
rect 105556 536897 105584 540110
rect 105542 536888 105598 536897
rect 105542 536823 105598 536832
rect 104254 491600 104310 491609
rect 104254 491535 104310 491544
rect 104268 489802 104296 491535
rect 104256 489796 104308 489802
rect 104256 489738 104308 489744
rect 104084 451246 104204 451274
rect 103518 450664 103574 450673
rect 103518 450599 103574 450608
rect 104084 445777 104112 451246
rect 104070 445768 104126 445777
rect 104070 445703 104126 445712
rect 104084 445233 104112 445703
rect 104070 445224 104126 445233
rect 104070 445159 104126 445168
rect 103520 445120 103572 445126
rect 103520 445062 103572 445068
rect 103532 444281 103560 445062
rect 104162 444408 104218 444417
rect 104162 444343 104218 444352
rect 103518 444272 103574 444281
rect 103518 444207 103574 444216
rect 104176 399566 104204 444343
rect 104164 399560 104216 399566
rect 104164 399502 104216 399508
rect 104268 394942 104296 489738
rect 105544 472252 105596 472258
rect 105544 472194 105596 472200
rect 105556 455530 105584 472194
rect 105544 455524 105596 455530
rect 105544 455466 105596 455472
rect 105556 451274 105584 455466
rect 105556 451246 105676 451274
rect 105544 445868 105596 445874
rect 105544 445810 105596 445816
rect 103704 394936 103756 394942
rect 103704 394878 103756 394884
rect 104256 394936 104308 394942
rect 104256 394878 104308 394884
rect 103426 394088 103482 394097
rect 103426 394023 103482 394032
rect 102048 391332 102100 391338
rect 102048 391274 102100 391280
rect 101404 389156 101456 389162
rect 101404 389098 101456 389104
rect 103612 389156 103664 389162
rect 103612 389098 103664 389104
rect 101864 388544 101916 388550
rect 101864 388486 101916 388492
rect 101876 385914 101904 388486
rect 103624 385914 103652 389098
rect 100772 385886 100970 385914
rect 101614 385886 101904 385914
rect 103546 385886 103652 385914
rect 103716 385914 103744 394878
rect 104532 389904 104584 389910
rect 104532 389846 104584 389852
rect 104544 385914 104572 389846
rect 105556 387258 105584 445810
rect 105648 396914 105676 451246
rect 105832 450634 105860 543759
rect 106094 540424 106150 540433
rect 106094 540359 106150 540368
rect 106108 536790 106136 540359
rect 106096 536784 106148 536790
rect 106096 536726 106148 536732
rect 106108 536110 106136 536726
rect 106096 536104 106148 536110
rect 106096 536046 106148 536052
rect 106200 460154 106228 552055
rect 106384 482934 106412 574631
rect 106476 486577 106504 578031
rect 107672 573345 107700 582694
rect 109130 582448 109186 582457
rect 109130 582383 109186 582392
rect 108946 580816 109002 580825
rect 108946 580751 109002 580760
rect 108854 580136 108910 580145
rect 108854 580071 108910 580080
rect 108868 579578 108896 580071
rect 108960 579698 108988 580751
rect 108948 579692 109000 579698
rect 108948 579634 109000 579640
rect 108868 579550 109080 579578
rect 108854 579456 108910 579465
rect 108854 579391 108910 579400
rect 108868 578338 108896 579391
rect 108946 578776 109002 578785
rect 108946 578711 109002 578720
rect 108856 578332 108908 578338
rect 108856 578274 108908 578280
rect 108960 578270 108988 578711
rect 108948 578264 109000 578270
rect 108948 578206 109000 578212
rect 108212 578196 108264 578202
rect 108212 578138 108264 578144
rect 108224 577561 108252 578138
rect 108210 577552 108266 577561
rect 108210 577487 108266 577496
rect 108854 576736 108910 576745
rect 108854 576671 108910 576680
rect 108868 575550 108896 576671
rect 108946 576056 109002 576065
rect 108946 575991 109002 576000
rect 108960 575618 108988 575991
rect 108948 575612 109000 575618
rect 108948 575554 109000 575560
rect 108856 575544 108908 575550
rect 108856 575486 108908 575492
rect 108948 574048 109000 574054
rect 108946 574016 108948 574025
rect 109000 574016 109002 574025
rect 108946 573951 109002 573960
rect 107658 573336 107714 573345
rect 107658 573271 107714 573280
rect 107842 573336 107898 573345
rect 107842 573271 107898 573280
rect 107856 572830 107884 573271
rect 108948 572892 109000 572898
rect 108948 572834 109000 572840
rect 107844 572824 107896 572830
rect 108960 572801 108988 572834
rect 107844 572766 107896 572772
rect 108946 572792 109002 572801
rect 108946 572727 109002 572736
rect 108946 571976 109002 571985
rect 108946 571911 109002 571920
rect 107934 571432 107990 571441
rect 108960 571402 108988 571911
rect 107934 571367 107990 571376
rect 108948 571396 109000 571402
rect 107750 563136 107806 563145
rect 107750 563071 107806 563080
rect 107658 560416 107714 560425
rect 107658 560351 107660 560360
rect 107712 560351 107714 560360
rect 107660 560322 107712 560328
rect 107658 556336 107714 556345
rect 107658 556271 107714 556280
rect 106922 551576 106978 551585
rect 106922 551511 106978 551520
rect 106936 528630 106964 551511
rect 107672 548282 107700 556271
rect 107660 548276 107712 548282
rect 107660 548218 107712 548224
rect 107658 542736 107714 542745
rect 107658 542671 107714 542680
rect 107566 540152 107622 540161
rect 107566 540087 107622 540096
rect 106924 528624 106976 528630
rect 106924 528566 106976 528572
rect 106462 486568 106518 486577
rect 106462 486503 106518 486512
rect 106372 482928 106424 482934
rect 106372 482870 106424 482876
rect 107476 482928 107528 482934
rect 107476 482870 107528 482876
rect 107488 482322 107516 482870
rect 107476 482316 107528 482322
rect 107476 482258 107528 482264
rect 107476 477624 107528 477630
rect 107476 477566 107528 477572
rect 107384 474768 107436 474774
rect 107384 474710 107436 474716
rect 107396 471986 107424 474710
rect 107384 471980 107436 471986
rect 107384 471922 107436 471928
rect 107396 471034 107424 471922
rect 107384 471028 107436 471034
rect 107384 470970 107436 470976
rect 107016 469872 107068 469878
rect 107016 469814 107068 469820
rect 106188 460148 106240 460154
rect 106188 460090 106240 460096
rect 106188 459536 106240 459542
rect 106188 459478 106240 459484
rect 106094 456784 106150 456793
rect 106094 456719 106150 456728
rect 106108 453422 106136 456719
rect 106096 453416 106148 453422
rect 106096 453358 106148 453364
rect 106200 451274 106228 459478
rect 106108 451246 106228 451274
rect 105820 450628 105872 450634
rect 105820 450570 105872 450576
rect 105728 447840 105780 447846
rect 105728 447782 105780 447788
rect 105740 440230 105768 447782
rect 106108 443698 106136 451246
rect 106188 449200 106240 449206
rect 106188 449142 106240 449148
rect 106200 448526 106228 449142
rect 106924 448588 106976 448594
rect 106924 448530 106976 448536
rect 106188 448520 106240 448526
rect 106188 448462 106240 448468
rect 106096 443692 106148 443698
rect 106096 443634 106148 443640
rect 105728 440224 105780 440230
rect 105728 440166 105780 440172
rect 106936 398138 106964 448530
rect 107028 438666 107056 469814
rect 107488 465050 107516 477566
rect 107476 465044 107528 465050
rect 107476 464986 107528 464992
rect 107580 460934 107608 540087
rect 107396 460906 107608 460934
rect 107396 448662 107424 460906
rect 107566 456104 107622 456113
rect 107566 456039 107622 456048
rect 107580 455394 107608 456039
rect 107568 455388 107620 455394
rect 107568 455330 107620 455336
rect 107672 451274 107700 542671
rect 107764 474774 107792 563071
rect 107842 548856 107898 548865
rect 107842 548791 107898 548800
rect 107856 548418 107884 548791
rect 107844 548412 107896 548418
rect 107844 548354 107896 548360
rect 107844 548276 107896 548282
rect 107844 548218 107896 548224
rect 107856 477630 107884 548218
rect 107948 535022 107976 571367
rect 108948 571338 109000 571344
rect 108854 570616 108910 570625
rect 108854 570551 108910 570560
rect 108868 570042 108896 570551
rect 108946 570072 109002 570081
rect 108856 570036 108908 570042
rect 108946 570007 109002 570016
rect 108856 569978 108908 569984
rect 108960 569974 108988 570007
rect 108948 569968 109000 569974
rect 108948 569910 109000 569916
rect 108946 569256 109002 569265
rect 108946 569191 109002 569200
rect 108960 568614 108988 569191
rect 108948 568608 109000 568614
rect 108948 568550 109000 568556
rect 108946 567896 109002 567905
rect 108946 567831 109002 567840
rect 108960 567594 108988 567831
rect 108948 567588 109000 567594
rect 108948 567530 109000 567536
rect 108948 567248 109000 567254
rect 108946 567216 108948 567225
rect 109000 567216 109002 567225
rect 108946 567151 109002 567160
rect 108854 566536 108910 566545
rect 108854 566471 108910 566480
rect 108868 565962 108896 566471
rect 108856 565956 108908 565962
rect 108856 565898 108908 565904
rect 108948 565888 109000 565894
rect 108946 565856 108948 565865
rect 109000 565856 109002 565865
rect 108946 565791 109002 565800
rect 108946 565176 109002 565185
rect 108946 565111 109002 565120
rect 108960 564466 108988 565111
rect 108948 564460 109000 564466
rect 108948 564402 109000 564408
rect 108946 563816 109002 563825
rect 108946 563751 108948 563760
rect 109000 563751 109002 563760
rect 108948 563722 109000 563728
rect 108946 561096 109002 561105
rect 108946 561031 109002 561040
rect 108960 560318 108988 561031
rect 108948 560312 109000 560318
rect 108948 560254 109000 560260
rect 108854 559736 108910 559745
rect 108854 559671 108910 559680
rect 108868 559026 108896 559671
rect 108946 559056 109002 559065
rect 108856 559020 108908 559026
rect 108946 558991 109002 559000
rect 108856 558962 108908 558968
rect 108960 558958 108988 558991
rect 108948 558952 109000 558958
rect 108948 558894 109000 558900
rect 108578 558376 108634 558385
rect 108578 558311 108634 558320
rect 108592 558074 108620 558311
rect 108580 558068 108632 558074
rect 108580 558010 108632 558016
rect 108946 557016 109002 557025
rect 108946 556951 109002 556960
rect 108960 556578 108988 556951
rect 108948 556572 109000 556578
rect 108948 556514 109000 556520
rect 108946 554296 109002 554305
rect 108946 554231 109002 554240
rect 108960 554062 108988 554231
rect 108948 554056 109000 554062
rect 108948 553998 109000 554004
rect 108946 553616 109002 553625
rect 108946 553551 109002 553560
rect 108960 553450 108988 553551
rect 108948 553444 109000 553450
rect 108948 553386 109000 553392
rect 108946 552936 109002 552945
rect 108946 552871 109002 552880
rect 108960 552090 108988 552871
rect 108948 552084 109000 552090
rect 108948 552026 109000 552032
rect 108946 550896 109002 550905
rect 108946 550831 109002 550840
rect 108960 550662 108988 550831
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108854 550216 108910 550225
rect 108854 550151 108910 550160
rect 108868 549302 108896 550151
rect 108946 549536 109002 549545
rect 108946 549471 109002 549480
rect 108960 549370 108988 549471
rect 108948 549364 109000 549370
rect 108948 549306 109000 549312
rect 108856 549296 108908 549302
rect 108856 549238 108908 549244
rect 108946 547496 109002 547505
rect 108946 547431 109002 547440
rect 108960 546514 108988 547431
rect 108948 546508 109000 546514
rect 108948 546450 109000 546456
rect 108946 546136 109002 546145
rect 108946 546071 109002 546080
rect 108960 545766 108988 546071
rect 108948 545760 109000 545766
rect 108948 545702 109000 545708
rect 108946 545456 109002 545465
rect 108946 545391 109002 545400
rect 108960 545154 108988 545391
rect 108948 545148 109000 545154
rect 108948 545090 109000 545096
rect 108946 544776 109002 544785
rect 108946 544711 109002 544720
rect 108960 544406 108988 544711
rect 108948 544400 109000 544406
rect 108948 544342 109000 544348
rect 108946 543416 109002 543425
rect 108946 543351 109002 543360
rect 108960 542434 108988 543351
rect 108948 542428 109000 542434
rect 108948 542370 109000 542376
rect 108946 542056 109002 542065
rect 108946 541991 109002 542000
rect 108960 541006 108988 541991
rect 108948 541000 109000 541006
rect 108948 540942 109000 540948
rect 107936 535016 107988 535022
rect 107936 534958 107988 534964
rect 109052 488442 109080 579550
rect 109144 491858 109172 582383
rect 109224 572348 109276 572354
rect 109224 572290 109276 572296
rect 109236 555801 109264 572290
rect 110340 563786 110368 702714
rect 111708 702636 111760 702642
rect 111708 702578 111760 702584
rect 111616 590708 111668 590714
rect 111616 590650 111668 590656
rect 110696 583840 110748 583846
rect 110696 583782 110748 583788
rect 110512 572824 110564 572830
rect 110512 572766 110564 572772
rect 110328 563780 110380 563786
rect 110328 563722 110380 563728
rect 109222 555792 109278 555801
rect 109222 555727 109278 555736
rect 109236 554810 109264 555727
rect 109224 554804 109276 554810
rect 109224 554746 109276 554752
rect 109684 546576 109736 546582
rect 109684 546518 109736 546524
rect 109696 538218 109724 546518
rect 109776 541680 109828 541686
rect 109776 541622 109828 541628
rect 109684 538212 109736 538218
rect 109684 538154 109736 538160
rect 109788 537985 109816 541622
rect 109774 537976 109830 537985
rect 109774 537911 109830 537920
rect 109224 532228 109276 532234
rect 109224 532170 109276 532176
rect 109236 499574 109264 532170
rect 109236 499546 109448 499574
rect 109144 491830 109356 491858
rect 109132 491564 109184 491570
rect 109132 491506 109184 491512
rect 109144 491230 109172 491506
rect 109132 491224 109184 491230
rect 109132 491166 109184 491172
rect 109328 491162 109356 491830
rect 109316 491156 109368 491162
rect 109316 491098 109368 491104
rect 109420 489914 109448 499546
rect 110420 495508 110472 495514
rect 110420 495450 110472 495456
rect 109684 490612 109736 490618
rect 109684 490554 109736 490560
rect 109236 489886 109448 489914
rect 109040 488436 109092 488442
rect 109040 488378 109092 488384
rect 109052 487898 109080 488378
rect 109130 488336 109186 488345
rect 109130 488271 109186 488280
rect 109040 487892 109092 487898
rect 109040 487834 109092 487840
rect 107844 477624 107896 477630
rect 107844 477566 107896 477572
rect 108396 476196 108448 476202
rect 108396 476138 108448 476144
rect 107752 474768 107804 474774
rect 107752 474710 107804 474716
rect 108304 471028 108356 471034
rect 108304 470970 108356 470976
rect 107752 458924 107804 458930
rect 107752 458866 107804 458872
rect 107764 457162 107792 458866
rect 107752 457156 107804 457162
rect 107752 457098 107804 457104
rect 107580 451246 107700 451274
rect 107580 450650 107608 451246
rect 107488 450622 107608 450650
rect 107488 449274 107516 450622
rect 107568 450560 107620 450566
rect 107568 450502 107620 450508
rect 107580 449886 107608 450502
rect 107568 449880 107620 449886
rect 107568 449822 107620 449828
rect 107476 449268 107528 449274
rect 107476 449210 107528 449216
rect 107384 448656 107436 448662
rect 107384 448598 107436 448604
rect 107396 448458 107424 448598
rect 107488 448594 107516 449210
rect 107476 448588 107528 448594
rect 107476 448530 107528 448536
rect 107384 448452 107436 448458
rect 107384 448394 107436 448400
rect 107016 438660 107068 438666
rect 107016 438602 107068 438608
rect 108316 402422 108344 470970
rect 108408 439074 108436 476138
rect 109144 467945 109172 488271
rect 109236 476202 109264 489886
rect 109224 476196 109276 476202
rect 109224 476138 109276 476144
rect 109130 467936 109186 467945
rect 109130 467871 109186 467880
rect 108488 458176 108540 458182
rect 108488 458118 108540 458124
rect 108396 439068 108448 439074
rect 108396 439010 108448 439016
rect 108500 438938 108528 458118
rect 108488 438932 108540 438938
rect 108488 438874 108540 438880
rect 108304 402416 108356 402422
rect 108304 402358 108356 402364
rect 108856 401668 108908 401674
rect 108856 401610 108908 401616
rect 106924 398132 106976 398138
rect 106924 398074 106976 398080
rect 105636 396908 105688 396914
rect 105636 396850 105688 396856
rect 106280 389292 106332 389298
rect 106280 389234 106332 389240
rect 106292 387818 106320 389234
rect 107016 388476 107068 388482
rect 107016 388418 107068 388424
rect 106200 387790 106320 387818
rect 105544 387252 105596 387258
rect 105544 387194 105596 387200
rect 106200 385914 106228 387790
rect 107028 385914 107056 388418
rect 108868 387122 108896 401610
rect 108948 389904 109000 389910
rect 108948 389846 109000 389852
rect 108856 387116 108908 387122
rect 108856 387058 108908 387064
rect 108960 385914 108988 389846
rect 109696 388142 109724 490554
rect 110326 490512 110382 490521
rect 110326 490447 110382 490456
rect 110340 489734 110368 490447
rect 110328 489728 110380 489734
rect 110328 489670 110380 489676
rect 109684 388136 109736 388142
rect 109684 388078 109736 388084
rect 109696 385914 109724 388078
rect 110340 386442 110368 489670
rect 110432 393990 110460 495450
rect 110524 481574 110552 572766
rect 110604 548412 110656 548418
rect 110604 548354 110656 548360
rect 110512 481568 110564 481574
rect 110512 481510 110564 481516
rect 110616 472258 110644 548354
rect 110708 493474 110736 583782
rect 111628 554062 111656 590650
rect 111720 578241 111748 702578
rect 111800 587172 111852 587178
rect 111800 587114 111852 587120
rect 111706 578232 111762 578241
rect 111706 578167 111708 578176
rect 111760 578167 111762 578176
rect 111708 578138 111760 578144
rect 111720 578107 111748 578138
rect 111616 554056 111668 554062
rect 111616 553998 111668 554004
rect 111812 537849 111840 587114
rect 111984 581800 112036 581806
rect 111984 581742 112036 581748
rect 111892 558068 111944 558074
rect 111892 558010 111944 558016
rect 111798 537840 111854 537849
rect 111798 537775 111854 537784
rect 111812 536586 111840 537775
rect 111800 536580 111852 536586
rect 111800 536522 111852 536528
rect 111800 532092 111852 532098
rect 111800 532034 111852 532040
rect 110696 493468 110748 493474
rect 110696 493410 110748 493416
rect 111064 492108 111116 492114
rect 111064 492050 111116 492056
rect 110604 472252 110656 472258
rect 110604 472194 110656 472200
rect 110420 393984 110472 393990
rect 110418 393952 110420 393961
rect 110472 393952 110474 393961
rect 110418 393887 110474 393896
rect 110420 392828 110472 392834
rect 110420 392770 110472 392776
rect 110432 392018 110460 392770
rect 111076 392018 111104 492050
rect 111708 481568 111760 481574
rect 111708 481510 111760 481516
rect 111720 480962 111748 481510
rect 111708 480956 111760 480962
rect 111708 480898 111760 480904
rect 111708 478304 111760 478310
rect 111708 478246 111760 478252
rect 110420 392012 110472 392018
rect 110420 391954 110472 391960
rect 110972 392012 111024 392018
rect 110972 391954 111024 391960
rect 111064 392012 111116 392018
rect 111064 391954 111116 391960
rect 110328 386436 110380 386442
rect 110328 386378 110380 386384
rect 110340 385914 110368 386378
rect 103716 385886 104190 385914
rect 104544 385886 104834 385914
rect 106122 385886 106228 385914
rect 106766 385886 107056 385914
rect 108698 385886 108988 385914
rect 109342 385886 109724 385914
rect 109986 385886 110368 385914
rect 110984 385914 111012 391954
rect 111720 388482 111748 478246
rect 111812 436082 111840 532034
rect 111904 466410 111932 558010
rect 111996 539102 112024 581742
rect 113100 544406 113128 702850
rect 115848 702704 115900 702710
rect 115848 702646 115900 702652
rect 113180 584044 113232 584050
rect 113180 583986 113232 583992
rect 113088 544400 113140 544406
rect 113088 544342 113140 544348
rect 111984 539096 112036 539102
rect 111984 539038 112036 539044
rect 111984 534880 112036 534886
rect 111984 534822 112036 534828
rect 111892 466404 111944 466410
rect 111892 466346 111944 466352
rect 111996 466313 112024 534822
rect 112076 494896 112128 494902
rect 112076 494838 112128 494844
rect 111982 466304 112038 466313
rect 111982 466239 112038 466248
rect 112088 447914 112116 494838
rect 113192 489734 113220 583986
rect 114560 583976 114612 583982
rect 114560 583918 114612 583924
rect 113364 572892 113416 572898
rect 113364 572834 113416 572840
rect 113272 556572 113324 556578
rect 113272 556514 113324 556520
rect 113180 489728 113232 489734
rect 113180 489670 113232 489676
rect 112168 485104 112220 485110
rect 112166 485072 112168 485081
rect 112220 485072 112222 485081
rect 112166 485007 112222 485016
rect 113086 485072 113142 485081
rect 113086 485007 113142 485016
rect 113100 484430 113128 485007
rect 113088 484424 113140 484430
rect 113088 484366 113140 484372
rect 112352 466404 112404 466410
rect 112352 466346 112404 466352
rect 112364 465730 112392 466346
rect 112352 465724 112404 465730
rect 112352 465666 112404 465672
rect 113088 463752 113140 463758
rect 113088 463694 113140 463700
rect 113284 463694 113312 556514
rect 113376 481642 113404 572834
rect 114572 494766 114600 583918
rect 114652 567588 114704 567594
rect 114652 567530 114704 567536
rect 114560 494760 114612 494766
rect 114560 494702 114612 494708
rect 114560 492788 114612 492794
rect 114560 492730 114612 492736
rect 113456 491972 113508 491978
rect 113456 491914 113508 491920
rect 113364 481636 113416 481642
rect 113364 481578 113416 481584
rect 113100 463666 113312 463694
rect 112076 447908 112128 447914
rect 112076 447850 112128 447856
rect 111800 436076 111852 436082
rect 111800 436018 111852 436024
rect 113100 393314 113128 463666
rect 113468 401674 113496 491914
rect 114466 488744 114522 488753
rect 114466 488679 114522 488688
rect 114480 488442 114508 488679
rect 114468 488436 114520 488442
rect 114468 488378 114520 488384
rect 113456 401668 113508 401674
rect 113456 401610 113508 401616
rect 113822 401296 113878 401305
rect 113822 401231 113878 401240
rect 113008 393286 113128 393314
rect 112076 392012 112128 392018
rect 112076 391954 112128 391960
rect 111708 388476 111760 388482
rect 111708 388418 111760 388424
rect 112088 387870 112116 391954
rect 112076 387864 112128 387870
rect 112076 387806 112128 387812
rect 112088 385914 112116 387806
rect 112904 386504 112956 386510
rect 112904 386446 112956 386452
rect 112916 385914 112944 386446
rect 110984 385886 111274 385914
rect 111918 385886 112116 385914
rect 112562 385886 112944 385914
rect 96264 385750 96462 385778
rect 113008 385762 113036 393286
rect 113088 392488 113140 392494
rect 113088 392430 113140 392436
rect 113100 388550 113128 392430
rect 113836 392018 113864 401231
rect 114480 393314 114508 488378
rect 114388 393286 114508 393314
rect 113824 392012 113876 392018
rect 113824 391954 113876 391960
rect 113836 389174 113864 391954
rect 114388 389230 114416 393286
rect 114572 392494 114600 492730
rect 114664 477494 114692 567530
rect 115204 554804 115256 554810
rect 115204 554746 115256 554752
rect 114744 536580 114796 536586
rect 114744 536522 114796 536528
rect 114756 485774 114784 536522
rect 114756 485746 114876 485774
rect 114652 477488 114704 477494
rect 114652 477430 114704 477436
rect 114652 460964 114704 460970
rect 114652 460906 114704 460912
rect 114664 459785 114692 460906
rect 114650 459776 114706 459785
rect 114650 459711 114706 459720
rect 114848 458182 114876 485746
rect 115216 463690 115244 554746
rect 115860 545766 115888 702646
rect 116308 584452 116360 584458
rect 116308 584394 116360 584400
rect 116124 582480 116176 582486
rect 116124 582422 116176 582428
rect 115940 567248 115992 567254
rect 115940 567190 115992 567196
rect 115848 545760 115900 545766
rect 115848 545702 115900 545708
rect 115952 475998 115980 567190
rect 116136 534954 116164 582422
rect 116124 534948 116176 534954
rect 116124 534890 116176 534896
rect 116216 528624 116268 528630
rect 116216 528566 116268 528572
rect 116032 493400 116084 493406
rect 116032 493342 116084 493348
rect 116044 478310 116072 493342
rect 116124 487892 116176 487898
rect 116124 487834 116176 487840
rect 116032 478304 116084 478310
rect 116032 478246 116084 478252
rect 116032 477556 116084 477562
rect 116032 477498 116084 477504
rect 116044 477465 116072 477498
rect 116030 477456 116086 477465
rect 116030 477391 116086 477400
rect 116032 476128 116084 476134
rect 116032 476070 116084 476076
rect 115940 475992 115992 475998
rect 115938 475960 115940 475969
rect 115992 475960 115994 475969
rect 115938 475895 115994 475904
rect 115204 463684 115256 463690
rect 115204 463626 115256 463632
rect 115480 460284 115532 460290
rect 115480 460226 115532 460232
rect 115296 460148 115348 460154
rect 115296 460090 115348 460096
rect 115202 458280 115258 458289
rect 115202 458215 115204 458224
rect 115256 458215 115258 458224
rect 115204 458186 115256 458192
rect 114836 458176 114888 458182
rect 114836 458118 114888 458124
rect 114560 392488 114612 392494
rect 114560 392430 114612 392436
rect 114376 389224 114428 389230
rect 113836 389146 113956 389174
rect 113088 388544 113140 388550
rect 113088 388486 113140 388492
rect 113088 387932 113140 387938
rect 113088 387874 113140 387880
rect 113100 387326 113128 387874
rect 113088 387320 113140 387326
rect 113088 387262 113140 387268
rect 113928 385914 113956 389146
rect 113850 385886 113956 385914
rect 114296 389172 114376 389174
rect 114296 389166 114428 389172
rect 114926 389192 114982 389201
rect 114296 389146 114416 389166
rect 114296 385778 114324 389146
rect 114388 389101 114416 389146
rect 114926 389127 114982 389136
rect 114940 385914 114968 389127
rect 114940 385886 115138 385914
rect 112996 385756 113048 385762
rect 114296 385750 114494 385778
rect 112996 385698 113048 385704
rect 86316 385620 86368 385626
rect 86316 385562 86368 385568
rect 77496 385354 77892 385370
rect 77484 385348 77892 385354
rect 77536 385342 77892 385348
rect 102258 385354 102640 385370
rect 107410 385354 107608 385370
rect 102258 385348 102652 385354
rect 102258 385342 102600 385348
rect 77484 385290 77536 385296
rect 107410 385348 107620 385354
rect 107410 385342 107568 385348
rect 102600 385290 102652 385296
rect 107568 385290 107620 385296
rect 70308 378820 70360 378826
rect 70308 378762 70360 378768
rect 69308 364306 69704 364334
rect 69204 361616 69256 361622
rect 69204 361558 69256 361564
rect 69216 360913 69244 361558
rect 69202 360904 69258 360913
rect 69202 360839 69258 360848
rect 69110 356960 69166 356969
rect 69110 356895 69166 356904
rect 69478 356960 69534 356969
rect 69478 356895 69534 356904
rect 69492 356114 69520 356895
rect 69480 356108 69532 356114
rect 69480 356050 69532 356056
rect 68742 352472 68798 352481
rect 68742 352407 68798 352416
rect 67730 351520 67786 351529
rect 67730 351455 67786 351464
rect 68282 351520 68338 351529
rect 68282 351455 68338 351464
rect 67744 351218 67772 351455
rect 67732 351212 67784 351218
rect 67732 351154 67784 351160
rect 67638 349888 67694 349897
rect 67638 349823 67694 349832
rect 68008 349852 68060 349858
rect 67652 349178 67680 349823
rect 68008 349794 68060 349800
rect 68020 349761 68048 349794
rect 68006 349752 68062 349761
rect 68006 349687 68062 349696
rect 67640 349172 67692 349178
rect 67640 349114 67692 349120
rect 68558 347168 68614 347177
rect 68558 347103 68614 347112
rect 68572 347070 68600 347103
rect 68560 347064 68612 347070
rect 68560 347006 68612 347012
rect 67638 346760 67694 346769
rect 67638 346695 67694 346704
rect 67652 346458 67680 346695
rect 67640 346452 67692 346458
rect 67640 346394 67692 346400
rect 67652 345030 67680 346394
rect 67730 345672 67786 345681
rect 67730 345607 67786 345616
rect 67744 345098 67772 345607
rect 67732 345092 67784 345098
rect 67732 345034 67784 345040
rect 67640 345024 67692 345030
rect 68572 345014 68600 347006
rect 68572 344986 68692 345014
rect 67640 344966 67692 344972
rect 67730 344448 67786 344457
rect 67730 344383 67786 344392
rect 67638 343768 67694 343777
rect 67744 343738 67772 344383
rect 67638 343703 67694 343712
rect 67732 343732 67784 343738
rect 67652 343670 67680 343703
rect 67732 343674 67784 343680
rect 67640 343664 67692 343670
rect 67640 343606 67692 343612
rect 67638 341728 67694 341737
rect 67638 341663 67694 341672
rect 67546 341592 67602 341601
rect 67546 341527 67602 341536
rect 67652 340950 67680 341663
rect 67640 340944 67692 340950
rect 67640 340886 67692 340892
rect 68664 334801 68692 344986
rect 68650 334792 68706 334801
rect 68650 334727 68706 334736
rect 68756 333305 68784 352407
rect 68926 349752 68982 349761
rect 68926 349687 68982 349696
rect 68848 348430 68876 348461
rect 68836 348424 68888 348430
rect 68834 348392 68836 348401
rect 68888 348392 68890 348401
rect 68834 348327 68890 348336
rect 68742 333296 68798 333305
rect 68742 333231 68798 333240
rect 67456 331900 67508 331906
rect 67456 331842 67508 331848
rect 68848 327758 68876 348327
rect 68836 327752 68888 327758
rect 68836 327694 68888 327700
rect 68652 326528 68704 326534
rect 68652 326470 68704 326476
rect 66904 322244 66956 322250
rect 66904 322186 66956 322192
rect 66166 320784 66222 320793
rect 66166 320719 66222 320728
rect 67548 318232 67600 318238
rect 67548 318174 67600 318180
rect 66168 303748 66220 303754
rect 66168 303690 66220 303696
rect 65984 302932 66036 302938
rect 65984 302874 66036 302880
rect 66180 289814 66208 303690
rect 67560 291122 67588 318174
rect 67638 291136 67694 291145
rect 67560 291094 67638 291122
rect 67638 291071 67694 291080
rect 67652 290494 67680 291071
rect 67640 290488 67692 290494
rect 67640 290430 67692 290436
rect 66168 289808 66220 289814
rect 66168 289750 66220 289756
rect 68192 289808 68244 289814
rect 68192 289750 68244 289756
rect 68204 289513 68232 289750
rect 68190 289504 68246 289513
rect 68190 289439 68246 289448
rect 67640 288380 67692 288386
rect 67640 288322 67692 288328
rect 67652 288153 67680 288322
rect 67638 288144 67694 288153
rect 67638 288079 67694 288088
rect 66902 287464 66958 287473
rect 66902 287399 66958 287408
rect 66076 271924 66128 271930
rect 66076 271866 66128 271872
rect 65984 258188 66036 258194
rect 65984 258130 66036 258136
rect 65892 247172 65944 247178
rect 65892 247114 65944 247120
rect 64788 244996 64840 245002
rect 64788 244938 64840 244944
rect 64800 236706 64828 244938
rect 64788 236700 64840 236706
rect 64788 236642 64840 236648
rect 65904 182986 65932 247114
rect 65996 239562 66024 258130
rect 65984 239556 66036 239562
rect 65984 239498 66036 239504
rect 66088 227089 66116 271866
rect 66916 244662 66944 287399
rect 68282 286512 68338 286521
rect 68282 286447 68338 286456
rect 67638 284472 67694 284481
rect 67638 284407 67694 284416
rect 67652 284374 67680 284407
rect 67640 284368 67692 284374
rect 67640 284310 67692 284316
rect 67732 284300 67784 284306
rect 67732 284242 67784 284248
rect 67744 283393 67772 284242
rect 67730 283384 67786 283393
rect 67730 283319 67786 283328
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 282169 67680 282814
rect 67638 282160 67694 282169
rect 67638 282095 67694 282104
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67640 280084 67692 280090
rect 67640 280026 67692 280032
rect 67652 279313 67680 280026
rect 67744 279993 67772 280094
rect 67730 279984 67786 279993
rect 67730 279919 67786 279928
rect 67638 279304 67694 279313
rect 67638 279239 67694 279248
rect 67730 277808 67786 277817
rect 67730 277743 67786 277752
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277506 67680 277607
rect 67640 277500 67692 277506
rect 67640 277442 67692 277448
rect 67744 277438 67772 277743
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67638 276448 67694 276457
rect 67638 276383 67694 276392
rect 67652 276078 67680 276383
rect 67640 276072 67692 276078
rect 67640 276014 67692 276020
rect 67822 275088 67878 275097
rect 67822 275023 67878 275032
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274786 67680 274887
rect 67640 274780 67692 274786
rect 67640 274722 67692 274728
rect 67836 274718 67864 275023
rect 67824 274712 67876 274718
rect 67824 274654 67876 274660
rect 67732 274644 67784 274650
rect 67732 274586 67784 274592
rect 67744 274553 67772 274586
rect 67730 274544 67786 274553
rect 67730 274479 67786 274488
rect 67638 273592 67694 273601
rect 67638 273527 67694 273536
rect 67652 273290 67680 273527
rect 67640 273284 67692 273290
rect 67640 273226 67692 273232
rect 67638 272232 67694 272241
rect 67638 272167 67694 272176
rect 67546 271960 67602 271969
rect 67652 271930 67680 272167
rect 67546 271895 67602 271904
rect 67640 271924 67692 271930
rect 67456 248940 67508 248946
rect 67456 248882 67508 248888
rect 66904 244656 66956 244662
rect 66904 244598 66956 244604
rect 67364 244384 67416 244390
rect 67364 244326 67416 244332
rect 66168 242956 66220 242962
rect 66168 242898 66220 242904
rect 66180 233918 66208 242898
rect 66168 233912 66220 233918
rect 66168 233854 66220 233860
rect 66074 227080 66130 227089
rect 66074 227015 66130 227024
rect 65892 182980 65944 182986
rect 65892 182922 65944 182928
rect 67376 182889 67404 244326
rect 67362 182880 67418 182889
rect 67362 182815 67418 182824
rect 67468 180033 67496 248882
rect 67560 196790 67588 271895
rect 67640 271866 67692 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271008 67694 271017
rect 67638 270943 67694 270952
rect 67652 270570 67680 270943
rect 67744 270881 67772 271798
rect 67730 270872 67786 270881
rect 67730 270807 67786 270816
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67730 269648 67786 269657
rect 67730 269583 67786 269592
rect 67638 269512 67694 269521
rect 67638 269447 67694 269456
rect 67652 269142 67680 269447
rect 67744 269210 67772 269583
rect 67732 269204 67784 269210
rect 67732 269146 67784 269152
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67640 268388 67692 268394
rect 67640 268330 67692 268336
rect 67652 268161 67680 268330
rect 67638 268152 67694 268161
rect 67638 268087 67694 268096
rect 67640 267708 67692 267714
rect 67640 267650 67692 267656
rect 67652 267481 67680 267650
rect 67732 267640 67784 267646
rect 67732 267582 67784 267588
rect 67638 267472 67694 267481
rect 67638 267407 67694 267416
rect 67744 267073 67772 267582
rect 67730 267064 67786 267073
rect 67730 266999 67786 267008
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265033 67680 266290
rect 67638 265024 67694 265033
rect 67638 264959 67694 264968
rect 67640 264920 67692 264926
rect 67638 264888 67640 264897
rect 67692 264888 67694 264897
rect 67638 264823 67694 264832
rect 67730 263664 67786 263673
rect 67730 263599 67732 263608
rect 67784 263599 67786 263608
rect 67732 263570 67784 263576
rect 67640 263560 67692 263566
rect 67638 263528 67640 263537
rect 67692 263528 67694 263537
rect 67638 263463 67694 263472
rect 67638 262304 67694 262313
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67638 261488 67694 261497
rect 67638 261423 67694 261432
rect 67652 260982 67680 261423
rect 67640 260976 67692 260982
rect 67640 260918 67692 260924
rect 67730 260944 67786 260953
rect 67730 260879 67732 260888
rect 67784 260879 67786 260888
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 259584 67694 259593
rect 67638 259519 67694 259528
rect 67652 259486 67680 259519
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 258632 67786 258641
rect 67730 258567 67786 258576
rect 67638 258224 67694 258233
rect 67638 258159 67640 258168
rect 67692 258159 67694 258168
rect 67640 258130 67692 258136
rect 67744 258126 67772 258567
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257961 67680 257994
rect 67638 257952 67694 257961
rect 67638 257887 67694 257896
rect 67638 256864 67694 256873
rect 67638 256799 67694 256808
rect 67652 256766 67680 256799
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 67730 255368 67786 255377
rect 67730 255303 67732 255312
rect 67784 255303 67786 255312
rect 67732 255274 67784 255280
rect 67640 255264 67692 255270
rect 67638 255232 67640 255241
rect 67692 255232 67694 255241
rect 67638 255167 67694 255176
rect 67730 254008 67786 254017
rect 67730 253943 67732 253952
rect 67784 253943 67786 253952
rect 67732 253914 67784 253920
rect 67640 253904 67692 253910
rect 67638 253872 67640 253881
rect 67692 253872 67694 253881
rect 67638 253807 67694 253816
rect 67638 252648 67694 252657
rect 67638 252583 67640 252592
rect 67692 252583 67694 252592
rect 67640 252554 67692 252560
rect 67730 249928 67786 249937
rect 67730 249863 67786 249872
rect 67744 249830 67772 249863
rect 67732 249824 67784 249830
rect 67638 249792 67694 249801
rect 67732 249766 67784 249772
rect 67638 249727 67640 249736
rect 67692 249727 67694 249736
rect 67640 249698 67692 249704
rect 67638 247752 67694 247761
rect 67638 247687 67694 247696
rect 67652 247178 67680 247687
rect 67730 247208 67786 247217
rect 67640 247172 67692 247178
rect 67730 247143 67786 247152
rect 67640 247114 67692 247120
rect 67744 247110 67772 247143
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67640 247036 67692 247042
rect 67640 246978 67692 246984
rect 67652 246673 67680 246978
rect 67638 246664 67694 246673
rect 67638 246599 67694 246608
rect 67640 245608 67692 245614
rect 67640 245550 67692 245556
rect 67652 245313 67680 245550
rect 67638 245304 67694 245313
rect 67638 245239 67694 245248
rect 67638 244624 67694 244633
rect 67638 244559 67694 244568
rect 67652 244322 67680 244559
rect 68296 244390 68324 286447
rect 68664 285433 68692 326470
rect 68940 326398 68968 349687
rect 69676 340082 69704 364306
rect 115216 354674 115244 458186
rect 115308 357406 115336 460090
rect 115492 459474 115520 460226
rect 115938 460184 115994 460193
rect 115938 460119 115994 460128
rect 115952 459785 115980 460119
rect 115938 459776 115994 459785
rect 115938 459711 115994 459720
rect 115480 459468 115532 459474
rect 115480 459410 115532 459416
rect 115388 391400 115440 391406
rect 115388 391342 115440 391348
rect 115400 385914 115428 391342
rect 115400 385886 115782 385914
rect 115296 357400 115348 357406
rect 115296 357342 115348 357348
rect 115216 354646 115336 354674
rect 115308 349217 115336 354646
rect 115952 353297 115980 459711
rect 116044 370297 116072 476070
rect 116136 384305 116164 487834
rect 116228 460290 116256 528566
rect 116320 492046 116348 584394
rect 116596 537538 116624 703054
rect 122748 683188 122800 683194
rect 122748 683130 122800 683136
rect 117504 586832 117556 586838
rect 117504 586774 117556 586780
rect 117320 578332 117372 578338
rect 117320 578274 117372 578280
rect 116584 537532 116636 537538
rect 116584 537474 116636 537480
rect 116308 492040 116360 492046
rect 116308 491982 116360 491988
rect 117332 488510 117360 578274
rect 117412 565956 117464 565962
rect 117412 565898 117464 565904
rect 117320 488504 117372 488510
rect 117320 488446 117372 488452
rect 117332 487898 117360 488446
rect 117320 487892 117372 487898
rect 117320 487834 117372 487840
rect 117318 484392 117374 484401
rect 117318 484327 117374 484336
rect 117228 466404 117280 466410
rect 117228 466346 117280 466352
rect 116216 460284 116268 460290
rect 116216 460226 116268 460232
rect 116122 384296 116178 384305
rect 116122 384231 116178 384240
rect 116674 384296 116730 384305
rect 116674 384231 116730 384240
rect 116688 383722 116716 384231
rect 116676 383716 116728 383722
rect 116676 383658 116728 383664
rect 116768 383648 116820 383654
rect 116122 383616 116178 383625
rect 116122 383551 116178 383560
rect 116766 383616 116768 383625
rect 116820 383616 116822 383625
rect 116766 383551 116822 383560
rect 116030 370288 116086 370297
rect 116030 370223 116086 370232
rect 116044 366994 116072 370223
rect 116032 366988 116084 366994
rect 116032 366930 116084 366936
rect 115938 353288 115994 353297
rect 115938 353223 115994 353232
rect 115294 349208 115350 349217
rect 115294 349143 115350 349152
rect 115296 342372 115348 342378
rect 115296 342314 115348 342320
rect 69676 340068 70058 340082
rect 69676 340054 70072 340068
rect 70044 338094 70072 340054
rect 70412 340054 70702 340082
rect 70032 338088 70084 338094
rect 70032 338030 70084 338036
rect 70412 335238 70440 340054
rect 71134 339960 71190 339969
rect 71134 339895 71190 339904
rect 70400 335232 70452 335238
rect 70400 335174 70452 335180
rect 70412 334014 70440 335174
rect 70400 334008 70452 334014
rect 70400 333950 70452 333956
rect 71044 334008 71096 334014
rect 71044 333950 71096 333956
rect 68928 326392 68980 326398
rect 68928 326334 68980 326340
rect 71056 305726 71084 333950
rect 71148 316742 71176 339895
rect 71332 338065 71360 340068
rect 71976 339522 72004 340068
rect 73264 339590 73292 340068
rect 73252 339584 73304 339590
rect 73252 339526 73304 339532
rect 71964 339516 72016 339522
rect 71964 339458 72016 339464
rect 71318 338056 71374 338065
rect 71318 337991 71374 338000
rect 71332 337521 71360 337991
rect 71318 337512 71374 337521
rect 71318 337447 71374 337456
rect 71976 336802 72004 339458
rect 72976 338088 73028 338094
rect 72976 338030 73028 338036
rect 71964 336796 72016 336802
rect 71964 336738 72016 336744
rect 72988 334665 73016 338030
rect 73264 335354 73292 339526
rect 73908 339386 73936 340068
rect 73896 339380 73948 339386
rect 73896 339322 73948 339328
rect 74448 339380 74500 339386
rect 74448 339322 74500 339328
rect 73172 335326 73292 335354
rect 72974 334656 73030 334665
rect 72974 334591 73030 334600
rect 72424 325032 72476 325038
rect 72424 324974 72476 324980
rect 71136 316736 71188 316742
rect 71136 316678 71188 316684
rect 71044 305720 71096 305726
rect 71044 305662 71096 305668
rect 71780 304292 71832 304298
rect 71780 304234 71832 304240
rect 71044 301504 71096 301510
rect 71044 301446 71096 301452
rect 70030 298208 70086 298217
rect 70030 298143 70086 298152
rect 69018 296848 69074 296857
rect 69018 296783 69074 296792
rect 68836 295452 68888 295458
rect 68836 295394 68888 295400
rect 68742 293992 68798 294001
rect 68742 293927 68798 293936
rect 68756 286113 68784 293927
rect 68848 290873 68876 295394
rect 68926 292768 68982 292777
rect 68926 292703 68982 292712
rect 68834 290864 68890 290873
rect 68834 290799 68890 290808
rect 68742 286104 68798 286113
rect 68742 286039 68798 286048
rect 68650 285424 68706 285433
rect 68650 285359 68706 285368
rect 68940 284073 68968 292703
rect 69032 289785 69060 296783
rect 70044 291924 70072 298143
rect 70676 294636 70728 294642
rect 70676 294578 70728 294584
rect 70688 291963 70716 294578
rect 71056 292369 71084 301446
rect 71792 294370 71820 304234
rect 71872 302252 71924 302258
rect 71872 302194 71924 302200
rect 71780 294364 71832 294370
rect 71780 294306 71832 294312
rect 71320 294296 71372 294302
rect 71320 294238 71372 294244
rect 71042 292360 71098 292369
rect 71042 292295 71098 292304
rect 71332 291963 71360 294238
rect 71884 291977 71912 302194
rect 72332 294364 72384 294370
rect 72332 294306 72384 294312
rect 72344 291977 72372 294306
rect 72436 294302 72464 324974
rect 73172 302841 73200 335326
rect 73344 324964 73396 324970
rect 73344 324906 73396 324912
rect 73158 302832 73214 302841
rect 73158 302767 73214 302776
rect 73252 298444 73304 298450
rect 73252 298386 73304 298392
rect 72424 294296 72476 294302
rect 72424 294238 72476 294244
rect 71884 291949 71990 291977
rect 72344 291949 72634 291977
rect 73264 291963 73292 298386
rect 73356 291977 73384 324906
rect 74460 309874 74488 339322
rect 74552 336734 74580 340068
rect 75840 339425 75868 340068
rect 75826 339416 75882 339425
rect 75826 339351 75882 339360
rect 75840 338094 75868 339351
rect 75828 338088 75880 338094
rect 75828 338030 75880 338036
rect 76484 337890 76512 340068
rect 77128 339454 77156 340068
rect 78432 339810 78460 340068
rect 78432 339782 78628 339810
rect 76656 339448 76708 339454
rect 76656 339390 76708 339396
rect 77116 339448 77168 339454
rect 77116 339390 77168 339396
rect 76472 337884 76524 337890
rect 76472 337826 76524 337832
rect 75184 336796 75236 336802
rect 75184 336738 75236 336744
rect 74540 336728 74592 336734
rect 74540 336670 74592 336676
rect 75196 318170 75224 336738
rect 75276 336728 75328 336734
rect 75276 336670 75328 336676
rect 75288 319462 75316 336670
rect 76484 335354 76512 337826
rect 76484 335326 76604 335354
rect 75276 319456 75328 319462
rect 75276 319398 75328 319404
rect 75184 318164 75236 318170
rect 75184 318106 75236 318112
rect 74448 309868 74500 309874
rect 74448 309810 74500 309816
rect 74632 307964 74684 307970
rect 74632 307906 74684 307912
rect 74644 306374 74672 307906
rect 74644 306346 75500 306374
rect 74540 300960 74592 300966
rect 74540 300902 74592 300908
rect 73356 291949 73922 291977
rect 74552 291963 74580 300902
rect 75184 298308 75236 298314
rect 75184 298250 75236 298256
rect 75196 291963 75224 298250
rect 75472 291938 75500 306346
rect 75920 303816 75972 303822
rect 75920 303758 75972 303764
rect 75932 291977 75960 303758
rect 76576 296041 76604 335326
rect 76668 315353 76696 339390
rect 77300 337408 77352 337414
rect 77300 337350 77352 337356
rect 78600 337362 78628 339782
rect 79060 339697 79088 340068
rect 79658 339810 79686 340068
rect 79336 339782 79686 339810
rect 79046 339688 79102 339697
rect 79046 339623 79102 339632
rect 79060 337385 79088 339623
rect 79046 337376 79102 337385
rect 76654 315344 76710 315353
rect 76654 315279 76710 315288
rect 77312 306374 77340 337350
rect 78600 337334 78720 337362
rect 78692 336666 78720 337334
rect 79046 337311 79102 337320
rect 78680 336660 78732 336666
rect 78680 336602 78732 336608
rect 78692 331809 78720 336602
rect 79336 336530 79364 339782
rect 80704 338836 80756 338842
rect 80704 338778 80756 338784
rect 79968 338088 80020 338094
rect 79968 338030 80020 338036
rect 79324 336524 79376 336530
rect 79324 336466 79376 336472
rect 78678 331800 78734 331809
rect 78678 331735 78734 331744
rect 78772 307828 78824 307834
rect 78772 307770 78824 307776
rect 78784 306374 78812 307770
rect 79336 307222 79364 336466
rect 79980 329118 80008 338030
rect 79968 329112 80020 329118
rect 79968 329054 80020 329060
rect 80060 312656 80112 312662
rect 80060 312598 80112 312604
rect 79324 307216 79376 307222
rect 79324 307158 79376 307164
rect 77312 306346 78076 306374
rect 78784 306346 79364 306374
rect 77760 297560 77812 297566
rect 77760 297502 77812 297508
rect 76562 296032 76618 296041
rect 76562 295967 76618 295976
rect 77116 292732 77168 292738
rect 77116 292674 77168 292680
rect 75932 291949 76498 291977
rect 77128 291963 77156 292674
rect 77772 291963 77800 297502
rect 78048 291938 78076 306346
rect 79048 294772 79100 294778
rect 79048 294714 79100 294720
rect 79060 291963 79088 294714
rect 79336 291938 79364 306346
rect 80072 291977 80100 312598
rect 80716 304366 80744 338778
rect 80992 337686 81020 340068
rect 80980 337680 81032 337686
rect 80980 337622 81032 337628
rect 81440 337680 81492 337686
rect 81440 337622 81492 337628
rect 81452 333946 81480 337622
rect 81636 336802 81664 340068
rect 82280 339250 82308 340068
rect 82268 339244 82320 339250
rect 82268 339186 82320 339192
rect 83568 338026 83596 340068
rect 83556 338020 83608 338026
rect 83556 337962 83608 337968
rect 81624 336796 81676 336802
rect 81624 336738 81676 336744
rect 81636 335306 81664 336738
rect 83568 335354 83596 337962
rect 84212 337958 84240 340068
rect 84810 339810 84838 340068
rect 84764 339782 84838 339810
rect 86160 339810 86188 340068
rect 86160 339782 86264 339810
rect 84200 337952 84252 337958
rect 84200 337894 84252 337900
rect 84764 336462 84792 339782
rect 84842 337512 84898 337521
rect 84842 337447 84898 337456
rect 84752 336456 84804 336462
rect 84752 336398 84804 336404
rect 83476 335326 83596 335354
rect 81624 335300 81676 335306
rect 81624 335242 81676 335248
rect 81440 333940 81492 333946
rect 81440 333882 81492 333888
rect 81452 332654 81480 333882
rect 81440 332648 81492 332654
rect 81440 332590 81492 332596
rect 82084 332648 82136 332654
rect 82084 332590 82136 332596
rect 82096 322153 82124 332590
rect 82082 322144 82138 322153
rect 82082 322079 82138 322088
rect 83476 309806 83504 335326
rect 84856 318102 84884 337447
rect 86236 333878 86264 339782
rect 86788 337822 86816 340068
rect 87432 339454 87460 340068
rect 88736 339810 88764 340068
rect 89318 339810 89346 340068
rect 88736 339782 89024 339810
rect 87420 339448 87472 339454
rect 87420 339390 87472 339396
rect 87604 339448 87656 339454
rect 87604 339390 87656 339396
rect 86776 337816 86828 337822
rect 86776 337758 86828 337764
rect 87616 335170 87644 339390
rect 88996 336598 89024 339782
rect 89088 339782 89346 339810
rect 90024 339810 90052 340068
rect 90024 339782 90404 339810
rect 88984 336592 89036 336598
rect 88984 336534 89036 336540
rect 87604 335164 87656 335170
rect 87604 335106 87656 335112
rect 86224 333872 86276 333878
rect 86224 333814 86276 333820
rect 84844 318096 84896 318102
rect 84844 318038 84896 318044
rect 83464 309800 83516 309806
rect 83464 309742 83516 309748
rect 81440 307896 81492 307902
rect 81440 307838 81492 307844
rect 80704 304360 80756 304366
rect 80704 304302 80756 304308
rect 80980 294092 81032 294098
rect 80980 294034 81032 294040
rect 80072 291949 80362 291977
rect 80992 291963 81020 294034
rect 81452 291977 81480 307838
rect 85580 303680 85632 303686
rect 85580 303622 85632 303628
rect 84200 301096 84252 301102
rect 84200 301038 84252 301044
rect 81900 299600 81952 299606
rect 81900 299542 81952 299548
rect 81452 291949 81650 291977
rect 81912 291938 81940 299542
rect 82912 298376 82964 298382
rect 82912 298318 82964 298324
rect 82924 291963 82952 298318
rect 83556 295588 83608 295594
rect 83556 295530 83608 295536
rect 83568 291963 83596 295530
rect 84212 291963 84240 301038
rect 84844 294772 84896 294778
rect 84844 294714 84896 294720
rect 84856 291963 84884 294714
rect 85488 294364 85540 294370
rect 85488 294306 85540 294312
rect 85500 291963 85528 294306
rect 85592 294302 85620 303622
rect 85672 302388 85724 302394
rect 85672 302330 85724 302336
rect 85580 294296 85632 294302
rect 85580 294238 85632 294244
rect 85684 291938 85712 302330
rect 86236 300286 86264 333814
rect 86316 323604 86368 323610
rect 86316 323546 86368 323552
rect 86224 300280 86276 300286
rect 86224 300222 86276 300228
rect 86328 294370 86356 323546
rect 88996 313954 89024 336534
rect 89088 333985 89116 339782
rect 89074 333976 89130 333985
rect 89074 333911 89130 333920
rect 88984 313948 89036 313954
rect 88984 313890 89036 313896
rect 89088 312594 89116 333911
rect 90376 332586 90404 339782
rect 91008 338156 91060 338162
rect 91008 338098 91060 338104
rect 90364 332580 90416 332586
rect 90364 332522 90416 332528
rect 89076 312588 89128 312594
rect 89076 312530 89128 312536
rect 88340 309188 88392 309194
rect 88340 309130 88392 309136
rect 88352 306374 88380 309130
rect 88352 306346 89116 306374
rect 87512 302456 87564 302462
rect 87512 302398 87564 302404
rect 87420 294840 87472 294846
rect 87420 294782 87472 294788
rect 86316 294364 86368 294370
rect 86316 294306 86368 294312
rect 86500 294296 86552 294302
rect 86500 294238 86552 294244
rect 86512 291977 86540 294238
rect 86512 291949 86802 291977
rect 87432 291963 87460 294782
rect 87524 291977 87552 302398
rect 88708 296948 88760 296954
rect 88708 296890 88760 296896
rect 87524 291949 88090 291977
rect 88720 291963 88748 296890
rect 89088 291977 89116 306346
rect 89720 305040 89772 305046
rect 89720 304982 89772 304988
rect 89732 291977 89760 304982
rect 90376 301578 90404 332522
rect 91020 324290 91048 338098
rect 91296 336734 91324 340068
rect 91940 338162 91968 340068
rect 91928 338156 91980 338162
rect 91928 338098 91980 338104
rect 92584 336870 92612 340068
rect 93228 339318 93256 340068
rect 93216 339312 93268 339318
rect 93216 339254 93268 339260
rect 92572 336864 92624 336870
rect 92572 336806 92624 336812
rect 91284 336728 91336 336734
rect 91284 336670 91336 336676
rect 92388 336728 92440 336734
rect 92388 336670 92440 336676
rect 91008 324284 91060 324290
rect 91008 324226 91060 324232
rect 91100 313336 91152 313342
rect 91100 313278 91152 313284
rect 91112 312662 91140 313278
rect 91100 312656 91152 312662
rect 91100 312598 91152 312604
rect 92400 307057 92428 336670
rect 93228 335354 93256 339254
rect 93136 335326 93256 335354
rect 92386 307048 92442 307057
rect 92386 306983 92442 306992
rect 90364 301572 90416 301578
rect 90364 301514 90416 301520
rect 93136 300354 93164 335326
rect 94516 332586 94544 340068
rect 95160 333946 95188 340068
rect 95804 337890 95832 340068
rect 95792 337884 95844 337890
rect 95792 337826 95844 337832
rect 95240 336864 95292 336870
rect 95240 336806 95292 336812
rect 95148 333940 95200 333946
rect 95148 333882 95200 333888
rect 95160 332654 95188 333882
rect 94596 332648 94648 332654
rect 94596 332590 94648 332596
rect 95148 332648 95200 332654
rect 95148 332590 95200 332596
rect 94504 332580 94556 332586
rect 94504 332522 94556 332528
rect 93952 320884 94004 320890
rect 93952 320826 94004 320832
rect 93216 316804 93268 316810
rect 93216 316746 93268 316752
rect 93124 300348 93176 300354
rect 93124 300290 93176 300296
rect 93228 300234 93256 316746
rect 92952 300206 93256 300234
rect 90638 298344 90694 298353
rect 90638 298279 90694 298288
rect 89088 291949 89378 291977
rect 89732 291949 90022 291977
rect 90652 291963 90680 298279
rect 91928 295724 91980 295730
rect 91928 295666 91980 295672
rect 91284 294704 91336 294710
rect 91284 294646 91336 294652
rect 91296 291963 91324 294646
rect 91940 291963 91968 295666
rect 92952 295390 92980 300206
rect 93216 296812 93268 296818
rect 93216 296754 93268 296760
rect 92572 295384 92624 295390
rect 92572 295326 92624 295332
rect 92940 295384 92992 295390
rect 92940 295326 92992 295332
rect 92584 291963 92612 295326
rect 93228 291963 93256 296754
rect 93964 294370 93992 320826
rect 94044 319524 94096 319530
rect 94044 319466 94096 319472
rect 93952 294364 94004 294370
rect 93952 294306 94004 294312
rect 93860 292800 93912 292806
rect 93860 292742 93912 292748
rect 93872 291963 93900 292742
rect 94056 291977 94084 319466
rect 94608 304201 94636 332590
rect 95252 330721 95280 336806
rect 96526 331120 96582 331129
rect 96526 331055 96582 331064
rect 96540 330721 96568 331055
rect 95238 330712 95294 330721
rect 95238 330647 95294 330656
rect 96526 330712 96582 330721
rect 96526 330647 96582 330656
rect 94594 304192 94650 304201
rect 94594 304127 94650 304136
rect 96540 300121 96568 330647
rect 97092 328438 97120 340068
rect 97264 338768 97316 338774
rect 97264 338710 97316 338716
rect 97080 328432 97132 328438
rect 97080 328374 97132 328380
rect 97276 312662 97304 338710
rect 97736 337958 97764 340068
rect 97724 337952 97776 337958
rect 97724 337894 97776 337900
rect 98380 337754 98408 340068
rect 98368 337748 98420 337754
rect 98368 337690 98420 337696
rect 99668 337414 99696 340068
rect 100312 339250 100340 340068
rect 100300 339244 100352 339250
rect 100300 339186 100352 339192
rect 99656 337408 99708 337414
rect 99656 337350 99708 337356
rect 100024 336796 100076 336802
rect 100024 336738 100076 336744
rect 98000 331968 98052 331974
rect 98000 331910 98052 331916
rect 97264 312656 97316 312662
rect 97264 312598 97316 312604
rect 96526 300112 96582 300121
rect 96526 300047 96582 300056
rect 94780 294364 94832 294370
rect 94780 294306 94832 294312
rect 94056 291949 94530 291977
rect 94792 291938 94820 294306
rect 95790 294128 95846 294137
rect 95790 294063 95846 294072
rect 95804 291963 95832 294063
rect 97080 293276 97132 293282
rect 97080 293218 97132 293224
rect 96436 292596 96488 292602
rect 96436 292538 96488 292544
rect 96448 291963 96476 292538
rect 97092 291963 97120 293218
rect 97724 292596 97776 292602
rect 97724 292538 97776 292544
rect 97736 291963 97764 292538
rect 98012 291977 98040 331910
rect 100036 305658 100064 336738
rect 100956 320142 100984 340068
rect 102244 339114 102272 340068
rect 102232 339108 102284 339114
rect 102232 339050 102284 339056
rect 102888 337278 102916 340068
rect 103336 339108 103388 339114
rect 103336 339050 103388 339056
rect 102876 337272 102928 337278
rect 102876 337214 102928 337220
rect 100944 320136 100996 320142
rect 100944 320078 100996 320084
rect 101404 318300 101456 318306
rect 101404 318242 101456 318248
rect 100024 305652 100076 305658
rect 100024 305594 100076 305600
rect 100944 296880 100996 296886
rect 100944 296822 100996 296828
rect 99656 295520 99708 295526
rect 99656 295462 99708 295468
rect 99010 292632 99066 292641
rect 99010 292567 99066 292576
rect 98012 291949 98394 291977
rect 99024 291963 99052 292567
rect 99668 291963 99696 295462
rect 100956 291963 100984 296822
rect 101416 294030 101444 318242
rect 103348 307086 103376 339050
rect 103428 337408 103480 337414
rect 103428 337350 103480 337356
rect 103336 307080 103388 307086
rect 103336 307022 103388 307028
rect 102140 299532 102192 299538
rect 102140 299474 102192 299480
rect 101404 294024 101456 294030
rect 101404 293966 101456 293972
rect 101588 294024 101640 294030
rect 101588 293966 101640 293972
rect 101600 291963 101628 293966
rect 102152 291977 102180 299474
rect 102876 298240 102928 298246
rect 102876 298182 102928 298188
rect 102152 291949 102258 291977
rect 102888 291963 102916 298182
rect 103440 298178 103468 337350
rect 103532 337074 103560 340068
rect 104164 338768 104216 338774
rect 104164 338710 104216 338716
rect 103520 337068 103572 337074
rect 103520 337010 103572 337016
rect 103428 298172 103480 298178
rect 103428 298114 103480 298120
rect 104176 294778 104204 338710
rect 104820 335238 104848 340068
rect 104900 337272 104952 337278
rect 104900 337214 104952 337220
rect 104808 335232 104860 335238
rect 104808 335174 104860 335180
rect 104820 334694 104848 335174
rect 104808 334688 104860 334694
rect 104808 334630 104860 334636
rect 104912 333878 104940 337214
rect 104900 333872 104952 333878
rect 104900 333814 104952 333820
rect 105464 331226 105492 340068
rect 105544 337748 105596 337754
rect 105544 337690 105596 337696
rect 105452 331220 105504 331226
rect 105452 331162 105504 331168
rect 105556 327826 105584 337690
rect 106108 327826 106136 340068
rect 107412 339810 107440 340068
rect 107412 339782 107608 339810
rect 107580 336734 107608 339782
rect 108040 338094 108068 340068
rect 108638 339810 108666 340068
rect 109926 339810 109954 340068
rect 108316 339782 108666 339810
rect 109880 339782 109954 339810
rect 108028 338088 108080 338094
rect 108028 338030 108080 338036
rect 108040 337754 108068 338030
rect 108028 337748 108080 337754
rect 108028 337690 108080 337696
rect 107568 336728 107620 336734
rect 107568 336670 107620 336676
rect 106280 331968 106332 331974
rect 106280 331910 106332 331916
rect 105544 327820 105596 327826
rect 105544 327762 105596 327768
rect 106096 327820 106148 327826
rect 106096 327762 106148 327768
rect 106188 326460 106240 326466
rect 106188 326402 106240 326408
rect 106200 298178 106228 326402
rect 106292 306374 106320 331910
rect 106292 306346 106872 306374
rect 104808 298172 104860 298178
rect 104808 298114 104860 298120
rect 106188 298172 106240 298178
rect 106188 298114 106240 298120
rect 104164 294772 104216 294778
rect 104164 294714 104216 294720
rect 104164 294024 104216 294030
rect 104164 293966 104216 293972
rect 103520 292664 103572 292670
rect 103520 292606 103572 292612
rect 103532 291963 103560 292606
rect 104176 291963 104204 293966
rect 104820 291963 104848 298114
rect 106200 296714 106228 298114
rect 106108 296686 106228 296714
rect 105452 294296 105504 294302
rect 105452 294238 105504 294244
rect 105464 291963 105492 294238
rect 106108 291963 106136 296686
rect 106740 294432 106792 294438
rect 106740 294374 106792 294380
rect 106752 291963 106780 294374
rect 106844 291977 106872 306346
rect 106924 301028 106976 301034
rect 106924 300970 106976 300976
rect 106936 294846 106964 300970
rect 107580 296177 107608 336670
rect 108316 335306 108344 339782
rect 109132 337068 109184 337074
rect 109132 337010 109184 337016
rect 109144 336054 109172 337010
rect 109880 336598 109908 339782
rect 109868 336592 109920 336598
rect 109868 336534 109920 336540
rect 109132 336048 109184 336054
rect 109132 335990 109184 335996
rect 108304 335300 108356 335306
rect 108304 335242 108356 335248
rect 107660 333328 107712 333334
rect 107660 333270 107712 333276
rect 107672 306374 107700 333270
rect 108316 325038 108344 335242
rect 109880 334626 109908 336534
rect 109868 334620 109920 334626
rect 109868 334562 109920 334568
rect 110616 329798 110644 340068
rect 111062 330440 111118 330449
rect 111062 330375 111118 330384
rect 110604 329792 110656 329798
rect 110604 329734 110656 329740
rect 108304 325032 108356 325038
rect 108304 324974 108356 324980
rect 107672 306346 108436 306374
rect 107566 296168 107622 296177
rect 107566 296103 107622 296112
rect 106924 294840 106976 294846
rect 106924 294782 106976 294788
rect 108028 294364 108080 294370
rect 108028 294306 108080 294312
rect 106844 291949 107410 291977
rect 108040 291963 108068 294306
rect 108408 291977 108436 306346
rect 109684 304292 109736 304298
rect 109684 304234 109736 304240
rect 109696 291977 109724 304234
rect 110972 300892 111024 300898
rect 110972 300834 111024 300840
rect 110604 296744 110656 296750
rect 110604 296686 110656 296692
rect 110420 294024 110472 294030
rect 110420 293966 110472 293972
rect 110432 293282 110460 293966
rect 110420 293276 110472 293282
rect 110420 293218 110472 293224
rect 108408 291949 108698 291977
rect 109696 291949 109986 291977
rect 110616 291963 110644 296686
rect 110984 291977 111012 300834
rect 111076 297401 111104 330375
rect 111260 320074 111288 340068
rect 112444 336796 112496 336802
rect 112444 336738 112496 336744
rect 111248 320068 111300 320074
rect 111248 320010 111300 320016
rect 112456 319530 112484 336738
rect 112548 335170 112576 340068
rect 113192 339318 113220 340068
rect 113836 339590 113864 340068
rect 115124 339658 115152 340068
rect 113916 339652 113968 339658
rect 113916 339594 113968 339600
rect 115112 339652 115164 339658
rect 115112 339594 115164 339600
rect 113824 339584 113876 339590
rect 113824 339526 113876 339532
rect 113180 339312 113232 339318
rect 113180 339254 113232 339260
rect 113836 336802 113864 339526
rect 113824 336796 113876 336802
rect 113824 336738 113876 336744
rect 113928 336682 113956 339594
rect 114008 339312 114060 339318
rect 114008 339254 114060 339260
rect 113836 336654 113956 336682
rect 112536 335164 112588 335170
rect 112536 335106 112588 335112
rect 113088 335164 113140 335170
rect 113088 335106 113140 335112
rect 112444 319524 112496 319530
rect 112444 319466 112496 319472
rect 113100 308446 113128 335106
rect 113836 316810 113864 336654
rect 114020 335354 114048 339254
rect 113928 335326 114048 335354
rect 113928 323610 113956 335326
rect 115204 333260 115256 333266
rect 115204 333202 115256 333208
rect 114468 327820 114520 327826
rect 114468 327762 114520 327768
rect 113916 323604 113968 323610
rect 113916 323546 113968 323552
rect 113824 316804 113876 316810
rect 113824 316746 113876 316752
rect 113088 308440 113140 308446
rect 113088 308382 113140 308388
rect 112444 302320 112496 302326
rect 112444 302262 112496 302268
rect 111062 297392 111118 297401
rect 111062 297327 111118 297336
rect 111892 295384 111944 295390
rect 111892 295326 111944 295332
rect 110984 291949 111274 291977
rect 111904 291963 111932 295326
rect 112456 294438 112484 302262
rect 114480 300801 114508 327762
rect 114560 319456 114612 319462
rect 114560 319398 114612 319404
rect 113178 300792 113234 300801
rect 113178 300727 113234 300736
rect 114466 300792 114522 300801
rect 114466 300727 114522 300736
rect 112444 294432 112496 294438
rect 112444 294374 112496 294380
rect 112536 294160 112588 294166
rect 112536 294102 112588 294108
rect 112548 291963 112576 294102
rect 113192 291963 113220 300727
rect 114480 299577 114508 300727
rect 114466 299568 114522 299577
rect 114466 299503 114522 299512
rect 113824 294228 113876 294234
rect 113824 294170 113876 294176
rect 113836 291963 113864 294170
rect 114572 291977 114600 319398
rect 115216 293350 115244 333202
rect 115308 318238 115336 342314
rect 115386 339552 115442 339561
rect 115386 339487 115442 339496
rect 115400 326534 115428 339487
rect 115768 338026 115796 340068
rect 115756 338020 115808 338026
rect 115756 337962 115808 337968
rect 115388 326528 115440 326534
rect 115388 326470 115440 326476
rect 116044 324970 116072 366930
rect 116136 326466 116164 383551
rect 117240 360330 117268 466346
rect 117332 385490 117360 484327
rect 117424 476066 117452 565898
rect 117516 532166 117544 586774
rect 118700 585404 118752 585410
rect 118700 585346 118752 585352
rect 117504 532160 117556 532166
rect 117504 532102 117556 532108
rect 117504 500268 117556 500274
rect 117504 500210 117556 500216
rect 117412 476060 117464 476066
rect 117412 476002 117464 476008
rect 117516 461553 117544 500210
rect 117596 497616 117648 497622
rect 117596 497558 117648 497564
rect 117502 461544 117558 461553
rect 117502 461479 117558 461488
rect 117502 459640 117558 459649
rect 117502 459575 117558 459584
rect 117412 443692 117464 443698
rect 117412 443634 117464 443640
rect 117320 385484 117372 385490
rect 117320 385426 117372 385432
rect 117318 385384 117374 385393
rect 117318 385319 117374 385328
rect 117332 384826 117360 385319
rect 117424 384946 117452 443634
rect 117516 384985 117544 459575
rect 117608 440910 117636 497558
rect 118712 489802 118740 585346
rect 121460 585200 121512 585206
rect 121460 585142 121512 585148
rect 118792 583908 118844 583914
rect 118792 583850 118844 583856
rect 118804 496806 118832 583850
rect 118976 582616 119028 582622
rect 118976 582558 119028 582564
rect 118884 497684 118936 497690
rect 118884 497626 118936 497632
rect 118792 496800 118844 496806
rect 118792 496742 118844 496748
rect 118792 494896 118844 494902
rect 118792 494838 118844 494844
rect 118804 494766 118832 494838
rect 118792 494760 118844 494766
rect 118792 494702 118844 494708
rect 118792 491428 118844 491434
rect 118792 491370 118844 491376
rect 118804 489938 118832 491370
rect 118792 489932 118844 489938
rect 118792 489874 118844 489880
rect 118700 489796 118752 489802
rect 118700 489738 118752 489744
rect 118792 482316 118844 482322
rect 118792 482258 118844 482264
rect 118700 480956 118752 480962
rect 118700 480898 118752 480904
rect 117780 476060 117832 476066
rect 117780 476002 117832 476008
rect 117792 475386 117820 476002
rect 117780 475380 117832 475386
rect 117780 475322 117832 475328
rect 117596 440904 117648 440910
rect 117596 440846 117648 440852
rect 117596 402416 117648 402422
rect 117596 402358 117648 402364
rect 117502 384976 117558 384985
rect 117412 384940 117464 384946
rect 117502 384911 117558 384920
rect 117412 384882 117464 384888
rect 117332 384798 117544 384826
rect 117412 384600 117464 384606
rect 117412 384542 117464 384548
rect 117318 382256 117374 382265
rect 117318 382191 117320 382200
rect 117372 382191 117374 382200
rect 117320 382162 117372 382168
rect 117318 380896 117374 380905
rect 117318 380831 117320 380840
rect 117372 380831 117374 380840
rect 117320 380802 117372 380808
rect 116676 360324 116728 360330
rect 116676 360266 116728 360272
rect 117228 360324 117280 360330
rect 117228 360266 117280 360272
rect 116688 359825 116716 360266
rect 116674 359816 116730 359825
rect 116674 359751 116730 359760
rect 117320 357400 117372 357406
rect 117320 357342 117372 357348
rect 116584 351348 116636 351354
rect 116584 351290 116636 351296
rect 116124 326460 116176 326466
rect 116124 326402 116176 326408
rect 116032 324964 116084 324970
rect 116032 324906 116084 324912
rect 115296 318232 115348 318238
rect 115296 318174 115348 318180
rect 115940 311160 115992 311166
rect 115940 311102 115992 311108
rect 115294 305688 115350 305697
rect 115294 305623 115350 305632
rect 115308 294273 115336 305623
rect 115846 295352 115902 295361
rect 115846 295287 115902 295296
rect 115860 294642 115888 295287
rect 115848 294636 115900 294642
rect 115848 294578 115900 294584
rect 115294 294264 115350 294273
rect 115294 294199 115350 294208
rect 115754 294264 115810 294273
rect 115754 294199 115810 294208
rect 115204 293344 115256 293350
rect 115204 293286 115256 293292
rect 114282 291952 114338 291961
rect 75472 291910 75842 291938
rect 78048 291910 78418 291938
rect 79336 291910 79706 291938
rect 81912 291910 82282 291938
rect 85684 291910 86146 291938
rect 94792 291910 95162 291938
rect 109592 291916 109644 291922
rect 109342 291864 109592 291870
rect 114572 291949 115138 291977
rect 115768 291963 115796 294199
rect 115952 291977 115980 311102
rect 116596 300218 116624 351290
rect 117332 350985 117360 357342
rect 117424 351665 117452 384542
rect 117516 373425 117544 384798
rect 117502 373416 117558 373425
rect 117502 373351 117504 373360
rect 117556 373351 117558 373360
rect 117504 373322 117556 373328
rect 117516 373291 117544 373322
rect 117608 363633 117636 402358
rect 117688 385484 117740 385490
rect 117688 385426 117740 385432
rect 117700 380186 117728 385426
rect 118238 384976 118294 384985
rect 118238 384911 118240 384920
rect 118292 384911 118294 384920
rect 118240 384882 118292 384888
rect 117688 380180 117740 380186
rect 117688 380122 117740 380128
rect 117700 379545 117728 380122
rect 117686 379536 117742 379545
rect 117686 379471 117742 379480
rect 118606 378856 118662 378865
rect 118606 378791 118608 378800
rect 118660 378791 118662 378800
rect 118608 378762 118660 378768
rect 118608 377460 118660 377466
rect 118608 377402 118660 377408
rect 118620 376825 118648 377402
rect 118606 376816 118662 376825
rect 118606 376751 118662 376760
rect 118606 376136 118662 376145
rect 118712 376122 118740 480898
rect 118804 378185 118832 482258
rect 118896 447846 118924 497626
rect 118988 494766 119016 582558
rect 120172 579692 120224 579698
rect 120172 579634 120224 579640
rect 120080 568608 120132 568614
rect 120080 568550 120132 568556
rect 119068 496800 119120 496806
rect 119068 496742 119120 496748
rect 118976 494760 119028 494766
rect 118976 494702 119028 494708
rect 119080 491434 119108 496742
rect 119986 495000 120042 495009
rect 119986 494935 120042 494944
rect 119068 491428 119120 491434
rect 119068 491370 119120 491376
rect 120000 467838 120028 494935
rect 120092 476066 120120 568550
rect 120184 488481 120212 579634
rect 120264 560380 120316 560386
rect 120264 560322 120316 560328
rect 120170 488472 120226 488481
rect 120170 488407 120226 488416
rect 120172 481636 120224 481642
rect 120172 481578 120224 481584
rect 120080 476060 120132 476066
rect 120080 476002 120132 476008
rect 119988 467832 120040 467838
rect 119988 467774 120040 467780
rect 119344 465724 119396 465730
rect 119344 465666 119396 465672
rect 118884 447840 118936 447846
rect 118884 447782 118936 447788
rect 118884 398268 118936 398274
rect 118884 398210 118936 398216
rect 118790 378176 118846 378185
rect 118790 378111 118846 378120
rect 118662 376094 118740 376122
rect 118606 376071 118608 376080
rect 118660 376071 118662 376080
rect 118608 376042 118660 376048
rect 118516 376032 118568 376038
rect 118516 375974 118568 375980
rect 118528 375465 118556 375974
rect 118514 375456 118570 375465
rect 118514 375391 118570 375400
rect 118608 375352 118660 375358
rect 118608 375294 118660 375300
rect 118620 374105 118648 375294
rect 118606 374096 118662 374105
rect 118606 374031 118662 374040
rect 118422 372736 118478 372745
rect 118422 372671 118478 372680
rect 118436 372638 118464 372671
rect 118424 372632 118476 372638
rect 118424 372574 118476 372580
rect 118606 371376 118662 371385
rect 118606 371311 118662 371320
rect 118620 371278 118648 371311
rect 118608 371272 118660 371278
rect 118608 371214 118660 371220
rect 118514 367976 118570 367985
rect 118514 367911 118570 367920
rect 118528 367130 118556 367911
rect 118606 367296 118662 367305
rect 118606 367231 118608 367240
rect 118660 367231 118662 367240
rect 118608 367202 118660 367208
rect 118516 367124 118568 367130
rect 118516 367066 118568 367072
rect 118608 367056 118660 367062
rect 118608 366998 118660 367004
rect 118620 365945 118648 366998
rect 118606 365936 118662 365945
rect 118606 365871 118662 365880
rect 118606 365256 118662 365265
rect 118606 365191 118662 365200
rect 118620 364818 118648 365191
rect 118700 365152 118752 365158
rect 118700 365094 118752 365100
rect 118608 364812 118660 364818
rect 118608 364754 118660 364760
rect 118606 364576 118662 364585
rect 118712 364562 118740 365094
rect 118662 364534 118740 364562
rect 118606 364511 118662 364520
rect 117594 363624 117650 363633
rect 117594 363559 117650 363568
rect 117964 362908 118016 362914
rect 117964 362850 118016 362856
rect 117976 362545 118004 362850
rect 117962 362536 118018 362545
rect 117962 362471 118018 362480
rect 118608 362228 118660 362234
rect 118608 362170 118660 362176
rect 118620 361865 118648 362170
rect 118606 361856 118662 361865
rect 118606 361791 118662 361800
rect 118606 361176 118662 361185
rect 118606 361111 118662 361120
rect 118620 360262 118648 361111
rect 118608 360256 118660 360262
rect 118608 360198 118660 360204
rect 118148 360188 118200 360194
rect 118148 360130 118200 360136
rect 118160 359145 118188 360130
rect 118146 359136 118202 359145
rect 118146 359071 118202 359080
rect 118608 358488 118660 358494
rect 118606 358456 118608 358465
rect 118660 358456 118662 358465
rect 118606 358391 118662 358400
rect 117686 357096 117742 357105
rect 117686 357031 117688 357040
rect 117740 357031 117742 357040
rect 117688 357002 117740 357008
rect 118608 356040 118660 356046
rect 118608 355982 118660 355988
rect 118620 355745 118648 355982
rect 118606 355736 118662 355745
rect 118606 355671 118662 355680
rect 118608 354680 118660 354686
rect 118608 354622 118660 354628
rect 118054 354376 118110 354385
rect 118054 354311 118110 354320
rect 118068 353326 118096 354311
rect 118620 353705 118648 354622
rect 118606 353696 118662 353705
rect 118606 353631 118662 353640
rect 118056 353320 118108 353326
rect 118056 353262 118108 353268
rect 117962 353016 118018 353025
rect 117962 352951 118018 352960
rect 117410 351656 117466 351665
rect 117410 351591 117466 351600
rect 117318 350976 117374 350985
rect 117318 350911 117374 350920
rect 117778 348936 117834 348945
rect 117778 348871 117834 348880
rect 117792 347818 117820 348871
rect 117780 347812 117832 347818
rect 117780 347754 117832 347760
rect 117412 347744 117464 347750
rect 117412 347686 117464 347692
rect 117424 347585 117452 347686
rect 117410 347576 117466 347585
rect 117410 347511 117466 347520
rect 116676 345092 116728 345098
rect 116676 345034 116728 345040
rect 116688 336666 116716 345034
rect 117780 340808 117832 340814
rect 117780 340750 117832 340756
rect 117792 340105 117820 340750
rect 117778 340096 117834 340105
rect 117778 340031 117834 340040
rect 116676 336660 116728 336666
rect 116676 336602 116728 336608
rect 116584 300212 116636 300218
rect 116584 300154 116636 300160
rect 117228 297424 117280 297430
rect 117228 297366 117280 297372
rect 117136 294364 117188 294370
rect 117136 294306 117188 294312
rect 117148 291990 117176 294306
rect 117240 294030 117268 297366
rect 117976 297022 118004 352951
rect 118514 351656 118570 351665
rect 118514 351591 118570 351600
rect 118424 351280 118476 351286
rect 118424 351222 118476 351228
rect 118436 350985 118464 351222
rect 118528 351218 118556 351591
rect 118516 351212 118568 351218
rect 118516 351154 118568 351160
rect 118422 350976 118478 350985
rect 118422 350911 118478 350920
rect 118606 350296 118662 350305
rect 118606 350231 118662 350240
rect 118620 349926 118648 350231
rect 118608 349920 118660 349926
rect 118608 349862 118660 349868
rect 118606 348256 118662 348265
rect 118606 348191 118662 348200
rect 118620 347886 118648 348191
rect 118608 347880 118660 347886
rect 118608 347822 118660 347828
rect 118608 346384 118660 346390
rect 118608 346326 118660 346332
rect 118330 346216 118386 346225
rect 118330 346151 118386 346160
rect 118344 345710 118372 346151
rect 118332 345704 118384 345710
rect 118332 345646 118384 345652
rect 118620 345545 118648 346326
rect 118606 345536 118662 345545
rect 118606 345471 118662 345480
rect 118608 345024 118660 345030
rect 118608 344966 118660 344972
rect 118620 344865 118648 344966
rect 118606 344856 118662 344865
rect 118606 344791 118662 344800
rect 118608 343596 118660 343602
rect 118608 343538 118660 343544
rect 118146 343496 118202 343505
rect 118146 343431 118202 343440
rect 118160 342310 118188 343431
rect 118620 342825 118648 343538
rect 118606 342816 118662 342825
rect 118606 342751 118662 342760
rect 118148 342304 118200 342310
rect 118148 342246 118200 342252
rect 118606 342136 118662 342145
rect 118606 342071 118662 342080
rect 118620 341562 118648 342071
rect 118608 341556 118660 341562
rect 118608 341498 118660 341504
rect 118056 340876 118108 340882
rect 118056 340818 118108 340824
rect 118068 340785 118096 340818
rect 118054 340776 118110 340785
rect 118054 340711 118110 340720
rect 118056 320544 118108 320550
rect 118056 320486 118108 320492
rect 117964 297016 118016 297022
rect 117964 296958 118016 296964
rect 118068 295798 118096 320486
rect 118056 295792 118108 295798
rect 118056 295734 118108 295740
rect 117688 295656 117740 295662
rect 117688 295598 117740 295604
rect 117228 294024 117280 294030
rect 117228 293966 117280 293972
rect 117136 291984 117188 291990
rect 115952 291949 116426 291977
rect 114338 291910 114482 291938
rect 117700 291963 117728 295598
rect 118068 291977 118096 295734
rect 118620 292913 118648 341498
rect 118712 331974 118740 364534
rect 118804 342378 118832 378111
rect 118896 370025 118924 398210
rect 119356 390726 119384 465666
rect 120080 450628 120132 450634
rect 120080 450570 120132 450576
rect 119344 390720 119396 390726
rect 119344 390662 119396 390668
rect 119356 389842 119384 390662
rect 119344 389836 119396 389842
rect 119344 389778 119396 389784
rect 119344 388136 119396 388142
rect 119344 388078 119396 388084
rect 119356 377369 119384 388078
rect 119342 377360 119398 377369
rect 119342 377295 119398 377304
rect 119988 371952 120040 371958
rect 119988 371894 120040 371900
rect 118882 370016 118938 370025
rect 118882 369951 118938 369960
rect 118974 368656 119030 368665
rect 118974 368591 119030 368600
rect 118988 368558 119016 368591
rect 118976 368552 119028 368558
rect 118976 368494 119028 368500
rect 119344 367804 119396 367810
rect 119344 367746 119396 367752
rect 119356 367266 119384 367746
rect 119344 367260 119396 367266
rect 119344 367202 119396 367208
rect 118792 342372 118844 342378
rect 118792 342314 118844 342320
rect 118792 340944 118844 340950
rect 118792 340886 118844 340892
rect 118700 331968 118752 331974
rect 118700 331910 118752 331916
rect 118804 314022 118832 340886
rect 118792 314016 118844 314022
rect 118792 313958 118844 313964
rect 119356 304298 119384 367202
rect 120000 356153 120028 371894
rect 119986 356144 120042 356153
rect 119986 356079 120042 356088
rect 120092 340950 120120 450570
rect 120184 376038 120212 481578
rect 120276 469198 120304 560322
rect 121472 494154 121500 585142
rect 121552 581052 121604 581058
rect 121552 580994 121604 581000
rect 121564 534818 121592 580994
rect 121644 578944 121696 578950
rect 121644 578886 121696 578892
rect 121656 538966 121684 578886
rect 121920 574048 121972 574054
rect 121920 573990 121972 573996
rect 121932 573374 121960 573990
rect 122760 573374 122788 683130
rect 129004 643136 129056 643142
rect 129004 643078 129056 643084
rect 123116 586764 123168 586770
rect 123116 586706 123168 586712
rect 122840 585336 122892 585342
rect 122840 585278 122892 585284
rect 121920 573368 121972 573374
rect 121920 573310 121972 573316
rect 122748 573368 122800 573374
rect 122748 573310 122800 573316
rect 121644 538960 121696 538966
rect 121644 538902 121696 538908
rect 122104 538892 122156 538898
rect 122104 538834 122156 538840
rect 121736 537736 121788 537742
rect 121736 537678 121788 537684
rect 121552 534812 121604 534818
rect 121552 534754 121604 534760
rect 121644 532024 121696 532030
rect 121644 531966 121696 531972
rect 121460 494148 121512 494154
rect 121460 494090 121512 494096
rect 120356 494080 120408 494086
rect 120356 494022 120408 494028
rect 120264 469192 120316 469198
rect 120264 469134 120316 469140
rect 120276 468586 120304 469134
rect 120264 468580 120316 468586
rect 120264 468522 120316 468528
rect 120368 442513 120396 494022
rect 120354 442504 120410 442513
rect 120354 442439 120410 442448
rect 120356 391332 120408 391338
rect 120356 391274 120408 391280
rect 120262 381032 120318 381041
rect 120262 380967 120318 380976
rect 120172 376032 120224 376038
rect 120172 375974 120224 375980
rect 120172 360256 120224 360262
rect 120172 360198 120224 360204
rect 120184 360126 120212 360198
rect 120172 360120 120224 360126
rect 120172 360062 120224 360068
rect 120080 340944 120132 340950
rect 120080 340886 120132 340892
rect 120276 320550 120304 380967
rect 120368 345014 120396 391274
rect 121472 391270 121500 494090
rect 121656 469878 121684 531966
rect 121644 469872 121696 469878
rect 121644 469814 121696 469820
rect 121642 463584 121698 463593
rect 121642 463519 121698 463528
rect 121550 439376 121606 439385
rect 121550 439311 121606 439320
rect 121564 439006 121592 439311
rect 121552 439000 121604 439006
rect 121552 438942 121604 438948
rect 121656 395350 121684 463519
rect 121748 438734 121776 537678
rect 122116 439385 122144 538834
rect 122852 489870 122880 585278
rect 123024 581120 123076 581126
rect 123024 581062 123076 581068
rect 122932 539028 122984 539034
rect 122932 538970 122984 538976
rect 122840 489864 122892 489870
rect 122840 489806 122892 489812
rect 122102 439376 122158 439385
rect 121920 439340 121972 439346
rect 122944 439346 122972 538970
rect 123036 488442 123064 581062
rect 123128 496194 123156 586706
rect 127072 586696 127124 586702
rect 127072 586638 127124 586644
rect 124312 586628 124364 586634
rect 124312 586570 124364 586576
rect 124220 583772 124272 583778
rect 124220 583714 124272 583720
rect 124232 497554 124260 583714
rect 124220 497548 124272 497554
rect 124220 497490 124272 497496
rect 123116 496188 123168 496194
rect 123116 496130 123168 496136
rect 124220 496188 124272 496194
rect 124220 496130 124272 496136
rect 123208 494828 123260 494834
rect 123208 494770 123260 494776
rect 123116 491224 123168 491230
rect 123116 491166 123168 491172
rect 123128 489977 123156 491166
rect 123114 489968 123170 489977
rect 123114 489903 123170 489912
rect 123024 488436 123076 488442
rect 123024 488378 123076 488384
rect 123024 467832 123076 467838
rect 123024 467774 123076 467780
rect 122102 439311 122158 439320
rect 122932 439340 122984 439346
rect 121920 439282 121972 439288
rect 122932 439282 122984 439288
rect 121932 438870 121960 439282
rect 121920 438864 121972 438870
rect 121920 438806 121972 438812
rect 122196 438864 122248 438870
rect 122196 438806 122248 438812
rect 121736 438728 121788 438734
rect 121736 438670 121788 438676
rect 122104 398200 122156 398206
rect 122104 398142 122156 398148
rect 121644 395344 121696 395350
rect 121644 395286 121696 395292
rect 121460 391264 121512 391270
rect 121460 391206 121512 391212
rect 120632 389156 120684 389162
rect 120632 389098 120684 389104
rect 120644 388074 120672 389098
rect 121918 388920 121974 388929
rect 121918 388855 121974 388864
rect 120632 388068 120684 388074
rect 120632 388010 120684 388016
rect 120644 387841 120672 388010
rect 121932 388006 121960 388855
rect 121920 388000 121972 388006
rect 121920 387942 121972 387948
rect 122116 387841 122144 398142
rect 120630 387832 120686 387841
rect 120630 387767 120686 387776
rect 122102 387832 122158 387841
rect 122102 387767 122158 387776
rect 122102 385248 122158 385257
rect 122102 385183 122158 385192
rect 121460 384940 121512 384946
rect 121460 384882 121512 384888
rect 121472 382974 121500 384882
rect 121460 382968 121512 382974
rect 121460 382910 121512 382916
rect 121460 377460 121512 377466
rect 121460 377402 121512 377408
rect 120724 360120 120776 360126
rect 120724 360062 120776 360068
rect 120368 344986 120488 345014
rect 120460 337822 120488 344986
rect 120736 338774 120764 360062
rect 120724 338768 120776 338774
rect 120724 338710 120776 338716
rect 120448 337816 120500 337822
rect 120448 337758 120500 337764
rect 120460 337521 120488 337758
rect 120446 337512 120502 337521
rect 120446 337447 120502 337456
rect 120264 320544 120316 320550
rect 120264 320486 120316 320492
rect 120724 315308 120776 315314
rect 120724 315250 120776 315256
rect 119712 309868 119764 309874
rect 119712 309810 119764 309816
rect 119724 306374 119752 309810
rect 120080 307216 120132 307222
rect 120080 307158 120132 307164
rect 119724 306346 119844 306374
rect 119344 304292 119396 304298
rect 119344 304234 119396 304240
rect 119620 294024 119672 294030
rect 119620 293966 119672 293972
rect 119344 293956 119396 293962
rect 119344 293898 119396 293904
rect 118606 292904 118662 292913
rect 118606 292839 118662 292848
rect 119356 291977 119384 293898
rect 118068 291949 118358 291977
rect 119002 291949 119384 291977
rect 117136 291926 117188 291932
rect 119632 291924 119660 293966
rect 117320 291916 117372 291922
rect 114282 291887 114338 291896
rect 109342 291858 109644 291864
rect 117070 291864 117320 291870
rect 117070 291858 117372 291864
rect 109342 291842 109632 291858
rect 117070 291842 117360 291858
rect 119816 289921 119844 306346
rect 119802 289912 119858 289921
rect 119802 289847 119858 289856
rect 69018 289776 69074 289785
rect 69018 289711 69074 289720
rect 68926 284064 68982 284073
rect 68926 283999 68982 284008
rect 68374 280528 68430 280537
rect 68374 280463 68430 280472
rect 68388 245002 68416 280463
rect 69110 268288 69166 268297
rect 69110 268223 69166 268232
rect 68834 251832 68890 251841
rect 68834 251767 68890 251776
rect 68848 248946 68876 251767
rect 68836 248940 68888 248946
rect 68836 248882 68888 248888
rect 69018 245712 69074 245721
rect 69018 245647 69074 245656
rect 68376 244996 68428 245002
rect 68376 244938 68428 244944
rect 68284 244384 68336 244390
rect 68284 244326 68336 244332
rect 67640 244316 67692 244322
rect 67640 244258 67692 244264
rect 67732 244248 67784 244254
rect 67732 244190 67784 244196
rect 67822 244216 67878 244225
rect 67744 243953 67772 244190
rect 67822 244151 67878 244160
rect 67730 243944 67786 243953
rect 67730 243879 67786 243888
rect 67836 242962 67864 244151
rect 67824 242956 67876 242962
rect 67824 242898 67876 242904
rect 67640 242888 67692 242894
rect 67640 242830 67692 242836
rect 67652 242593 67680 242830
rect 67638 242584 67694 242593
rect 67638 242519 67694 242528
rect 67638 241904 67694 241913
rect 67638 241839 67694 241848
rect 67652 241534 67680 241839
rect 67640 241528 67692 241534
rect 67640 241470 67692 241476
rect 67638 240544 67694 240553
rect 67638 240479 67694 240488
rect 67652 240174 67680 240479
rect 67640 240168 67692 240174
rect 67640 240110 67692 240116
rect 67548 196784 67600 196790
rect 67548 196726 67600 196732
rect 69032 184210 69060 245647
rect 69124 206378 69152 268223
rect 120092 256465 120120 307158
rect 120170 292904 120226 292913
rect 120170 292839 120226 292848
rect 120078 256456 120134 256465
rect 120078 256391 120134 256400
rect 69294 255912 69350 255921
rect 69294 255847 69350 255856
rect 69308 236774 69336 255847
rect 120078 251016 120134 251025
rect 120078 250951 120134 250960
rect 119986 240952 120042 240961
rect 119986 240887 120042 240896
rect 119896 240168 119948 240174
rect 69676 240094 70058 240122
rect 119646 240116 119896 240122
rect 119646 240110 119948 240116
rect 119646 240094 119936 240110
rect 69296 236768 69348 236774
rect 69296 236710 69348 236716
rect 69676 219434 69704 240094
rect 70400 239828 70452 239834
rect 70400 239770 70452 239776
rect 69216 219406 69704 219434
rect 69112 206372 69164 206378
rect 69112 206314 69164 206320
rect 69020 184204 69072 184210
rect 69020 184146 69072 184152
rect 69216 180130 69244 219406
rect 70412 191146 70440 239770
rect 70688 238754 70716 240037
rect 71320 239834 71348 240037
rect 71964 239850 71992 240037
rect 71308 239828 71360 239834
rect 71308 239770 71360 239776
rect 71884 239822 71992 239850
rect 70504 238726 70716 238754
rect 70504 195294 70532 238726
rect 71884 224262 71912 239822
rect 72620 238542 72648 240037
rect 73252 239850 73280 240037
rect 73896 239850 73924 240037
rect 73172 239822 73280 239850
rect 73816 239822 73924 239850
rect 72608 238536 72660 238542
rect 72608 238478 72660 238484
rect 71872 224256 71924 224262
rect 71872 224198 71924 224204
rect 73172 198014 73200 239822
rect 73816 219434 73844 239822
rect 74552 238754 74580 240037
rect 74552 238726 74672 238754
rect 74540 233980 74592 233986
rect 74540 233922 74592 233928
rect 73264 219406 73844 219434
rect 73264 215966 73292 219406
rect 73252 215960 73304 215966
rect 73252 215902 73304 215908
rect 73160 198008 73212 198014
rect 74552 197985 74580 233922
rect 74644 217394 74672 238726
rect 75196 233986 75224 240037
rect 75840 238649 75868 240037
rect 75920 239828 75972 239834
rect 75920 239770 75972 239776
rect 75826 238640 75882 238649
rect 75826 238575 75882 238584
rect 75184 233980 75236 233986
rect 75184 233922 75236 233928
rect 75932 228313 75960 239770
rect 76484 238754 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 77772 238754 77800 240037
rect 78404 239816 78432 240037
rect 76024 238726 76512 238754
rect 77312 238726 77800 238754
rect 78324 239788 78432 239816
rect 78680 239828 78732 239834
rect 76024 230450 76052 238726
rect 76012 230444 76064 230450
rect 76012 230386 76064 230392
rect 75918 228304 75974 228313
rect 75918 228239 75974 228248
rect 74632 217388 74684 217394
rect 74632 217330 74684 217336
rect 73160 197950 73212 197956
rect 74538 197976 74594 197985
rect 74538 197911 74594 197920
rect 70492 195288 70544 195294
rect 70492 195230 70544 195236
rect 70400 191140 70452 191146
rect 70400 191082 70452 191088
rect 77312 189689 77340 238726
rect 78324 219434 78352 239788
rect 78680 239770 78732 239776
rect 77404 219406 78352 219434
rect 77404 211818 77432 219406
rect 77392 211812 77444 211818
rect 77392 211754 77444 211760
rect 78692 192545 78720 239770
rect 79060 238754 79088 240037
rect 79692 239834 79720 240037
rect 79680 239828 79732 239834
rect 79680 239770 79732 239776
rect 80348 238754 80376 240037
rect 80980 239816 81008 240037
rect 78784 238726 79088 238754
rect 80072 238726 80376 238754
rect 80900 239788 81008 239816
rect 78784 227050 78812 238726
rect 78772 227044 78824 227050
rect 78772 226986 78824 226992
rect 78678 192536 78734 192545
rect 78678 192471 78734 192480
rect 77298 189680 77354 189689
rect 77298 189615 77354 189624
rect 80072 182850 80100 238726
rect 80900 219434 80928 239788
rect 81636 234530 81664 240037
rect 82280 238882 82308 240037
rect 82912 239816 82940 240037
rect 83556 239816 83584 240037
rect 82832 239788 82940 239816
rect 83476 239788 83584 239816
rect 82268 238876 82320 238882
rect 82268 238818 82320 238824
rect 81624 234524 81676 234530
rect 81624 234466 81676 234472
rect 82832 226302 82860 239788
rect 83476 233238 83504 239788
rect 84212 239442 84240 240037
rect 84212 239414 84424 239442
rect 84292 239352 84344 239358
rect 84292 239294 84344 239300
rect 83464 233232 83516 233238
rect 83464 233174 83516 233180
rect 82820 226296 82872 226302
rect 82820 226238 82872 226244
rect 80164 219406 80928 219434
rect 80164 184278 80192 219406
rect 83476 203590 83504 233174
rect 84108 231872 84160 231878
rect 84160 231826 84240 231854
rect 84108 231814 84160 231820
rect 83464 203584 83516 203590
rect 83464 203526 83516 203532
rect 84212 185638 84240 231826
rect 84304 195430 84332 239294
rect 84396 226953 84424 239414
rect 84856 231878 84884 240037
rect 85500 239358 85528 240037
rect 85488 239352 85540 239358
rect 85488 239294 85540 239300
rect 86144 238754 86172 240037
rect 86144 238726 86264 238754
rect 86236 238513 86264 238726
rect 86222 238504 86278 238513
rect 86222 238439 86278 238448
rect 84844 231872 84896 231878
rect 84844 231814 84896 231820
rect 84382 226944 84438 226953
rect 84382 226879 84438 226888
rect 86236 196654 86264 238439
rect 86788 237250 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86776 237244 86828 237250
rect 86776 237186 86828 237192
rect 86224 196648 86276 196654
rect 86224 196590 86276 196596
rect 84292 195424 84344 195430
rect 84292 195366 84344 195372
rect 84200 185632 84252 185638
rect 84200 185574 84252 185580
rect 80152 184272 80204 184278
rect 80152 184214 80204 184220
rect 80060 182844 80112 182850
rect 80060 182786 80112 182792
rect 86972 181626 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 88720 238754 88748 240037
rect 87064 238726 87460 238754
rect 88352 238726 88748 238754
rect 87064 209001 87092 238726
rect 88352 216034 88380 238726
rect 89364 238474 89392 240037
rect 89720 239828 89772 239834
rect 89720 239770 89772 239776
rect 89352 238468 89404 238474
rect 89352 238410 89404 238416
rect 88340 216028 88392 216034
rect 88340 215970 88392 215976
rect 87050 208992 87106 209001
rect 87050 208927 87106 208936
rect 89732 188426 89760 239770
rect 90008 238754 90036 240037
rect 90640 239834 90668 240037
rect 90628 239828 90680 239834
rect 90628 239770 90680 239776
rect 89824 238726 90036 238754
rect 89824 209098 89852 238726
rect 91296 235890 91324 240037
rect 91940 238678 91968 240037
rect 91928 238672 91980 238678
rect 91928 238614 91980 238620
rect 91940 238513 91968 238614
rect 91926 238504 91982 238513
rect 91926 238439 91982 238448
rect 91284 235884 91336 235890
rect 91284 235826 91336 235832
rect 92584 232558 92612 240037
rect 93216 239816 93244 240037
rect 93136 239788 93244 239816
rect 92572 232552 92624 232558
rect 92572 232494 92624 232500
rect 93136 219434 93164 239788
rect 92492 219406 93164 219434
rect 89812 209092 89864 209098
rect 89812 209034 89864 209040
rect 92492 196722 92520 219406
rect 93872 199578 93900 240037
rect 93952 239828 94004 239834
rect 93952 239770 94004 239776
rect 93964 203658 93992 239770
rect 94516 238754 94544 240037
rect 95148 239834 95176 240037
rect 95136 239828 95188 239834
rect 95136 239770 95188 239776
rect 94056 238726 94544 238754
rect 94056 231130 94084 238726
rect 95804 238610 95832 240037
rect 95792 238604 95844 238610
rect 95792 238546 95844 238552
rect 96448 238066 96476 240037
rect 97092 238754 97120 240037
rect 97724 239816 97752 240037
rect 96632 238726 97120 238754
rect 97644 239788 97752 239816
rect 96436 238060 96488 238066
rect 96436 238002 96488 238008
rect 94044 231124 94096 231130
rect 94044 231066 94096 231072
rect 93952 203652 94004 203658
rect 93952 203594 94004 203600
rect 96632 199714 96660 238726
rect 97644 229770 97672 239788
rect 98380 238746 98408 240037
rect 98368 238740 98420 238746
rect 98368 238682 98420 238688
rect 99024 238542 99052 240037
rect 99380 239828 99432 239834
rect 99380 239770 99432 239776
rect 99012 238536 99064 238542
rect 99012 238478 99064 238484
rect 97632 229764 97684 229770
rect 97632 229706 97684 229712
rect 96620 199708 96672 199714
rect 96620 199650 96672 199656
rect 93860 199572 93912 199578
rect 93860 199514 93912 199520
rect 92480 196716 92532 196722
rect 92480 196658 92532 196664
rect 89720 188420 89772 188426
rect 89720 188362 89772 188368
rect 99392 188358 99420 239770
rect 99668 238754 99696 240037
rect 100300 239834 100328 240037
rect 100944 239884 100972 240037
rect 100864 239856 100972 239884
rect 100288 239828 100340 239834
rect 100288 239770 100340 239776
rect 100760 239828 100812 239834
rect 100760 239770 100812 239776
rect 99484 238726 99696 238754
rect 99484 213217 99512 238726
rect 99470 213208 99526 213217
rect 99470 213143 99526 213152
rect 100772 202230 100800 239770
rect 100864 206446 100892 239856
rect 101588 239834 101616 240037
rect 102232 239884 102260 240037
rect 102152 239856 102260 239884
rect 101576 239828 101628 239834
rect 101576 239770 101628 239776
rect 100852 206440 100904 206446
rect 100852 206382 100904 206388
rect 102152 206310 102180 239856
rect 102888 237454 102916 240037
rect 103532 238882 103560 240037
rect 103520 238876 103572 238882
rect 103520 238818 103572 238824
rect 103518 238776 103574 238785
rect 104176 238754 104204 240037
rect 104820 238785 104848 240037
rect 104900 239828 104952 239834
rect 104900 239770 104952 239776
rect 103518 238711 103574 238720
rect 103624 238726 104204 238754
rect 104806 238776 104862 238785
rect 102876 237448 102928 237454
rect 102876 237390 102928 237396
rect 102140 206304 102192 206310
rect 102140 206246 102192 206252
rect 100760 202224 100812 202230
rect 100760 202166 100812 202172
rect 103532 191350 103560 238711
rect 103624 220114 103652 238726
rect 104806 238711 104862 238720
rect 103612 220108 103664 220114
rect 103612 220050 103664 220056
rect 104912 207738 104940 239770
rect 105464 238134 105492 240037
rect 106096 239834 106124 240037
rect 106084 239828 106136 239834
rect 106084 239770 106136 239776
rect 106752 238814 106780 240037
rect 106740 238808 106792 238814
rect 106740 238750 106792 238756
rect 105452 238128 105504 238134
rect 105452 238070 105504 238076
rect 105544 237448 105596 237454
rect 105544 237390 105596 237396
rect 104900 207732 104952 207738
rect 104900 207674 104952 207680
rect 105556 205018 105584 237390
rect 107396 237386 107424 240037
rect 107660 239828 107712 239834
rect 107660 239770 107712 239776
rect 107384 237380 107436 237386
rect 107384 237322 107436 237328
rect 105544 205012 105596 205018
rect 105544 204954 105596 204960
rect 107672 195362 107700 239770
rect 108040 238754 108068 240037
rect 108672 239834 108700 240037
rect 108660 239828 108712 239834
rect 108660 239770 108712 239776
rect 107764 238726 108068 238754
rect 107764 199510 107792 238726
rect 109040 234592 109092 234598
rect 109040 234534 109092 234540
rect 109052 234190 109080 234534
rect 109972 234190 110000 240037
rect 110616 237386 110644 240037
rect 111260 238754 111288 240037
rect 111892 239850 111920 240037
rect 110984 238726 111288 238754
rect 111812 239822 111920 239850
rect 110604 237380 110656 237386
rect 110604 237322 110656 237328
rect 110616 236842 110644 237322
rect 110604 236836 110656 236842
rect 110604 236778 110656 236784
rect 109040 234184 109092 234190
rect 109040 234126 109092 234132
rect 109960 234184 110012 234190
rect 109960 234126 110012 234132
rect 107752 199504 107804 199510
rect 107752 199446 107804 199452
rect 107660 195356 107712 195362
rect 107660 195298 107712 195304
rect 103520 191344 103572 191350
rect 103520 191286 103572 191292
rect 105544 189100 105596 189106
rect 105544 189042 105596 189048
rect 99380 188352 99432 188358
rect 99380 188294 99432 188300
rect 101956 187808 102008 187814
rect 101956 187750 102008 187756
rect 99288 186380 99340 186386
rect 99288 186322 99340 186328
rect 97724 182232 97776 182238
rect 97724 182174 97776 182180
rect 86960 181620 87012 181626
rect 86960 181562 87012 181568
rect 69204 180124 69256 180130
rect 69204 180066 69256 180072
rect 67454 180024 67510 180033
rect 67454 179959 67510 179968
rect 97736 177721 97764 182174
rect 99300 177721 99328 186322
rect 100668 183592 100720 183598
rect 100668 183534 100720 183540
rect 97722 177712 97778 177721
rect 97722 177647 97778 177656
rect 99286 177712 99342 177721
rect 99286 177647 99342 177656
rect 100680 176769 100708 183534
rect 101968 177721 101996 187750
rect 104808 187740 104860 187746
rect 104808 187682 104860 187688
rect 102048 177880 102100 177886
rect 102048 177822 102100 177828
rect 101954 177712 102010 177721
rect 101954 177647 102010 177656
rect 102060 176769 102088 177822
rect 104820 177721 104848 187682
rect 105556 177886 105584 189042
rect 109052 185842 109080 234126
rect 110984 219434 111012 238726
rect 111064 236836 111116 236842
rect 111064 236778 111116 236784
rect 110432 219406 111012 219434
rect 110432 194070 110460 219406
rect 110420 194064 110472 194070
rect 110420 194006 110472 194012
rect 109040 185836 109092 185842
rect 109040 185778 109092 185784
rect 110142 179480 110198 179489
rect 110142 179415 110198 179424
rect 105544 177880 105596 177886
rect 105544 177822 105596 177828
rect 104806 177712 104862 177721
rect 104806 177647 104862 177656
rect 110156 177041 110184 179415
rect 110142 177032 110198 177041
rect 107016 176996 107068 177002
rect 110142 176967 110198 176976
rect 107016 176938 107068 176944
rect 105728 176928 105780 176934
rect 105728 176870 105780 176876
rect 103336 176860 103388 176866
rect 103336 176802 103388 176808
rect 103348 176769 103376 176802
rect 105740 176769 105768 176870
rect 107028 176769 107056 176938
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 102046 176760 102102 176769
rect 102046 176695 102102 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 105726 176760 105782 176769
rect 105726 176695 105782 176704
rect 107014 176760 107070 176769
rect 107014 176695 107070 176704
rect 108118 176760 108174 176769
rect 108118 176695 108120 176704
rect 108172 176695 108174 176704
rect 108120 176666 108172 176672
rect 110696 176180 110748 176186
rect 110696 176122 110748 176128
rect 110708 175409 110736 176122
rect 111076 175982 111104 236778
rect 111812 191282 111840 239822
rect 112548 235958 112576 240037
rect 112536 235952 112588 235958
rect 112536 235894 112588 235900
rect 113192 203590 113220 240037
rect 113836 238610 113864 240037
rect 113824 238604 113876 238610
rect 113824 238546 113876 238552
rect 114480 235958 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 235952 114520 235958
rect 114468 235894 114520 235900
rect 113180 203584 113232 203590
rect 113180 203526 113232 203532
rect 111800 191276 111852 191282
rect 111800 191218 111852 191224
rect 114572 191214 114600 239770
rect 115124 238882 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 115112 238876 115164 238882
rect 115112 238818 115164 238824
rect 116412 238754 116440 240037
rect 115952 238726 116440 238754
rect 114560 191208 114612 191214
rect 114560 191150 114612 191156
rect 114468 184952 114520 184958
rect 114468 184894 114520 184900
rect 114100 180872 114152 180878
rect 114100 180814 114152 180820
rect 114112 177721 114140 180814
rect 114480 177721 114508 184894
rect 115952 184346 115980 238726
rect 117056 237318 117084 240037
rect 117044 237312 117096 237318
rect 117044 237254 117096 237260
rect 117700 237182 117728 240037
rect 118344 238746 118372 240037
rect 118988 239970 119016 240037
rect 120000 239970 120028 240887
rect 118976 239964 119028 239970
rect 118976 239906 119028 239912
rect 119988 239964 120040 239970
rect 119988 239906 120040 239912
rect 118332 238740 118384 238746
rect 118332 238682 118384 238688
rect 117688 237176 117740 237182
rect 117688 237118 117740 237124
rect 117700 235278 117728 237118
rect 117688 235272 117740 235278
rect 117688 235214 117740 235220
rect 120092 202842 120120 250951
rect 120184 244905 120212 292839
rect 120736 257145 120764 315250
rect 121472 266778 121500 377402
rect 122116 367713 122144 385183
rect 122102 367704 122158 367713
rect 122102 367639 122158 367648
rect 121552 365084 121604 365090
rect 121552 365026 121604 365032
rect 121564 364818 121592 365026
rect 121552 364812 121604 364818
rect 121552 364754 121604 364760
rect 121564 286770 121592 364754
rect 122104 362228 122156 362234
rect 122104 362170 122156 362176
rect 121644 357060 121696 357066
rect 121644 357002 121696 357008
rect 121656 354006 121684 357002
rect 121644 354000 121696 354006
rect 121644 353942 121696 353948
rect 121642 314256 121698 314265
rect 121642 314191 121698 314200
rect 121656 313342 121684 314191
rect 121644 313336 121696 313342
rect 121644 313278 121696 313284
rect 121644 292528 121696 292534
rect 121644 292470 121696 292476
rect 121656 291825 121684 292470
rect 121642 291816 121698 291825
rect 121642 291751 121698 291760
rect 121642 290456 121698 290465
rect 121642 290391 121698 290400
rect 121656 289882 121684 290391
rect 121644 289876 121696 289882
rect 121644 289818 121696 289824
rect 121734 289096 121790 289105
rect 121734 289031 121790 289040
rect 121748 288454 121776 289031
rect 121736 288448 121788 288454
rect 121736 288390 121788 288396
rect 121826 288416 121882 288425
rect 121644 288380 121696 288386
rect 121826 288351 121882 288360
rect 121644 288322 121696 288328
rect 121656 287745 121684 288322
rect 121642 287736 121698 287745
rect 121642 287671 121698 287680
rect 121840 287094 121868 288351
rect 121828 287088 121880 287094
rect 121642 287056 121698 287065
rect 121828 287030 121880 287036
rect 121642 286991 121698 287000
rect 121656 286890 121684 286991
rect 121736 286952 121788 286958
rect 121736 286894 121788 286900
rect 121644 286884 121696 286890
rect 121644 286826 121696 286832
rect 121564 286742 121684 286770
rect 121552 286680 121604 286686
rect 121552 286622 121604 286628
rect 121564 286385 121592 286622
rect 121550 286376 121606 286385
rect 121550 286311 121606 286320
rect 121656 285138 121684 286742
rect 121748 285705 121776 286894
rect 121734 285696 121790 285705
rect 121734 285631 121790 285640
rect 121564 285110 121684 285138
rect 121564 284753 121592 285110
rect 121642 285016 121698 285025
rect 121642 284951 121698 284960
rect 121550 284744 121606 284753
rect 121550 284679 121606 284688
rect 121656 284374 121684 284951
rect 121644 284368 121696 284374
rect 121644 284310 121696 284316
rect 121552 284300 121604 284306
rect 121552 284242 121604 284248
rect 121564 283665 121592 284242
rect 121550 283656 121606 283665
rect 121550 283591 121606 283600
rect 121550 282976 121606 282985
rect 121550 282911 121552 282920
rect 121604 282911 121606 282920
rect 121552 282882 121604 282888
rect 121642 282296 121698 282305
rect 121642 282231 121698 282240
rect 121656 281654 121684 282231
rect 121644 281648 121696 281654
rect 121550 281616 121606 281625
rect 121644 281590 121696 281596
rect 121550 281551 121552 281560
rect 121604 281551 121606 281560
rect 121552 281522 121604 281528
rect 121550 280936 121606 280945
rect 121550 280871 121606 280880
rect 121564 280226 121592 280871
rect 121552 280220 121604 280226
rect 121552 280162 121604 280168
rect 121642 279576 121698 279585
rect 121642 279511 121698 279520
rect 121550 278896 121606 278905
rect 121550 278831 121552 278840
rect 121604 278831 121606 278840
rect 121552 278802 121604 278808
rect 121656 278798 121684 279511
rect 121644 278792 121696 278798
rect 121644 278734 121696 278740
rect 121642 278216 121698 278225
rect 121642 278151 121698 278160
rect 121550 277536 121606 277545
rect 121550 277471 121552 277480
rect 121604 277471 121606 277480
rect 121552 277442 121604 277448
rect 121656 277438 121684 278151
rect 121644 277432 121696 277438
rect 121644 277374 121696 277380
rect 121550 276856 121606 276865
rect 121550 276791 121606 276800
rect 121564 276690 121592 276791
rect 121552 276684 121604 276690
rect 121552 276626 121604 276632
rect 121734 276176 121790 276185
rect 121734 276111 121790 276120
rect 121550 274816 121606 274825
rect 121550 274751 121606 274760
rect 121564 274718 121592 274751
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121644 274644 121696 274650
rect 121644 274586 121696 274592
rect 121656 274145 121684 274586
rect 121642 274136 121698 274145
rect 121642 274071 121698 274080
rect 121748 273970 121776 276111
rect 121826 275496 121882 275505
rect 121826 275431 121882 275440
rect 121736 273964 121788 273970
rect 121736 273906 121788 273912
rect 121550 273456 121606 273465
rect 121550 273391 121606 273400
rect 121564 273290 121592 273391
rect 121552 273284 121604 273290
rect 121552 273226 121604 273232
rect 121644 273216 121696 273222
rect 121644 273158 121696 273164
rect 121656 272785 121684 273158
rect 121642 272776 121698 272785
rect 121642 272711 121698 272720
rect 121550 272096 121606 272105
rect 121550 272031 121606 272040
rect 121564 271930 121592 272031
rect 121552 271924 121604 271930
rect 121552 271866 121604 271872
rect 121550 271416 121606 271425
rect 121550 271351 121606 271360
rect 121564 270570 121592 271351
rect 121552 270564 121604 270570
rect 121552 270506 121604 270512
rect 121550 270056 121606 270065
rect 121550 269991 121606 270000
rect 121564 269210 121592 269991
rect 121840 269822 121868 275431
rect 121828 269816 121880 269822
rect 121828 269758 121880 269764
rect 121642 269376 121698 269385
rect 121642 269311 121698 269320
rect 121552 269204 121604 269210
rect 121552 269146 121604 269152
rect 121656 269142 121684 269311
rect 121644 269136 121696 269142
rect 121644 269078 121696 269084
rect 121552 269068 121604 269074
rect 121552 269010 121604 269016
rect 121564 268705 121592 269010
rect 121550 268696 121606 268705
rect 121550 268631 121606 268640
rect 121550 268016 121606 268025
rect 121550 267951 121606 267960
rect 121564 267782 121592 267951
rect 121552 267776 121604 267782
rect 121552 267718 121604 267724
rect 121734 267336 121790 267345
rect 121734 267271 121790 267280
rect 121472 266750 121684 266778
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266490 121500 266591
rect 121460 266484 121512 266490
rect 121460 266426 121512 266432
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121460 264920 121512 264926
rect 121460 264862 121512 264868
rect 121472 264625 121500 264862
rect 121458 264616 121514 264625
rect 121458 264551 121514 264560
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121552 262200 121604 262206
rect 121552 262142 121604 262148
rect 121564 261225 121592 262142
rect 121550 261216 121606 261225
rect 121550 261151 121606 261160
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121460 259344 121512 259350
rect 121460 259286 121512 259292
rect 121472 258505 121500 259286
rect 121550 259176 121606 259185
rect 121550 259111 121606 259120
rect 121458 258496 121514 258505
rect 121458 258431 121514 258440
rect 121564 258126 121592 259111
rect 121552 258120 121604 258126
rect 121552 258062 121604 258068
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 120722 257136 120778 257145
rect 120722 257071 120778 257080
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121460 256692 121512 256698
rect 121460 256634 121512 256640
rect 121472 255785 121500 256634
rect 121458 255776 121514 255785
rect 121458 255711 121514 255720
rect 121550 255096 121606 255105
rect 121550 255031 121606 255040
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 253978 121500 254351
rect 121564 254250 121592 255031
rect 121552 254244 121604 254250
rect 121552 254186 121604 254192
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121564 251870 121592 253671
rect 121656 252385 121684 266750
rect 121748 266422 121776 267271
rect 121736 266416 121788 266422
rect 121736 266358 121788 266364
rect 121734 261896 121790 261905
rect 121734 261831 121790 261840
rect 121748 260914 121776 261831
rect 121736 260908 121788 260914
rect 121736 260850 121788 260856
rect 121642 252376 121698 252385
rect 121642 252311 121698 252320
rect 121552 251864 121604 251870
rect 121552 251806 121604 251812
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121460 249756 121512 249762
rect 121460 249698 121512 249704
rect 121472 249665 121500 249698
rect 121458 249656 121514 249665
rect 121458 249591 121514 249600
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121550 245576 121606 245585
rect 121550 245511 121606 245520
rect 120170 244896 120226 244905
rect 120170 244831 120226 244840
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121550 244216 121606 244225
rect 121472 243545 121500 244190
rect 121550 244151 121606 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121564 242962 121592 244151
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121458 242791 121514 242800
rect 121552 242820 121604 242826
rect 121552 242762 121604 242768
rect 121564 242185 121592 242762
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 122116 241602 122144 362170
rect 122208 356794 122236 438806
rect 122840 389292 122892 389298
rect 122840 389234 122892 389240
rect 122288 388544 122340 388550
rect 122288 388486 122340 388492
rect 122300 376009 122328 388486
rect 122286 376000 122342 376009
rect 122286 375935 122342 375944
rect 122196 356788 122248 356794
rect 122196 356730 122248 356736
rect 122746 247616 122802 247625
rect 122852 247602 122880 389234
rect 123036 388929 123064 467774
rect 123116 396772 123168 396778
rect 123116 396714 123168 396720
rect 123022 388920 123078 388929
rect 123022 388855 123078 388864
rect 122932 385756 122984 385762
rect 122932 385698 122984 385704
rect 122944 371958 122972 385698
rect 122932 371952 122984 371958
rect 122932 371894 122984 371900
rect 122932 366988 122984 366994
rect 122932 366930 122984 366936
rect 122944 365022 122972 366930
rect 122932 365016 122984 365022
rect 122932 364958 122984 364964
rect 122932 345704 122984 345710
rect 122932 345646 122984 345652
rect 122944 251025 122972 345646
rect 123128 337414 123156 396714
rect 123220 392834 123248 494770
rect 123208 392828 123260 392834
rect 123208 392770 123260 392776
rect 124232 392601 124260 496130
rect 124324 494018 124352 586570
rect 125600 585268 125652 585274
rect 125600 585210 125652 585216
rect 124496 583024 124548 583030
rect 124496 582966 124548 582972
rect 124404 545760 124456 545766
rect 124404 545702 124456 545708
rect 124312 494012 124364 494018
rect 124312 493954 124364 493960
rect 124312 489932 124364 489938
rect 124312 489874 124364 489880
rect 124324 422278 124352 489874
rect 124416 454034 124444 545702
rect 124508 491230 124536 582966
rect 125612 491298 125640 585210
rect 126244 575612 126296 575618
rect 126244 575554 126296 575560
rect 125876 565888 125928 565894
rect 125876 565830 125928 565836
rect 125784 534744 125836 534750
rect 125784 534686 125836 534692
rect 125600 491292 125652 491298
rect 125600 491234 125652 491240
rect 124496 491224 124548 491230
rect 124496 491166 124548 491172
rect 125508 491224 125560 491230
rect 125508 491166 125560 491172
rect 125520 490618 125548 491166
rect 125508 490612 125560 490618
rect 125508 490554 125560 490560
rect 125612 490346 125640 491234
rect 125600 490340 125652 490346
rect 125600 490282 125652 490288
rect 125692 487892 125744 487898
rect 125692 487834 125744 487840
rect 125600 483676 125652 483682
rect 125600 483618 125652 483624
rect 124404 454028 124456 454034
rect 124404 453970 124456 453976
rect 124312 422272 124364 422278
rect 124312 422214 124364 422220
rect 124312 402280 124364 402286
rect 124312 402222 124364 402228
rect 124218 392592 124274 392601
rect 124218 392527 124274 392536
rect 124220 390720 124272 390726
rect 124220 390662 124272 390668
rect 124128 390040 124180 390046
rect 124128 389982 124180 389988
rect 124140 389298 124168 389982
rect 124128 389292 124180 389298
rect 124128 389234 124180 389240
rect 123852 373380 123904 373386
rect 123852 373322 123904 373328
rect 123864 369073 123892 373322
rect 123850 369064 123906 369073
rect 123850 368999 123906 369008
rect 124232 358494 124260 390662
rect 124220 358488 124272 358494
rect 124220 358430 124272 358436
rect 123116 337408 123168 337414
rect 123116 337350 123168 337356
rect 123116 300144 123168 300150
rect 123116 300086 123168 300092
rect 123024 297016 123076 297022
rect 123024 296958 123076 296964
rect 122930 251016 122986 251025
rect 122930 250951 122986 250960
rect 122802 247574 122880 247602
rect 122746 247551 122802 247560
rect 122104 241596 122156 241602
rect 122104 241538 122156 241544
rect 121460 241528 121512 241534
rect 122116 241505 122144 241538
rect 121460 241470 121512 241476
rect 122102 241496 122158 241505
rect 121472 240825 121500 241470
rect 122102 241431 122158 241440
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 122378 240136 122434 240145
rect 122378 240071 122434 240080
rect 122392 233986 122420 240071
rect 123036 238746 123064 296958
rect 123128 286686 123156 300086
rect 123116 286680 123168 286686
rect 123116 286622 123168 286628
rect 123484 254244 123536 254250
rect 123484 254186 123536 254192
rect 123024 238740 123076 238746
rect 123024 238682 123076 238688
rect 122380 233980 122432 233986
rect 122380 233922 122432 233928
rect 123496 211886 123524 254186
rect 124232 238542 124260 358430
rect 124324 345098 124352 402222
rect 124956 388476 125008 388482
rect 124956 388418 125008 388424
rect 124864 378208 124916 378214
rect 124864 378150 124916 378156
rect 124404 349920 124456 349926
rect 124404 349862 124456 349868
rect 124312 345092 124364 345098
rect 124312 345034 124364 345040
rect 124310 324320 124366 324329
rect 124310 324255 124312 324264
rect 124364 324255 124366 324264
rect 124312 324226 124364 324232
rect 124312 300280 124364 300286
rect 124312 300222 124364 300228
rect 124220 238536 124272 238542
rect 124220 238478 124272 238484
rect 124324 235958 124352 300222
rect 124416 297498 124444 349862
rect 124876 339386 124904 378150
rect 124968 356726 124996 388418
rect 125612 378842 125640 483618
rect 125704 383654 125732 487834
rect 125796 437442 125824 534686
rect 125888 474706 125916 565830
rect 126256 563718 126284 575554
rect 126244 563712 126296 563718
rect 126244 563654 126296 563660
rect 126256 483682 126284 563654
rect 127084 496126 127112 586638
rect 128360 571396 128412 571402
rect 128360 571338 128412 571344
rect 127256 553444 127308 553450
rect 127256 553386 127308 553392
rect 127164 537804 127216 537810
rect 127164 537746 127216 537752
rect 127072 496120 127124 496126
rect 127072 496062 127124 496068
rect 127072 490340 127124 490346
rect 127072 490282 127124 490288
rect 126244 483676 126296 483682
rect 126244 483618 126296 483624
rect 125876 474700 125928 474706
rect 125876 474642 125928 474648
rect 126980 460284 127032 460290
rect 126980 460226 127032 460232
rect 125784 437436 125836 437442
rect 125784 437378 125836 437384
rect 125876 392760 125928 392766
rect 125876 392702 125928 392708
rect 125784 387184 125836 387190
rect 125784 387126 125836 387132
rect 125692 383648 125744 383654
rect 125692 383590 125744 383596
rect 125612 378826 125732 378842
rect 125612 378820 125744 378826
rect 125612 378814 125692 378820
rect 125692 378762 125744 378768
rect 124956 356720 125008 356726
rect 124956 356662 125008 356668
rect 124864 339380 124916 339386
rect 124864 339322 124916 339328
rect 125600 339244 125652 339250
rect 125600 339186 125652 339192
rect 124404 297492 124456 297498
rect 124404 297434 124456 297440
rect 125508 294296 125560 294302
rect 125508 294238 125560 294244
rect 125520 293962 125548 294238
rect 125508 293956 125560 293962
rect 125508 293898 125560 293904
rect 125520 292890 125548 293898
rect 125428 292862 125548 292890
rect 125232 292732 125284 292738
rect 125232 292674 125284 292680
rect 125244 290442 125272 292674
rect 125428 292346 125456 292862
rect 125508 292732 125560 292738
rect 125508 292674 125560 292680
rect 125520 292466 125548 292674
rect 125508 292460 125560 292466
rect 125508 292402 125560 292408
rect 125428 292318 125548 292346
rect 125244 290414 125456 290442
rect 125428 259418 125456 290414
rect 125416 259412 125468 259418
rect 125416 259354 125468 259360
rect 125520 254590 125548 292318
rect 125612 263566 125640 339186
rect 125704 320890 125732 378762
rect 125796 337890 125824 387126
rect 125888 339250 125916 392702
rect 126244 380180 126296 380186
rect 126244 380122 126296 380128
rect 126256 349858 126284 380122
rect 126992 349926 127020 460226
rect 127084 389162 127112 490282
rect 127176 442882 127204 537746
rect 127268 460193 127296 553386
rect 128372 480214 128400 571338
rect 128636 559564 128688 559570
rect 128636 559506 128688 559512
rect 128648 559026 128676 559506
rect 128636 559020 128688 559026
rect 128636 558962 128688 558968
rect 128544 537600 128596 537606
rect 128544 537542 128596 537548
rect 128452 484424 128504 484430
rect 128452 484366 128504 484372
rect 128360 480208 128412 480214
rect 128360 480150 128412 480156
rect 128372 479534 128400 480150
rect 128360 479528 128412 479534
rect 128360 479470 128412 479476
rect 128360 474700 128412 474706
rect 128360 474642 128412 474648
rect 127254 460184 127310 460193
rect 127254 460119 127310 460128
rect 127164 442876 127216 442882
rect 127164 442818 127216 442824
rect 127440 442876 127492 442882
rect 127440 442818 127492 442824
rect 127452 442270 127480 442818
rect 127440 442264 127492 442270
rect 127440 442206 127492 442212
rect 127164 402348 127216 402354
rect 127164 402290 127216 402296
rect 127072 389156 127124 389162
rect 127072 389098 127124 389104
rect 127072 368552 127124 368558
rect 127072 368494 127124 368500
rect 126980 349920 127032 349926
rect 126980 349862 127032 349868
rect 126244 349852 126296 349858
rect 126244 349794 126296 349800
rect 125876 339244 125928 339250
rect 125876 339186 125928 339192
rect 125784 337884 125836 337890
rect 125784 337826 125836 337832
rect 126888 337884 126940 337890
rect 126888 337826 126940 337832
rect 126900 337414 126928 337826
rect 126888 337408 126940 337414
rect 126888 337350 126940 337356
rect 126980 336660 127032 336666
rect 126980 336602 127032 336608
rect 126992 336054 127020 336602
rect 126980 336048 127032 336054
rect 126980 335990 127032 335996
rect 125784 332580 125836 332586
rect 125784 332522 125836 332528
rect 125796 332489 125824 332522
rect 125782 332480 125838 332489
rect 125782 332415 125838 332424
rect 125692 320884 125744 320890
rect 125692 320826 125744 320832
rect 125784 312656 125836 312662
rect 125784 312598 125836 312604
rect 126888 312656 126940 312662
rect 126888 312598 126940 312604
rect 125692 293344 125744 293350
rect 125692 293286 125744 293292
rect 125600 263560 125652 263566
rect 125600 263502 125652 263508
rect 125508 254584 125560 254590
rect 125508 254526 125560 254532
rect 125704 244254 125732 293286
rect 125796 274650 125824 312598
rect 126900 311914 126928 312598
rect 126888 311908 126940 311914
rect 126888 311850 126940 311856
rect 125876 300348 125928 300354
rect 125876 300290 125928 300296
rect 125888 286958 125916 300290
rect 125876 286952 125928 286958
rect 125876 286894 125928 286900
rect 125888 286346 125916 286894
rect 125876 286340 125928 286346
rect 125876 286282 125928 286288
rect 125784 274644 125836 274650
rect 125784 274586 125836 274592
rect 126992 273222 127020 335990
rect 127084 318306 127112 368494
rect 127176 339182 127204 402290
rect 127256 396840 127308 396846
rect 127256 396782 127308 396788
rect 127164 339176 127216 339182
rect 127164 339118 127216 339124
rect 127268 333946 127296 396782
rect 128372 367810 128400 474642
rect 128464 380866 128492 484366
rect 128556 438802 128584 537542
rect 128648 466410 128676 558962
rect 129016 553450 129044 643078
rect 136652 596834 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 155224 700392 155276 700398
rect 155224 700334 155276 700340
rect 136640 596828 136692 596834
rect 136640 596770 136692 596776
rect 155236 587178 155264 700334
rect 170324 697610 170352 703520
rect 202800 703254 202828 703520
rect 201500 703248 201552 703254
rect 201500 703190 201552 703196
rect 202788 703248 202840 703254
rect 202788 703190 202840 703196
rect 170312 697604 170364 697610
rect 170312 697546 170364 697552
rect 133236 587172 133288 587178
rect 133236 587114 133288 587120
rect 155224 587172 155276 587178
rect 155224 587114 155276 587120
rect 133248 586566 133276 587114
rect 133236 586560 133288 586566
rect 133236 586502 133288 586508
rect 129740 582548 129792 582554
rect 129740 582490 129792 582496
rect 129004 553444 129056 553450
rect 129004 553386 129056 553392
rect 129752 493950 129780 582490
rect 129832 575544 129884 575550
rect 129832 575486 129884 575492
rect 129740 493944 129792 493950
rect 129740 493886 129792 493892
rect 129752 493338 129780 493886
rect 129740 493332 129792 493338
rect 129740 493274 129792 493280
rect 129844 484401 129872 575486
rect 131764 573368 131816 573374
rect 131764 573310 131816 573316
rect 131028 564460 131080 564466
rect 131028 564402 131080 564408
rect 130016 494760 130068 494766
rect 130016 494702 130068 494708
rect 129830 484392 129886 484401
rect 129830 484327 129886 484336
rect 129924 468580 129976 468586
rect 129924 468522 129976 468528
rect 128636 466404 128688 466410
rect 128636 466346 128688 466352
rect 129832 454028 129884 454034
rect 129832 453970 129884 453976
rect 128544 438796 128596 438802
rect 128544 438738 128596 438744
rect 128452 380860 128504 380866
rect 128452 380802 128504 380808
rect 128464 379574 128492 380802
rect 128452 379568 128504 379574
rect 128452 379510 128504 379516
rect 128452 376100 128504 376106
rect 128452 376042 128504 376048
rect 128360 367804 128412 367810
rect 128360 367746 128412 367752
rect 128360 356788 128412 356794
rect 128360 356730 128412 356736
rect 128372 335238 128400 356730
rect 128464 351354 128492 376042
rect 128452 351348 128504 351354
rect 128452 351290 128504 351296
rect 128450 338056 128506 338065
rect 128450 337991 128506 338000
rect 128464 337958 128492 337991
rect 128452 337952 128504 337958
rect 128452 337894 128504 337900
rect 128464 336802 128492 337894
rect 128452 336796 128504 336802
rect 128452 336738 128504 336744
rect 128556 336666 128584 438738
rect 128636 387184 128688 387190
rect 128636 387126 128688 387132
rect 128648 386510 128676 387126
rect 128636 386504 128688 386510
rect 128636 386446 128688 386452
rect 128544 336660 128596 336666
rect 128544 336602 128596 336608
rect 128360 335232 128412 335238
rect 128360 335174 128412 335180
rect 127256 333940 127308 333946
rect 127256 333882 127308 333888
rect 128648 333334 128676 386446
rect 129740 379568 129792 379574
rect 129740 379510 129792 379516
rect 128728 342984 128780 342990
rect 128728 342926 128780 342932
rect 128740 342310 128768 342926
rect 128728 342304 128780 342310
rect 128728 342246 128780 342252
rect 128636 333328 128688 333334
rect 128636 333270 128688 333276
rect 128452 332580 128504 332586
rect 128452 332522 128504 332528
rect 127072 318300 127124 318306
rect 127072 318242 127124 318248
rect 127164 298784 127216 298790
rect 127164 298726 127216 298732
rect 127070 296168 127126 296177
rect 127070 296103 127126 296112
rect 126980 273216 127032 273222
rect 126980 273158 127032 273164
rect 125692 244248 125744 244254
rect 125692 244190 125744 244196
rect 127084 237318 127112 296103
rect 127176 259350 127204 298726
rect 127164 259344 127216 259350
rect 127164 259286 127216 259292
rect 128464 238754 128492 332522
rect 128544 324284 128596 324290
rect 128544 324226 128596 324232
rect 128556 256698 128584 324226
rect 128544 256692 128596 256698
rect 128544 256634 128596 256640
rect 128372 238726 128492 238754
rect 127072 237312 127124 237318
rect 127072 237254 127124 237260
rect 124312 235952 124364 235958
rect 124312 235894 124364 235900
rect 128372 230450 128400 238726
rect 128740 238610 128768 342246
rect 129752 242826 129780 379510
rect 129844 342990 129872 453970
rect 129936 360126 129964 468522
rect 130028 392698 130056 494702
rect 130108 494012 130160 494018
rect 130108 493954 130160 493960
rect 130016 392692 130068 392698
rect 130016 392634 130068 392640
rect 130120 389978 130148 493954
rect 131040 474586 131068 564402
rect 131120 550656 131172 550662
rect 131120 550598 131172 550604
rect 131132 485081 131160 550598
rect 131212 493944 131264 493950
rect 131212 493886 131264 493892
rect 131118 485072 131174 485081
rect 131118 485007 131174 485016
rect 131040 474558 131160 474586
rect 131132 472802 131160 474558
rect 131120 472796 131172 472802
rect 131120 472738 131172 472744
rect 130108 389972 130160 389978
rect 130108 389914 130160 389920
rect 130016 383716 130068 383722
rect 130016 383658 130068 383664
rect 129924 360120 129976 360126
rect 129924 360062 129976 360068
rect 129832 342984 129884 342990
rect 129832 342926 129884 342932
rect 129832 328432 129884 328438
rect 129830 328400 129832 328409
rect 129884 328400 129886 328409
rect 129830 328335 129886 328344
rect 129832 304360 129884 304366
rect 129832 304302 129884 304308
rect 129740 242820 129792 242826
rect 129740 242762 129792 242768
rect 129844 240961 129872 304302
rect 129922 297392 129978 297401
rect 129922 297327 129978 297336
rect 129936 276690 129964 297327
rect 130028 293962 130056 383658
rect 131132 367062 131160 472738
rect 131224 389910 131252 493886
rect 131776 483002 131804 573310
rect 132500 570036 132552 570042
rect 132500 569978 132552 569984
rect 131764 482996 131816 483002
rect 131764 482938 131816 482944
rect 132512 477465 132540 569978
rect 133144 546576 133196 546582
rect 133144 546518 133196 546524
rect 132592 537668 132644 537674
rect 132592 537610 132644 537616
rect 132498 477456 132554 477465
rect 132498 477391 132554 477400
rect 132500 475380 132552 475386
rect 132500 475322 132552 475328
rect 131304 396908 131356 396914
rect 131304 396850 131356 396856
rect 131212 389904 131264 389910
rect 131212 389846 131264 389852
rect 131212 387252 131264 387258
rect 131212 387194 131264 387200
rect 131120 367056 131172 367062
rect 131120 366998 131172 367004
rect 131132 365770 131160 366998
rect 131120 365764 131172 365770
rect 131120 365706 131172 365712
rect 131224 335170 131252 387194
rect 131316 345710 131344 396850
rect 132512 368490 132540 475322
rect 132604 445058 132632 537610
rect 133156 445194 133184 546518
rect 133248 497486 133276 586502
rect 134064 578264 134116 578270
rect 134064 578206 134116 578212
rect 133972 554056 134024 554062
rect 133972 553998 134024 554004
rect 133788 547188 133840 547194
rect 133788 547130 133840 547136
rect 133800 546582 133828 547130
rect 133788 546576 133840 546582
rect 133788 546518 133840 546524
rect 133236 497480 133288 497486
rect 133236 497422 133288 497428
rect 133880 496120 133932 496126
rect 133880 496062 133932 496068
rect 133788 455388 133840 455394
rect 133788 455330 133840 455336
rect 133144 445188 133196 445194
rect 133144 445130 133196 445136
rect 132592 445052 132644 445058
rect 132592 444994 132644 445000
rect 132592 387320 132644 387326
rect 132592 387262 132644 387268
rect 131672 368484 131724 368490
rect 131672 368426 131724 368432
rect 132500 368484 132552 368490
rect 132500 368426 132552 368432
rect 131684 367130 131712 368426
rect 131672 367124 131724 367130
rect 131672 367066 131724 367072
rect 131684 364334 131712 367066
rect 132500 365764 132552 365770
rect 132500 365706 132552 365712
rect 131684 364306 131804 364334
rect 131304 345704 131356 345710
rect 131304 345646 131356 345652
rect 131212 335164 131264 335170
rect 131212 335106 131264 335112
rect 130568 328432 130620 328438
rect 130568 328374 130620 328380
rect 130580 327146 130608 328374
rect 130568 327140 130620 327146
rect 130568 327082 130620 327088
rect 131120 302932 131172 302938
rect 131120 302874 131172 302880
rect 130016 293956 130068 293962
rect 130016 293898 130068 293904
rect 129924 276684 129976 276690
rect 129924 276626 129976 276632
rect 129936 276078 129964 276626
rect 129924 276072 129976 276078
rect 129924 276014 129976 276020
rect 130384 276072 130436 276078
rect 130384 276014 130436 276020
rect 130396 247722 130424 276014
rect 131132 249762 131160 302874
rect 131776 267734 131804 364306
rect 131684 267706 131804 267734
rect 131684 260846 131712 267706
rect 131672 260840 131724 260846
rect 131672 260782 131724 260788
rect 131684 260166 131712 260782
rect 131672 260160 131724 260166
rect 131672 260102 131724 260108
rect 131120 249756 131172 249762
rect 131120 249698 131172 249704
rect 130384 247716 130436 247722
rect 130384 247658 130436 247664
rect 129830 240952 129886 240961
rect 129830 240887 129886 240896
rect 132512 238882 132540 365706
rect 132604 262206 132632 387262
rect 132684 360256 132736 360262
rect 132684 360198 132736 360204
rect 132696 286890 132724 360198
rect 133800 347750 133828 455330
rect 133892 385082 133920 496062
rect 133984 462398 134012 553998
rect 134076 487830 134104 578206
rect 135352 569968 135404 569974
rect 135352 569910 135404 569916
rect 134156 536104 134208 536110
rect 134156 536046 134208 536052
rect 134064 487824 134116 487830
rect 134064 487766 134116 487772
rect 133972 462392 134024 462398
rect 133972 462334 134024 462340
rect 133880 385076 133932 385082
rect 133880 385018 133932 385024
rect 133984 354686 134012 462334
rect 134168 449206 134196 536046
rect 135260 497548 135312 497554
rect 135260 497490 135312 497496
rect 135168 472728 135220 472734
rect 135168 472670 135220 472676
rect 135180 471306 135208 472670
rect 135168 471300 135220 471306
rect 135168 471242 135220 471248
rect 134156 449200 134208 449206
rect 134156 449142 134208 449148
rect 134064 445188 134116 445194
rect 134064 445130 134116 445136
rect 133972 354680 134024 354686
rect 133972 354622 134024 354628
rect 133984 353394 134012 354622
rect 133972 353388 134024 353394
rect 133972 353330 134024 353336
rect 133880 353320 133932 353326
rect 133880 353262 133932 353268
rect 133788 347744 133840 347750
rect 133788 347686 133840 347692
rect 133800 347138 133828 347686
rect 133788 347132 133840 347138
rect 133788 347074 133840 347080
rect 133144 329792 133196 329798
rect 133142 329760 133144 329769
rect 133788 329792 133840 329798
rect 133196 329760 133198 329769
rect 133788 329734 133840 329740
rect 133142 329695 133198 329704
rect 133800 329089 133828 329734
rect 133786 329080 133842 329089
rect 133786 329015 133842 329024
rect 133144 292800 133196 292806
rect 133144 292742 133196 292748
rect 132684 286884 132736 286890
rect 132684 286826 132736 286832
rect 132592 262200 132644 262206
rect 132592 262142 132644 262148
rect 132500 238876 132552 238882
rect 132500 238818 132552 238824
rect 128728 238604 128780 238610
rect 128728 238546 128780 238552
rect 128360 230444 128412 230450
rect 128360 230386 128412 230392
rect 128372 229838 128400 230386
rect 128360 229832 128412 229838
rect 128360 229774 128412 229780
rect 123484 211880 123536 211886
rect 123484 211822 123536 211828
rect 120080 202836 120132 202842
rect 120080 202778 120132 202784
rect 133156 200870 133184 292742
rect 133892 238474 133920 353262
rect 134076 336598 134104 445130
rect 135272 390046 135300 497490
rect 135364 474065 135392 569910
rect 136824 563780 136876 563786
rect 136824 563722 136876 563728
rect 136640 552084 136692 552090
rect 136640 552026 136692 552032
rect 135444 545148 135496 545154
rect 135444 545090 135496 545096
rect 135350 474056 135406 474065
rect 135350 473991 135406 474000
rect 135456 457473 135484 545090
rect 136652 459542 136680 552026
rect 136732 544400 136784 544406
rect 136732 544342 136784 544348
rect 136640 459536 136692 459542
rect 136640 459478 136692 459484
rect 135442 457464 135498 457473
rect 135442 457399 135498 457408
rect 136744 452606 136772 544342
rect 136836 472666 136864 563722
rect 139492 560312 139544 560318
rect 139492 560254 139544 560260
rect 138112 558952 138164 558958
rect 138112 558894 138164 558900
rect 138020 497480 138072 497486
rect 138020 497422 138072 497428
rect 136824 472660 136876 472666
rect 136824 472602 136876 472608
rect 136824 463752 136876 463758
rect 136824 463694 136876 463700
rect 136732 452600 136784 452606
rect 136732 452542 136784 452548
rect 136732 445052 136784 445058
rect 136732 444994 136784 445000
rect 135352 399492 135404 399498
rect 135352 399434 135404 399440
rect 135260 390040 135312 390046
rect 135260 389982 135312 389988
rect 134156 389904 134208 389910
rect 134156 389846 134208 389852
rect 134064 336592 134116 336598
rect 134064 336534 134116 336540
rect 133970 323776 134026 323785
rect 133970 323711 134026 323720
rect 133984 264926 134012 323711
rect 134168 301510 134196 389846
rect 135260 386368 135312 386374
rect 135260 386310 135312 386316
rect 134614 385656 134670 385665
rect 134614 385591 134670 385600
rect 134628 385082 134656 385591
rect 135272 385150 135300 386310
rect 135260 385144 135312 385150
rect 135260 385086 135312 385092
rect 134616 385076 134668 385082
rect 134616 385018 134668 385024
rect 134156 301504 134208 301510
rect 134156 301446 134208 301452
rect 133972 264920 134024 264926
rect 133972 264862 134024 264868
rect 133880 238468 133932 238474
rect 133880 238410 133932 238416
rect 135272 234530 135300 385086
rect 135364 320142 135392 399434
rect 135444 392624 135496 392630
rect 135444 392566 135496 392572
rect 135456 333878 135484 392566
rect 136640 386436 136692 386442
rect 136640 386378 136692 386384
rect 135444 333872 135496 333878
rect 135444 333814 135496 333820
rect 135456 333266 135484 333814
rect 135444 333260 135496 333266
rect 135444 333202 135496 333208
rect 135352 320136 135404 320142
rect 135352 320078 135404 320084
rect 136548 320136 136600 320142
rect 136548 320078 136600 320084
rect 136560 319530 136588 320078
rect 136548 319524 136600 319530
rect 136548 319466 136600 319472
rect 136652 237386 136680 386378
rect 136744 335306 136772 444994
rect 136836 353326 136864 463694
rect 137100 452600 137152 452606
rect 137100 452542 137152 452548
rect 137112 451314 137140 452542
rect 137100 451308 137152 451314
rect 137100 451250 137152 451256
rect 136916 439136 136968 439142
rect 136916 439078 136968 439084
rect 136824 353320 136876 353326
rect 136824 353262 136876 353268
rect 136732 335300 136784 335306
rect 136732 335242 136784 335248
rect 136928 331226 136956 439078
rect 138032 386374 138060 497422
rect 138124 468518 138152 558894
rect 139400 549364 139452 549370
rect 139400 549306 139452 549312
rect 138112 468512 138164 468518
rect 138112 468454 138164 468460
rect 139412 455394 139440 549306
rect 139504 470626 139532 560254
rect 201512 559570 201540 703190
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 595474 266400 697546
rect 266360 595468 266412 595474
rect 266360 595410 266412 595416
rect 282932 585818 282960 702406
rect 282920 585812 282972 585818
rect 282920 585754 282972 585760
rect 201500 559564 201552 559570
rect 201500 559506 201552 559512
rect 140964 549296 141016 549302
rect 140964 549238 141016 549244
rect 140780 541000 140832 541006
rect 140780 540942 140832 540948
rect 139492 470620 139544 470626
rect 139492 470562 139544 470568
rect 139400 455388 139452 455394
rect 139400 455330 139452 455336
rect 138112 440292 138164 440298
rect 138112 440234 138164 440240
rect 138020 386368 138072 386374
rect 138020 386310 138072 386316
rect 138020 353388 138072 353394
rect 138020 353330 138072 353336
rect 136916 331220 136968 331226
rect 136916 331162 136968 331168
rect 137192 331220 137244 331226
rect 137192 331162 137244 331168
rect 137204 330546 137232 331162
rect 137192 330540 137244 330546
rect 137192 330482 137244 330488
rect 138032 238649 138060 353330
rect 138124 327826 138152 440234
rect 138204 399560 138256 399566
rect 138204 399502 138256 399508
rect 138112 327820 138164 327826
rect 138112 327762 138164 327768
rect 138216 320074 138244 399502
rect 139400 390652 139452 390658
rect 139400 390594 139452 390600
rect 138204 320068 138256 320074
rect 138204 320010 138256 320016
rect 138664 320068 138716 320074
rect 138664 320010 138716 320016
rect 138676 319462 138704 320010
rect 138664 319456 138716 319462
rect 138664 319398 138716 319404
rect 139412 238814 139440 390594
rect 139504 362234 139532 470562
rect 140792 450566 140820 540942
rect 140872 472660 140924 472666
rect 140872 472602 140924 472608
rect 140780 450560 140832 450566
rect 140780 450502 140832 450508
rect 140792 449954 140820 450502
rect 140780 449948 140832 449954
rect 140780 449890 140832 449896
rect 140780 449200 140832 449206
rect 140780 449142 140832 449148
rect 139584 441652 139636 441658
rect 139584 441594 139636 441600
rect 139492 362228 139544 362234
rect 139492 362170 139544 362176
rect 139596 336734 139624 441594
rect 140792 339590 140820 449142
rect 140884 365158 140912 472602
rect 140976 458862 141004 549238
rect 299492 547194 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703186 332548 703520
rect 332508 703180 332560 703186
rect 332508 703122 332560 703128
rect 348804 702545 348832 703520
rect 364996 703050 365024 703520
rect 397472 703118 397500 703520
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 527192 702574 527220 703520
rect 527180 702568 527232 702574
rect 348790 702536 348846 702545
rect 527180 702510 527232 702516
rect 543476 702506 543504 703520
rect 559668 702642 559696 703520
rect 559656 702636 559708 702642
rect 559656 702578 559708 702584
rect 348790 702471 348846 702480
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 411904 616888 411956 616894
rect 411904 616830 411956 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 386328 582412 386380 582418
rect 386328 582354 386380 582360
rect 386340 578202 386368 582354
rect 386328 578196 386380 578202
rect 386328 578138 386380 578144
rect 299480 547188 299532 547194
rect 299480 547130 299532 547136
rect 142344 546508 142396 546514
rect 142344 546450 142396 546456
rect 142160 542428 142212 542434
rect 142160 542370 142212 542376
rect 140964 458856 141016 458862
rect 140964 458798 141016 458804
rect 142172 451926 142200 542370
rect 142252 465112 142304 465118
rect 142252 465054 142304 465060
rect 142160 451920 142212 451926
rect 142160 451862 142212 451868
rect 141056 398132 141108 398138
rect 141056 398074 141108 398080
rect 140964 392692 141016 392698
rect 140964 392634 141016 392640
rect 140872 365152 140924 365158
rect 140872 365094 140924 365100
rect 140872 347880 140924 347886
rect 140872 347822 140924 347828
rect 140884 347750 140912 347822
rect 140872 347744 140924 347750
rect 140872 347686 140924 347692
rect 140870 341456 140926 341465
rect 140870 341391 140926 341400
rect 140884 340950 140912 341391
rect 140872 340944 140924 340950
rect 140872 340886 140924 340892
rect 140780 339584 140832 339590
rect 140780 339526 140832 339532
rect 139584 336728 139636 336734
rect 139584 336670 139636 336676
rect 139400 238808 139452 238814
rect 139400 238750 139452 238756
rect 138018 238640 138074 238649
rect 138018 238575 138074 238584
rect 136640 237380 136692 237386
rect 136640 237322 136692 237328
rect 140884 235890 140912 340886
rect 140976 288386 141004 392634
rect 141068 338026 141096 398074
rect 142160 394868 142212 394874
rect 142160 394810 142212 394816
rect 141056 338020 141108 338026
rect 141056 337962 141108 337968
rect 141332 338020 141384 338026
rect 141332 337962 141384 337968
rect 141344 337482 141372 337962
rect 141332 337476 141384 337482
rect 141332 337418 141384 337424
rect 141424 295724 141476 295730
rect 141424 295666 141476 295672
rect 140964 288380 141016 288386
rect 140964 288322 141016 288328
rect 140872 235884 140924 235890
rect 140872 235826 140924 235832
rect 135260 234524 135312 234530
rect 135260 234466 135312 234472
rect 133880 226296 133932 226302
rect 133878 226264 133880 226273
rect 135168 226296 135220 226302
rect 133932 226264 133934 226273
rect 135168 226238 135220 226244
rect 133878 226199 133934 226208
rect 135180 225010 135208 226238
rect 135168 225004 135220 225010
rect 135168 224946 135220 224952
rect 133144 200864 133196 200870
rect 133144 200806 133196 200812
rect 141436 191049 141464 295666
rect 141608 288380 141660 288386
rect 141608 288322 141660 288328
rect 141620 287706 141648 288322
rect 141608 287700 141660 287706
rect 141608 287642 141660 287648
rect 142172 242894 142200 394810
rect 142264 356046 142292 465054
rect 142356 458930 142384 546450
rect 411916 538898 411944 616830
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579804 578196 579856 578202
rect 579804 578138 579856 578144
rect 579816 577697 579844 578138
rect 579802 577688 579858 577697
rect 579802 577623 579858 577632
rect 413284 564460 413336 564466
rect 413284 564402 413336 564408
rect 413296 538898 413324 564402
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563718 580212 564295
rect 580172 563712 580224 563718
rect 580172 563654 580224 563660
rect 580276 541686 580304 630799
rect 580264 541680 580316 541686
rect 580264 541622 580316 541628
rect 411904 538892 411956 538898
rect 411904 538834 411956 538840
rect 413284 538892 413336 538898
rect 413284 538834 413336 538840
rect 580908 538892 580960 538898
rect 580908 538834 580960 538840
rect 580920 537849 580948 538834
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580356 492720 580408 492726
rect 580356 492662 580408 492668
rect 143540 491972 143592 491978
rect 143540 491914 143592 491920
rect 142344 458924 142396 458930
rect 142344 458866 142396 458872
rect 142344 451308 142396 451314
rect 142344 451250 142396 451256
rect 142252 356040 142304 356046
rect 142252 355982 142304 355988
rect 142356 341562 142384 451250
rect 142436 389224 142488 389230
rect 142436 389166 142488 389172
rect 142344 341556 142396 341562
rect 142344 341498 142396 341504
rect 142448 292466 142476 389166
rect 143552 387190 143580 491914
rect 580264 490612 580316 490618
rect 580264 490554 580316 490560
rect 145012 487824 145064 487830
rect 145012 487766 145064 487772
rect 143632 449948 143684 449954
rect 143632 449890 143684 449896
rect 143540 387184 143592 387190
rect 143540 387126 143592 387132
rect 143540 376032 143592 376038
rect 143540 375974 143592 375980
rect 143448 356040 143500 356046
rect 143448 355982 143500 355988
rect 143460 355366 143488 355982
rect 143448 355360 143500 355366
rect 143448 355302 143500 355308
rect 142436 292460 142488 292466
rect 142436 292402 142488 292408
rect 142160 242888 142212 242894
rect 142160 242830 142212 242836
rect 143552 233238 143580 375974
rect 143644 339658 143672 449890
rect 144920 448588 144972 448594
rect 144920 448530 144972 448536
rect 143816 442264 143868 442270
rect 143816 442206 143868 442212
rect 143724 390584 143776 390590
rect 143724 390526 143776 390532
rect 143632 339652 143684 339658
rect 143632 339594 143684 339600
rect 143736 284306 143764 390526
rect 143828 338094 143856 442206
rect 144932 339318 144960 448530
rect 145024 382226 145052 487766
rect 146484 483064 146536 483070
rect 146484 483006 146536 483012
rect 146392 458924 146444 458930
rect 146392 458866 146444 458872
rect 146300 389972 146352 389978
rect 146300 389914 146352 389920
rect 145012 382220 145064 382226
rect 145012 382162 145064 382168
rect 145024 381546 145052 382162
rect 145012 381540 145064 381546
rect 145012 381482 145064 381488
rect 144920 339312 144972 339318
rect 144920 339254 144972 339260
rect 143816 338088 143868 338094
rect 143816 338030 143868 338036
rect 145564 307964 145616 307970
rect 145564 307906 145616 307912
rect 143724 284300 143776 284306
rect 143724 284242 143776 284248
rect 143540 233232 143592 233238
rect 143540 233174 143592 233180
rect 142804 220176 142856 220182
rect 142804 220118 142856 220124
rect 142816 192574 142844 220118
rect 145576 194138 145604 307906
rect 146312 269074 146340 389914
rect 146404 346390 146432 458866
rect 146496 377466 146524 483006
rect 151912 479528 151964 479534
rect 151912 479470 151964 479476
rect 147772 471300 147824 471306
rect 147772 471242 147824 471248
rect 147784 470626 147812 471242
rect 151818 471200 151874 471209
rect 151818 471135 151874 471144
rect 147772 470620 147824 470626
rect 147772 470562 147824 470568
rect 147680 468512 147732 468518
rect 147680 468454 147732 468460
rect 146484 377460 146536 377466
rect 146484 377402 146536 377408
rect 147692 360194 147720 468454
rect 147784 365090 147812 470562
rect 149152 458856 149204 458862
rect 149152 458798 149204 458804
rect 149058 456104 149114 456113
rect 149058 456039 149114 456048
rect 147864 391264 147916 391270
rect 147864 391206 147916 391212
rect 147772 365084 147824 365090
rect 147772 365026 147824 365032
rect 147680 360188 147732 360194
rect 147680 360130 147732 360136
rect 147692 359514 147720 360130
rect 147680 359508 147732 359514
rect 147680 359450 147732 359456
rect 146392 346384 146444 346390
rect 146392 346326 146444 346332
rect 146760 346384 146812 346390
rect 146760 346326 146812 346332
rect 146772 345710 146800 346326
rect 146760 345704 146812 345710
rect 146760 345646 146812 345652
rect 147876 292534 147904 391206
rect 149072 345030 149100 456039
rect 149164 364334 149192 458798
rect 150438 457464 150494 457473
rect 150438 457399 150494 457408
rect 149164 364306 149284 364334
rect 149256 347750 149284 364306
rect 149244 347744 149296 347750
rect 149244 347686 149296 347692
rect 149256 347070 149284 347686
rect 149244 347064 149296 347070
rect 149244 347006 149296 347012
rect 149060 345024 149112 345030
rect 149060 344966 149112 344972
rect 149072 344350 149100 344966
rect 149060 344344 149112 344350
rect 149060 344286 149112 344292
rect 150452 343602 150480 457399
rect 150532 451920 150584 451926
rect 150532 451862 150584 451868
rect 150440 343596 150492 343602
rect 150440 343538 150492 343544
rect 150452 342922 150480 343538
rect 150440 342916 150492 342922
rect 150440 342858 150492 342864
rect 150544 340882 150572 451862
rect 151832 362914 151860 471135
rect 151924 375358 151952 479470
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580276 458153 580304 490554
rect 580368 484673 580396 492662
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 431254 580212 431559
rect 580172 431248 580224 431254
rect 580172 431190 580224 431196
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 160742 401704 160798 401713
rect 160742 401639 160798 401648
rect 152004 393440 152056 393446
rect 152004 393382 152056 393388
rect 151912 375352 151964 375358
rect 151912 375294 151964 375300
rect 151820 362908 151872 362914
rect 151820 362850 151872 362856
rect 150532 340876 150584 340882
rect 150532 340818 150584 340824
rect 151544 340876 151596 340882
rect 151544 340818 151596 340824
rect 151556 340202 151584 340818
rect 151544 340196 151596 340202
rect 151544 340138 151596 340144
rect 152016 315994 152044 393382
rect 159364 393372 159416 393378
rect 159364 393314 159416 393320
rect 153108 375352 153160 375358
rect 153108 375294 153160 375300
rect 153120 374678 153148 375294
rect 153108 374672 153160 374678
rect 153108 374614 153160 374620
rect 153108 362908 153160 362914
rect 153108 362850 153160 362856
rect 153120 362273 153148 362850
rect 153106 362264 153162 362273
rect 153106 362199 153162 362208
rect 152004 315988 152056 315994
rect 152004 315930 152056 315936
rect 152016 315314 152044 315930
rect 152004 315308 152056 315314
rect 152004 315250 152056 315256
rect 155224 307896 155276 307902
rect 155224 307838 155276 307844
rect 151084 296948 151136 296954
rect 151084 296890 151136 296896
rect 147864 292528 147916 292534
rect 147864 292470 147916 292476
rect 146300 269068 146352 269074
rect 146300 269010 146352 269016
rect 151096 202162 151124 296890
rect 152464 294228 152516 294234
rect 152464 294170 152516 294176
rect 151084 202156 151136 202162
rect 151084 202098 151136 202104
rect 152476 200802 152504 294170
rect 152464 200796 152516 200802
rect 152464 200738 152516 200744
rect 145564 194132 145616 194138
rect 145564 194074 145616 194080
rect 142804 192568 142856 192574
rect 142804 192510 142856 192516
rect 141422 191040 141478 191049
rect 141422 190975 141478 190984
rect 155236 186998 155264 307838
rect 157984 298444 158036 298450
rect 157984 298386 158036 298392
rect 157996 198082 158024 298386
rect 157984 198076 158036 198082
rect 157984 198018 158036 198024
rect 155224 186992 155276 186998
rect 155224 186934 155276 186940
rect 128268 186448 128320 186454
rect 128268 186390 128320 186396
rect 119988 185020 120040 185026
rect 119988 184962 120040 184968
rect 115940 184340 115992 184346
rect 115940 184282 115992 184288
rect 118424 182300 118476 182306
rect 118424 182242 118476 182248
rect 115848 178220 115900 178226
rect 115848 178162 115900 178168
rect 114098 177712 114154 177721
rect 114098 177647 114154 177656
rect 114466 177712 114522 177721
rect 114466 177647 114522 177656
rect 115860 176769 115888 178162
rect 118436 177721 118464 182242
rect 120000 177721 120028 184962
rect 122656 180940 122708 180946
rect 122656 180882 122708 180888
rect 122668 177721 122696 180882
rect 126796 179444 126848 179450
rect 126796 179386 126848 179392
rect 123760 178288 123812 178294
rect 123760 178230 123812 178236
rect 118422 177712 118478 177721
rect 118422 177647 118478 177656
rect 119986 177712 120042 177721
rect 119986 177647 120042 177656
rect 122654 177712 122710 177721
rect 122654 177647 122710 177656
rect 123772 176769 123800 178230
rect 126808 177041 126836 179386
rect 128280 177721 128308 186390
rect 159376 183122 159404 393314
rect 159364 183116 159416 183122
rect 159364 183058 159416 183064
rect 129464 181008 129516 181014
rect 129464 180950 129516 180956
rect 129476 177721 129504 180950
rect 133144 179512 133196 179518
rect 133144 179454 133196 179460
rect 132408 178356 132460 178362
rect 132408 178298 132460 178304
rect 130752 178084 130804 178090
rect 130752 178026 130804 178032
rect 128266 177712 128322 177721
rect 128266 177647 128322 177656
rect 129462 177712 129518 177721
rect 129462 177647 129518 177656
rect 128176 177064 128228 177070
rect 126794 177032 126850 177041
rect 128176 177006 128228 177012
rect 126794 176967 126850 176976
rect 128188 176769 128216 177006
rect 130764 176769 130792 178026
rect 132420 176769 132448 178298
rect 133156 177041 133184 179454
rect 134800 178424 134852 178430
rect 134800 178366 134852 178372
rect 133142 177032 133198 177041
rect 133142 176967 133198 176976
rect 134812 176769 134840 178366
rect 148232 178152 148284 178158
rect 148232 178094 148284 178100
rect 136088 176792 136140 176798
rect 115846 176760 115902 176769
rect 115846 176695 115902 176704
rect 123758 176760 123814 176769
rect 123758 176695 123814 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 130750 176760 130806 176769
rect 130750 176695 130806 176704
rect 132406 176760 132462 176769
rect 132406 176695 132462 176704
rect 134798 176760 134854 176769
rect 134798 176695 134854 176704
rect 136086 176760 136088 176769
rect 148244 176769 148272 178094
rect 160756 177449 160784 401639
rect 264242 400344 264298 400353
rect 264242 400279 264298 400288
rect 162124 400240 162176 400246
rect 162124 400182 162176 400188
rect 162136 180266 162164 400182
rect 220084 397588 220136 397594
rect 220084 397530 220136 397536
rect 166264 396092 166316 396098
rect 166264 396034 166316 396040
rect 163504 303816 163556 303822
rect 163504 303758 163556 303764
rect 163516 205086 163544 303758
rect 164882 291952 164938 291961
rect 164882 291887 164938 291896
rect 163504 205080 163556 205086
rect 163504 205022 163556 205028
rect 164896 181393 164924 291887
rect 164882 181384 164938 181393
rect 164882 181319 164938 181328
rect 166276 180334 166304 396034
rect 170404 394800 170456 394806
rect 170404 394742 170456 394748
rect 169024 303748 169076 303754
rect 169024 303690 169076 303696
rect 166356 291916 166408 291922
rect 166356 291858 166408 291864
rect 166368 199646 166396 291858
rect 166356 199640 166408 199646
rect 166356 199582 166408 199588
rect 167644 183592 167696 183598
rect 167644 183534 167696 183540
rect 166356 182300 166408 182306
rect 166356 182242 166408 182248
rect 166264 180328 166316 180334
rect 166264 180270 166316 180276
rect 162124 180260 162176 180266
rect 162124 180202 162176 180208
rect 165068 179512 165120 179518
rect 165068 179454 165120 179460
rect 160742 177440 160798 177449
rect 160742 177375 160798 177384
rect 164424 176996 164476 177002
rect 164424 176938 164476 176944
rect 136140 176760 136142 176769
rect 136086 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158904 176316 158956 176322
rect 158904 176258 158956 176264
rect 124496 176112 124548 176118
rect 124496 176054 124548 176060
rect 120816 176044 120868 176050
rect 120816 175986 120868 175992
rect 111064 175976 111116 175982
rect 111064 175918 111116 175924
rect 116952 175976 117004 175982
rect 116952 175918 117004 175924
rect 116964 175545 116992 175918
rect 120828 175545 120856 175986
rect 124508 175545 124536 176054
rect 158916 175545 158944 176258
rect 164436 176254 164464 176938
rect 164424 176248 164476 176254
rect 164424 176190 164476 176196
rect 116950 175536 117006 175545
rect 116950 175471 117006 175480
rect 120814 175536 120870 175545
rect 120814 175471 120870 175480
rect 124494 175536 124550 175545
rect 124494 175471 124550 175480
rect 158902 175536 158958 175545
rect 158902 175471 158958 175480
rect 110694 175400 110750 175409
rect 110694 175335 110750 175344
rect 165080 175234 165108 179454
rect 165528 178424 165580 178430
rect 165528 178366 165580 178372
rect 165436 178356 165488 178362
rect 165436 178298 165488 178304
rect 165068 175228 165120 175234
rect 165068 175170 165120 175176
rect 165448 173874 165476 178298
rect 165540 175166 165568 178366
rect 166264 176316 166316 176322
rect 166264 176258 166316 176264
rect 165528 175160 165580 175166
rect 165528 175102 165580 175108
rect 165436 173868 165488 173874
rect 165436 173810 165488 173816
rect 166276 149054 166304 176258
rect 166368 166870 166396 182242
rect 166448 181008 166500 181014
rect 166448 180950 166500 180956
rect 166460 172514 166488 180950
rect 166540 179444 166592 179450
rect 166540 179386 166592 179392
rect 166448 172508 166500 172514
rect 166448 172450 166500 172456
rect 166552 171086 166580 179386
rect 167550 171592 167606 171601
rect 167550 171527 167606 171536
rect 167564 171358 167592 171527
rect 167552 171352 167604 171358
rect 167552 171294 167604 171300
rect 166540 171080 166592 171086
rect 166540 171022 166592 171028
rect 166356 166864 166408 166870
rect 166356 166806 166408 166812
rect 167656 157350 167684 183534
rect 167920 180940 167972 180946
rect 167920 180882 167972 180888
rect 167828 178220 167880 178226
rect 167828 178162 167880 178168
rect 167736 176860 167788 176866
rect 167736 176802 167788 176808
rect 167748 160750 167776 176802
rect 167840 165578 167868 178162
rect 167932 168366 167960 180882
rect 169036 178838 169064 303690
rect 169116 182232 169168 182238
rect 169116 182174 169168 182180
rect 169024 178832 169076 178838
rect 169024 178774 169076 178780
rect 169024 176928 169076 176934
rect 169024 176870 169076 176876
rect 167920 168360 167972 168366
rect 167920 168302 167972 168308
rect 167828 165572 167880 165578
rect 167828 165514 167880 165520
rect 167736 160744 167788 160750
rect 167736 160686 167788 160692
rect 169036 160070 169064 176870
rect 169024 160064 169076 160070
rect 169024 160006 169076 160012
rect 167644 157344 167696 157350
rect 167644 157286 167696 157292
rect 169128 155922 169156 182174
rect 169208 180872 169260 180878
rect 169208 180814 169260 180820
rect 169220 164218 169248 180814
rect 169300 178288 169352 178294
rect 169300 178230 169352 178236
rect 169312 169726 169340 178230
rect 169760 177064 169812 177070
rect 169760 177006 169812 177012
rect 169772 172446 169800 177006
rect 169760 172440 169812 172446
rect 169760 172382 169812 172388
rect 169300 169720 169352 169726
rect 169300 169662 169352 169668
rect 169666 168464 169722 168473
rect 169666 168399 169722 168408
rect 169208 164212 169260 164218
rect 169208 164154 169260 164160
rect 169116 155916 169168 155922
rect 169116 155858 169168 155864
rect 167644 153264 167696 153270
rect 167644 153206 167696 153212
rect 166264 149048 166316 149054
rect 166264 148990 166316 148996
rect 67454 129296 67510 129305
rect 67454 129231 67510 129240
rect 66166 128072 66222 128081
rect 66166 128007 66222 128016
rect 65522 125216 65578 125225
rect 65522 125151 65578 125160
rect 65536 124234 65564 125151
rect 65524 124228 65576 124234
rect 65524 124170 65576 124176
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 66088 91089 66116 122567
rect 66180 94897 66208 128007
rect 67362 120864 67418 120873
rect 67362 120799 67418 120808
rect 66166 94888 66222 94897
rect 66166 94823 66222 94832
rect 66074 91080 66130 91089
rect 66074 91015 66130 91024
rect 67376 89690 67404 120799
rect 67468 93809 67496 129231
rect 67546 126304 67602 126313
rect 67546 126239 67602 126248
rect 67454 93800 67510 93809
rect 67454 93735 67510 93744
rect 67560 91050 67588 126239
rect 166264 125656 166316 125662
rect 166264 125598 166316 125604
rect 67638 102368 67694 102377
rect 67638 102303 67694 102312
rect 67548 91044 67600 91050
rect 67548 90986 67600 90992
rect 67364 89684 67416 89690
rect 67364 89626 67416 89632
rect 67652 85542 67680 102303
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67640 85536 67692 85542
rect 67640 85478 67692 85484
rect 67744 85474 67772 100671
rect 164884 98048 164936 98054
rect 164884 97990 164936 97996
rect 94962 94752 95018 94761
rect 94962 94687 95018 94696
rect 104346 94752 104402 94761
rect 104346 94687 104402 94696
rect 116674 94752 116730 94761
rect 116674 94687 116730 94696
rect 120630 94752 120686 94761
rect 120630 94687 120686 94696
rect 133142 94752 133198 94761
rect 133142 94687 133198 94696
rect 151726 94752 151782 94761
rect 151726 94687 151782 94696
rect 94976 93906 95004 94687
rect 104360 94042 104388 94687
rect 104348 94036 104400 94042
rect 104348 93978 104400 93984
rect 116688 93974 116716 94687
rect 120644 94110 120672 94687
rect 133156 94178 133184 94687
rect 133144 94172 133196 94178
rect 133144 94114 133196 94120
rect 120632 94104 120684 94110
rect 120632 94046 120684 94052
rect 116676 93968 116728 93974
rect 116676 93910 116728 93916
rect 94964 93900 95016 93906
rect 94964 93842 95016 93848
rect 85670 93528 85726 93537
rect 85670 93463 85726 93472
rect 107750 93528 107806 93537
rect 107750 93463 107806 93472
rect 115846 93528 115902 93537
rect 115846 93463 115902 93472
rect 122102 93528 122158 93537
rect 151740 93498 151768 94687
rect 122102 93463 122158 93472
rect 151728 93492 151780 93498
rect 85684 93226 85712 93463
rect 107764 93294 107792 93463
rect 115860 93362 115888 93463
rect 122116 93430 122144 93463
rect 151728 93434 151780 93440
rect 122104 93424 122156 93430
rect 122104 93366 122156 93372
rect 115848 93356 115900 93362
rect 115848 93298 115900 93304
rect 107752 93288 107804 93294
rect 103426 93256 103482 93265
rect 85672 93220 85724 93226
rect 107752 93230 107804 93236
rect 110234 93256 110290 93265
rect 103426 93191 103482 93200
rect 164896 93226 164924 97990
rect 110234 93191 110290 93200
rect 164884 93220 164936 93226
rect 85672 93162 85724 93168
rect 85118 92440 85174 92449
rect 85118 92375 85174 92384
rect 88062 92440 88118 92449
rect 88062 92375 88118 92384
rect 99286 92440 99342 92449
rect 99286 92375 99342 92384
rect 100022 92440 100078 92449
rect 100022 92375 100078 92384
rect 75826 91216 75882 91225
rect 75826 91151 75882 91160
rect 67732 85468 67784 85474
rect 67732 85410 67784 85416
rect 75840 84182 75868 91151
rect 85132 91118 85160 92375
rect 86866 91216 86922 91225
rect 88076 91186 88104 92375
rect 99102 91352 99158 91361
rect 99300 91322 99328 92375
rect 99102 91287 99158 91296
rect 99288 91316 99340 91322
rect 89074 91216 89130 91225
rect 86866 91151 86922 91160
rect 88064 91180 88116 91186
rect 85120 91112 85172 91118
rect 85120 91054 85172 91060
rect 75828 84176 75880 84182
rect 75828 84118 75880 84124
rect 86880 79966 86908 91151
rect 89074 91151 89130 91160
rect 90638 91216 90694 91225
rect 90638 91151 90694 91160
rect 91926 91216 91982 91225
rect 91926 91151 91982 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97078 91216 97134 91225
rect 97078 91151 97134 91160
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 88064 91122 88116 91128
rect 89088 88330 89116 91151
rect 89076 88324 89128 88330
rect 89076 88266 89128 88272
rect 90652 86902 90680 91151
rect 90640 86896 90692 86902
rect 90640 86838 90692 86844
rect 91940 85406 91968 91151
rect 91928 85400 91980 85406
rect 91928 85342 91980 85348
rect 93780 81326 93808 91151
rect 93768 81320 93820 81326
rect 93768 81262 93820 81268
rect 86868 79960 86920 79966
rect 86868 79902 86920 79908
rect 95160 79898 95188 91151
rect 95148 79892 95200 79898
rect 95148 79834 95200 79840
rect 96540 78674 96568 91151
rect 97092 88233 97120 91151
rect 97078 88224 97134 88233
rect 97078 88159 97134 88168
rect 97920 82686 97948 91151
rect 97908 82680 97960 82686
rect 97908 82622 97960 82628
rect 96528 78668 96580 78674
rect 96528 78610 96580 78616
rect 99116 75818 99144 91287
rect 99288 91258 99340 91264
rect 100036 91254 100064 92375
rect 101862 91760 101918 91769
rect 101862 91695 101918 91704
rect 100024 91248 100076 91254
rect 99194 91216 99250 91225
rect 100024 91190 100076 91196
rect 100574 91216 100630 91225
rect 99194 91151 99250 91160
rect 100574 91151 100630 91160
rect 99208 79830 99236 91151
rect 100588 81190 100616 91151
rect 101876 89554 101904 91695
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 101864 89548 101916 89554
rect 101864 89490 101916 89496
rect 101968 84153 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 103334 91216 103390 91225
rect 103334 91151 103390 91160
rect 101954 84144 102010 84153
rect 101954 84079 102010 84088
rect 100576 81184 100628 81190
rect 100576 81126 100628 81132
rect 99196 79824 99248 79830
rect 99196 79766 99248 79772
rect 102060 78577 102088 91151
rect 103348 84114 103376 91151
rect 103336 84108 103388 84114
rect 103336 84050 103388 84056
rect 103440 82618 103468 93191
rect 105726 92440 105782 92449
rect 105726 92375 105728 92384
rect 105780 92375 105782 92384
rect 106830 92440 106886 92449
rect 106830 92375 106886 92384
rect 105728 92346 105780 92352
rect 106844 92206 106872 92375
rect 109682 92304 109738 92313
rect 109682 92239 109738 92248
rect 106832 92200 106884 92206
rect 106832 92142 106884 92148
rect 106924 91316 106976 91322
rect 106924 91258 106976 91264
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 105726 91216 105782 91225
rect 105726 91151 105782 91160
rect 103428 82612 103480 82618
rect 103428 82554 103480 82560
rect 104820 81258 104848 91151
rect 105740 86970 105768 91151
rect 105728 86964 105780 86970
rect 105728 86906 105780 86912
rect 104808 81252 104860 81258
rect 104808 81194 104860 81200
rect 102046 78568 102102 78577
rect 102046 78503 102102 78512
rect 106936 75886 106964 91258
rect 107106 91216 107162 91225
rect 107106 91151 107162 91160
rect 108762 91216 108818 91225
rect 108762 91151 108818 91160
rect 107120 88194 107148 91151
rect 107108 88188 107160 88194
rect 107108 88130 107160 88136
rect 108776 86737 108804 91151
rect 109696 90710 109724 92239
rect 109684 90704 109736 90710
rect 109684 90646 109736 90652
rect 108762 86728 108818 86737
rect 108762 86663 108818 86672
rect 110248 82822 110276 93191
rect 164884 93162 164936 93168
rect 129740 93152 129792 93158
rect 129740 93094 129792 93100
rect 114468 92472 114520 92478
rect 114466 92440 114468 92449
rect 114520 92440 114522 92449
rect 114466 92375 114522 92384
rect 120262 92440 120318 92449
rect 120262 92375 120318 92384
rect 123206 92440 123262 92449
rect 123206 92375 123262 92384
rect 124126 92440 124182 92449
rect 124126 92375 124182 92384
rect 125414 92440 125470 92449
rect 125414 92375 125470 92384
rect 120276 92342 120304 92375
rect 120264 92336 120316 92342
rect 120264 92278 120316 92284
rect 123220 92274 123248 92375
rect 123208 92268 123260 92274
rect 123208 92210 123260 92216
rect 112718 91624 112774 91633
rect 112718 91559 112774 91568
rect 119526 91624 119582 91633
rect 119526 91559 119582 91568
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 111062 91216 111118 91225
rect 111062 91151 111118 91160
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 110236 82816 110288 82822
rect 110236 82758 110288 82764
rect 110340 78470 110368 91151
rect 111076 85338 111104 91151
rect 111064 85332 111116 85338
rect 111064 85274 111116 85280
rect 111720 81394 111748 91151
rect 112732 89486 112760 91559
rect 114466 91352 114522 91361
rect 114466 91287 114522 91296
rect 115846 91352 115902 91361
rect 115846 91287 115902 91296
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 114374 91216 114430 91225
rect 114374 91151 114430 91160
rect 112720 89480 112772 89486
rect 112720 89422 112772 89428
rect 111708 81388 111760 81394
rect 111708 81330 111760 81336
rect 113100 79762 113128 91151
rect 114388 84017 114416 91151
rect 114374 84008 114430 84017
rect 114374 83943 114430 83952
rect 114480 82754 114508 91287
rect 115754 91216 115810 91225
rect 115754 91151 115810 91160
rect 114468 82748 114520 82754
rect 114468 82690 114520 82696
rect 115768 80034 115796 91151
rect 115756 80028 115808 80034
rect 115756 79970 115808 79976
rect 113088 79756 113140 79762
rect 113088 79698 113140 79704
rect 110328 78464 110380 78470
rect 110328 78406 110380 78412
rect 115860 77217 115888 91287
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 118238 91216 118294 91225
rect 118238 91151 118294 91160
rect 117240 84046 117268 91151
rect 118252 88058 118280 91151
rect 119540 89418 119568 91559
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 119710 91216 119766 91225
rect 122286 91216 122342 91225
rect 119710 91151 119766 91160
rect 120080 91180 120132 91186
rect 119528 89412 119580 89418
rect 119528 89354 119580 89360
rect 118240 88052 118292 88058
rect 118240 87994 118292 88000
rect 119724 86834 119752 91151
rect 122286 91151 122342 91160
rect 120080 91122 120132 91128
rect 120092 90914 120120 91122
rect 120080 90908 120132 90914
rect 120080 90850 120132 90856
rect 119712 86828 119764 86834
rect 119712 86770 119764 86776
rect 122300 85202 122328 91151
rect 122852 88262 122880 91423
rect 123484 91248 123536 91254
rect 123484 91190 123536 91196
rect 122840 88256 122892 88262
rect 122840 88198 122892 88204
rect 122288 85196 122340 85202
rect 122288 85138 122340 85144
rect 117228 84040 117280 84046
rect 117228 83982 117280 83988
rect 123496 78538 123524 91190
rect 124140 90846 124168 92375
rect 124128 90840 124180 90846
rect 124128 90782 124180 90788
rect 125428 90778 125456 92375
rect 129752 92206 129780 93094
rect 134430 92440 134486 92449
rect 134430 92375 134486 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152094 92440 152150 92449
rect 152094 92375 152150 92384
rect 134444 92206 134472 92375
rect 129740 92200 129792 92206
rect 129740 92142 129792 92148
rect 134432 92200 134484 92206
rect 134432 92142 134484 92148
rect 126886 91760 126942 91769
rect 126886 91695 126942 91704
rect 126794 91352 126850 91361
rect 126794 91287 126850 91296
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 126702 91216 126758 91225
rect 126702 91151 126758 91160
rect 125416 90772 125468 90778
rect 125416 90714 125468 90720
rect 125520 82550 125548 91151
rect 125508 82544 125560 82550
rect 125508 82486 125560 82492
rect 126716 81122 126744 91151
rect 126808 83978 126836 91287
rect 126900 89622 126928 91695
rect 136270 91624 136326 91633
rect 136270 91559 136326 91568
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 129462 91216 129518 91225
rect 129462 91151 129518 91160
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 126888 89616 126940 89622
rect 126888 89558 126940 89564
rect 126796 83972 126848 83978
rect 126796 83914 126848 83920
rect 126704 81116 126756 81122
rect 126704 81058 126756 81064
rect 128280 78606 128308 91151
rect 129476 87990 129504 91151
rect 129464 87984 129516 87990
rect 129464 87926 129516 87932
rect 130764 85270 130792 91151
rect 132420 86601 132448 91151
rect 133144 91112 133196 91118
rect 133144 91054 133196 91060
rect 132406 86592 132462 86601
rect 132406 86527 132462 86536
rect 130752 85264 130804 85270
rect 130752 85206 130804 85212
rect 128268 78600 128320 78606
rect 128268 78542 128320 78548
rect 123484 78532 123536 78538
rect 123484 78474 123536 78480
rect 133156 77246 133184 91054
rect 136284 89350 136312 91559
rect 136272 89344 136324 89350
rect 136272 89286 136324 89292
rect 151556 88126 151584 92375
rect 152108 92138 152136 92375
rect 152096 92132 152148 92138
rect 152096 92074 152148 92080
rect 151726 91216 151782 91225
rect 151726 91151 151782 91160
rect 151544 88120 151596 88126
rect 151544 88062 151596 88068
rect 151740 86766 151768 91151
rect 166276 90778 166304 125598
rect 166356 111852 166408 111858
rect 166356 111794 166408 111800
rect 166264 90772 166316 90778
rect 166264 90714 166316 90720
rect 151728 86760 151780 86766
rect 151728 86702 151780 86708
rect 166368 81190 166396 111794
rect 166540 99408 166592 99414
rect 166540 99350 166592 99356
rect 166448 98116 166500 98122
rect 166448 98058 166500 98064
rect 166356 81184 166408 81190
rect 166356 81126 166408 81132
rect 166460 79966 166488 98058
rect 166552 88330 166580 99350
rect 167656 93498 167684 153206
rect 167736 142860 167788 142866
rect 167736 142802 167788 142808
rect 167644 93492 167696 93498
rect 167644 93434 167696 93440
rect 167748 92206 167776 142802
rect 169024 140820 169076 140826
rect 169024 140762 169076 140768
rect 167828 122868 167880 122874
rect 167828 122810 167880 122816
rect 167840 94110 167868 122810
rect 168196 113688 168248 113694
rect 168196 113630 168248 113636
rect 168208 110129 168236 113630
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 168194 110120 168250 110129
rect 168194 110055 168250 110064
rect 167920 108996 167972 109002
rect 167920 108938 167972 108944
rect 167932 108769 167960 108938
rect 167918 108760 167974 108769
rect 167918 108695 167974 108704
rect 167920 106344 167972 106350
rect 167920 106286 167972 106292
rect 167828 94104 167880 94110
rect 167828 94046 167880 94052
rect 167736 92200 167788 92206
rect 167736 92142 167788 92148
rect 166540 88324 166592 88330
rect 166540 88266 166592 88272
rect 167932 85406 167960 106286
rect 167920 85400 167972 85406
rect 167920 85342 167972 85348
rect 169036 82550 169064 140762
rect 169116 140072 169168 140078
rect 169116 140014 169168 140020
rect 169128 111790 169156 140014
rect 169680 116618 169708 168399
rect 170416 123486 170444 394742
rect 214564 394732 214616 394738
rect 214564 394674 214616 394680
rect 177304 392012 177356 392018
rect 177304 391954 177356 391960
rect 171784 305040 171836 305046
rect 171784 304982 171836 304988
rect 171796 187105 171824 304982
rect 173900 271924 173952 271930
rect 173900 271866 173952 271872
rect 171876 187808 171928 187814
rect 171876 187750 171928 187756
rect 171782 187096 171838 187105
rect 171782 187031 171838 187040
rect 170496 185020 170548 185026
rect 170496 184962 170548 184968
rect 170508 166938 170536 184962
rect 170588 176180 170640 176186
rect 170588 176122 170640 176128
rect 170496 166932 170548 166938
rect 170496 166874 170548 166880
rect 170600 162858 170628 176122
rect 170680 171352 170732 171358
rect 170680 171294 170732 171300
rect 170588 162852 170640 162858
rect 170588 162794 170640 162800
rect 170692 158030 170720 171294
rect 170680 158024 170732 158030
rect 170680 157966 170732 157972
rect 171888 157282 171916 187750
rect 171968 186448 172020 186454
rect 171968 186390 172020 186396
rect 171980 171018 172008 186390
rect 171968 171012 172020 171018
rect 171968 170954 172020 170960
rect 171876 157276 171928 157282
rect 171876 157218 171928 157224
rect 171784 151836 171836 151842
rect 171784 151778 171836 151784
rect 170588 139460 170640 139466
rect 170588 139402 170640 139408
rect 170496 138032 170548 138038
rect 170496 137974 170548 137980
rect 170404 123480 170456 123486
rect 170404 123422 170456 123428
rect 169668 116612 169720 116618
rect 169668 116554 169720 116560
rect 169300 116000 169352 116006
rect 169300 115942 169352 115948
rect 169208 111920 169260 111926
rect 169208 111862 169260 111868
rect 169116 111784 169168 111790
rect 169116 111726 169168 111732
rect 169116 109064 169168 109070
rect 169116 109006 169168 109012
rect 169128 82686 169156 109006
rect 169220 89554 169248 111862
rect 169312 93294 169340 115942
rect 170404 106412 170456 106418
rect 170404 106354 170456 106360
rect 169300 93288 169352 93294
rect 169300 93230 169352 93236
rect 169208 89548 169260 89554
rect 169208 89490 169260 89496
rect 169116 82680 169168 82686
rect 169116 82622 169168 82628
rect 169024 82544 169076 82550
rect 169024 82486 169076 82492
rect 170416 81326 170444 106354
rect 170508 89418 170536 137974
rect 170600 93430 170628 139402
rect 170680 124228 170732 124234
rect 170680 124170 170732 124176
rect 170588 93424 170640 93430
rect 170588 93366 170640 93372
rect 170692 90846 170720 124170
rect 171796 92138 171824 151778
rect 173348 150476 173400 150482
rect 173348 150418 173400 150424
rect 171876 146328 171928 146334
rect 171876 146270 171928 146276
rect 171888 94178 171916 146270
rect 173164 133952 173216 133958
rect 173164 133894 173216 133900
rect 171968 128376 172020 128382
rect 171968 128318 172020 128324
rect 171876 94172 171928 94178
rect 171876 94114 171928 94120
rect 171784 92132 171836 92138
rect 171784 92074 171836 92080
rect 170680 90840 170732 90846
rect 170680 90782 170732 90788
rect 170496 89412 170548 89418
rect 170496 89354 170548 89360
rect 170404 81320 170456 81326
rect 170404 81262 170456 81268
rect 166448 79960 166500 79966
rect 166448 79902 166500 79908
rect 171980 79830 172008 128318
rect 172060 114572 172112 114578
rect 172060 114514 172112 114520
rect 172072 88194 172100 114514
rect 172060 88188 172112 88194
rect 172060 88130 172112 88136
rect 171968 79824 172020 79830
rect 171968 79766 172020 79772
rect 173176 78470 173204 133894
rect 173256 122936 173308 122942
rect 173256 122878 173308 122884
rect 173268 85202 173296 122878
rect 173360 113694 173388 150418
rect 173440 120148 173492 120154
rect 173440 120090 173492 120096
rect 173348 113688 173400 113694
rect 173348 113630 173400 113636
rect 173452 93362 173480 120090
rect 173440 93356 173492 93362
rect 173440 93298 173492 93304
rect 173256 85196 173308 85202
rect 173256 85138 173308 85144
rect 173164 78464 173216 78470
rect 173164 78406 173216 78412
rect 133144 77240 133196 77246
rect 115846 77208 115902 77217
rect 133144 77182 133196 77188
rect 115846 77143 115902 77152
rect 118700 76628 118752 76634
rect 118700 76570 118752 76576
rect 106924 75880 106976 75886
rect 106924 75822 106976 75828
rect 99104 75812 99156 75818
rect 99104 75754 99156 75760
rect 67640 75268 67692 75274
rect 67640 75210 67692 75216
rect 64696 75200 64748 75206
rect 64696 75142 64748 75148
rect 64604 73840 64656 73846
rect 64604 73782 64656 73788
rect 64420 71052 64472 71058
rect 64420 70994 64472 71000
rect 64880 65544 64932 65550
rect 64880 65486 64932 65492
rect 64892 16574 64920 65486
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 53380 3596 53432 3602
rect 53380 3538 53432 3544
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3538
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 59636 6248 59688 6254
rect 59636 6190 59688 6196
rect 59648 480 59676 6190
rect 60844 480 60872 16546
rect 63224 13184 63276 13190
rect 63224 13126 63276 13132
rect 62028 4820 62080 4826
rect 62028 4762 62080 4768
rect 62040 480 62068 4762
rect 63236 480 63264 13126
rect 64340 480 64368 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 7608 66772 7614
rect 66720 7550 66772 7556
rect 66732 480 66760 7550
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 75210
rect 80060 72480 80112 72486
rect 80060 72422 80112 72428
rect 74540 71120 74592 71126
rect 74540 71062 74592 71068
rect 69020 64184 69072 64190
rect 69020 64126 69072 64132
rect 69032 16574 69060 64126
rect 71780 29708 71832 29714
rect 71780 29650 71832 29656
rect 70398 24168 70454 24177
rect 70398 24103 70454 24112
rect 70412 16574 70440 24103
rect 71792 16574 71820 29650
rect 74552 16574 74580 71062
rect 77300 69692 77352 69698
rect 77300 69634 77352 69640
rect 75920 62824 75972 62830
rect 75920 62766 75972 62772
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 69124 480 69152 16546
rect 69848 15904 69900 15910
rect 69848 15846 69900 15852
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 15846
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 73804 6180 73856 6186
rect 73804 6122 73856 6128
rect 73816 480 73844 6122
rect 75012 480 75040 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 62766
rect 77312 3602 77340 69634
rect 78680 61396 78732 61402
rect 78680 61338 78732 61344
rect 77392 17332 77444 17338
rect 77392 17274 77444 17280
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77404 480 77432 17274
rect 78692 16574 78720 61338
rect 80072 16574 80100 72422
rect 81440 68400 81492 68406
rect 81440 68342 81492 68348
rect 81452 16574 81480 68342
rect 85580 66972 85632 66978
rect 85580 66914 85632 66920
rect 82820 60104 82872 60110
rect 82820 60046 82872 60052
rect 82832 16574 82860 60046
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3538
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 85592 6914 85620 66914
rect 88340 65612 88392 65618
rect 88340 65554 88392 65560
rect 85672 58744 85724 58750
rect 85672 58686 85724 58692
rect 85684 16574 85712 58686
rect 86960 46232 87012 46238
rect 86960 46174 87012 46180
rect 86972 16574 87000 46174
rect 88352 16574 88380 65554
rect 92478 64152 92534 64161
rect 92478 64087 92534 64096
rect 89720 57316 89772 57322
rect 89720 57258 89772 57264
rect 89732 16574 89760 57258
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 85592 6886 85712 6914
rect 84476 2100 84528 2106
rect 84476 2042 84528 2048
rect 84488 480 84516 2042
rect 85684 480 85712 6886
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 10396 91612 10402
rect 91560 10338 91612 10344
rect 91572 480 91600 10338
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 64087
rect 96620 55956 96672 55962
rect 96620 55898 96672 55904
rect 93860 33856 93912 33862
rect 93860 33798 93912 33804
rect 93872 16574 93900 33798
rect 96632 16574 96660 55898
rect 100760 54596 100812 54602
rect 100760 54538 100812 54544
rect 98642 43480 98698 43489
rect 98642 43415 98698 43424
rect 98000 19984 98052 19990
rect 98000 19926 98052 19932
rect 98012 16574 98040 19926
rect 93872 16546 93992 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 93964 480 93992 16546
rect 95148 9036 95200 9042
rect 95148 8978 95200 8984
rect 95160 480 95188 8978
rect 96252 4888 96304 4894
rect 96252 4830 96304 4836
rect 96264 480 96292 4830
rect 97460 480 97488 16546
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 98656 3534 98684 43415
rect 99840 3596 99892 3602
rect 99840 3538 99892 3544
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99852 480 99880 3538
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 54538
rect 103520 53168 103572 53174
rect 103520 53110 103572 53116
rect 102140 22908 102192 22914
rect 102140 22850 102192 22856
rect 102152 3534 102180 22850
rect 103532 16574 103560 53110
rect 107660 51740 107712 51746
rect 107660 51682 107712 51688
rect 106280 50448 106332 50454
rect 106280 50390 106332 50396
rect 104900 18692 104952 18698
rect 104900 18634 104952 18640
rect 104912 16574 104940 18634
rect 106292 16574 106320 50390
rect 107672 16574 107700 51682
rect 110420 47660 110472 47666
rect 110420 47602 110472 47608
rect 109040 32496 109092 32502
rect 109040 32438 109092 32444
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102232 14544 102284 14550
rect 102232 14486 102284 14492
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 102244 480 102272 14486
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 32438
rect 110432 3602 110460 47602
rect 113180 44940 113232 44946
rect 113180 44882 113232 44888
rect 110512 26988 110564 26994
rect 110512 26930 110564 26936
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 110524 480 110552 26930
rect 113192 16574 113220 44882
rect 114560 31068 114612 31074
rect 114560 31010 114612 31016
rect 114572 16574 114600 31010
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 112812 7676 112864 7682
rect 112812 7618 112864 7624
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111628 480 111656 3538
rect 112824 480 112852 7618
rect 114020 480 114048 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 117318 11656 117374 11665
rect 117318 11591 117374 11600
rect 116400 2168 116452 2174
rect 116400 2110 116452 2116
rect 116412 480 116440 2110
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 11591
rect 118712 3602 118740 76570
rect 124220 73908 124272 73914
rect 124220 73850 124272 73856
rect 118792 49088 118844 49094
rect 118792 49030 118844 49036
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 118804 480 118832 49030
rect 122840 46300 122892 46306
rect 122840 46242 122892 46248
rect 120080 25560 120132 25566
rect 120080 25502 120132 25508
rect 120092 16574 120120 25502
rect 122852 16574 122880 46242
rect 124232 16574 124260 73850
rect 120092 16546 120672 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 119908 480 119936 3538
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122288 15972 122340 15978
rect 122288 15914 122340 15920
rect 122300 480 122328 15914
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 132960 9104 133012 9110
rect 132960 9046 133012 9052
rect 129372 6316 129424 6322
rect 129372 6258 129424 6264
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 125888 480 125916 3538
rect 129384 480 129412 6258
rect 132972 480 133000 9046
rect 136456 7744 136508 7750
rect 136456 7686 136508 7692
rect 136468 480 136496 7686
rect 173912 3602 173940 271866
rect 174636 144220 174688 144226
rect 174636 144162 174688 144168
rect 174544 129804 174596 129810
rect 174544 129746 174596 129752
rect 174556 82618 174584 129746
rect 174648 109002 174676 144162
rect 176016 140888 176068 140894
rect 176016 140830 176068 140836
rect 175924 131164 175976 131170
rect 175924 131106 175976 131112
rect 174820 113212 174872 113218
rect 174820 113154 174872 113160
rect 174636 108996 174688 109002
rect 174636 108938 174688 108944
rect 174728 107704 174780 107710
rect 174728 107646 174780 107652
rect 174544 82612 174596 82618
rect 174544 82554 174596 82560
rect 174740 79898 174768 107646
rect 174832 94042 174860 113154
rect 174820 94036 174872 94042
rect 174820 93978 174872 93984
rect 175936 81258 175964 131106
rect 176028 92274 176056 140830
rect 177316 119406 177344 391954
rect 188344 387864 188396 387870
rect 188344 387806 188396 387812
rect 180064 336796 180116 336802
rect 180064 336738 180116 336744
rect 178776 298376 178828 298382
rect 178776 298318 178828 298324
rect 178682 294128 178738 294137
rect 178682 294063 178738 294072
rect 177396 235272 177448 235278
rect 177396 235214 177448 235220
rect 177304 119400 177356 119406
rect 177304 119342 177356 119348
rect 176108 104916 176160 104922
rect 176108 104858 176160 104864
rect 176016 92268 176068 92274
rect 176016 92210 176068 92216
rect 176120 86902 176148 104858
rect 176108 86896 176160 86902
rect 176108 86838 176160 86844
rect 175924 81252 175976 81258
rect 175924 81194 175976 81200
rect 174728 79892 174780 79898
rect 174728 79834 174780 79840
rect 177408 46918 177436 235214
rect 177488 134020 177540 134026
rect 177488 133962 177540 133968
rect 177500 85338 177528 133962
rect 177580 121508 177632 121514
rect 177580 121450 177632 121456
rect 177592 88058 177620 121450
rect 177672 118856 177724 118862
rect 177672 118798 177724 118804
rect 177684 89486 177712 118798
rect 178696 95169 178724 294063
rect 178788 178906 178816 298318
rect 178776 178900 178828 178906
rect 178776 178842 178828 178848
rect 178776 120216 178828 120222
rect 178776 120158 178828 120164
rect 178682 95160 178738 95169
rect 178682 95095 178738 95104
rect 177672 89480 177724 89486
rect 177672 89422 177724 89428
rect 177580 88052 177632 88058
rect 177580 87994 177632 88000
rect 177488 85332 177540 85338
rect 177488 85274 177540 85280
rect 178788 84046 178816 120158
rect 178868 110492 178920 110498
rect 178868 110434 178920 110440
rect 178776 84040 178828 84046
rect 178776 83982 178828 83988
rect 178880 75818 178908 110434
rect 178960 107772 179012 107778
rect 178960 107714 179012 107720
rect 178972 93906 179000 107714
rect 178960 93900 179012 93906
rect 178960 93842 179012 93848
rect 180076 80714 180104 336738
rect 186964 305720 187016 305726
rect 186964 305662 187016 305668
rect 180156 301096 180208 301102
rect 180156 301038 180208 301044
rect 180168 183054 180196 301038
rect 182824 296880 182876 296886
rect 182824 296822 182876 296828
rect 185582 296848 185638 296857
rect 181444 295588 181496 295594
rect 181444 295530 181496 295536
rect 180248 191344 180300 191350
rect 180248 191286 180300 191292
rect 180156 183048 180208 183054
rect 180156 182990 180208 182996
rect 180260 90982 180288 191286
rect 181456 177313 181484 295530
rect 182836 180198 182864 296822
rect 185582 296783 185638 296792
rect 184204 238128 184256 238134
rect 184204 238070 184256 238076
rect 182824 180192 182876 180198
rect 182824 180134 182876 180140
rect 181442 177304 181498 177313
rect 181442 177239 181498 177248
rect 182824 143608 182876 143614
rect 182824 143550 182876 143556
rect 181444 138712 181496 138718
rect 181444 138654 181496 138660
rect 180340 125724 180392 125730
rect 180340 125666 180392 125672
rect 180248 90976 180300 90982
rect 180248 90918 180300 90924
rect 180352 83978 180380 125666
rect 181456 92342 181484 138654
rect 181536 116068 181588 116074
rect 181536 116010 181588 116016
rect 181444 92336 181496 92342
rect 181444 92278 181496 92284
rect 181548 90710 181576 116010
rect 181536 90704 181588 90710
rect 181536 90646 181588 90652
rect 182836 87990 182864 143550
rect 184216 95198 184244 238070
rect 184296 187740 184348 187746
rect 184296 187682 184348 187688
rect 184308 160002 184336 187682
rect 184296 159996 184348 160002
rect 184296 159938 184348 159944
rect 184296 142180 184348 142186
rect 184296 142122 184348 142128
rect 184204 95192 184256 95198
rect 184204 95134 184256 95140
rect 182824 87984 182876 87990
rect 182824 87926 182876 87932
rect 180340 83972 180392 83978
rect 180340 83914 180392 83920
rect 180156 83496 180208 83502
rect 180156 83438 180208 83444
rect 180064 80708 180116 80714
rect 180064 80650 180116 80656
rect 178868 75812 178920 75818
rect 178868 75754 178920 75760
rect 177396 46912 177448 46918
rect 177396 46854 177448 46860
rect 173900 3596 173952 3602
rect 173900 3538 173952 3544
rect 180168 3466 180196 83438
rect 184308 81122 184336 142122
rect 184388 121576 184440 121582
rect 184388 121518 184440 121524
rect 184400 86834 184428 121518
rect 185596 95033 185624 296783
rect 185676 135312 185728 135318
rect 185676 135254 185728 135260
rect 185582 95024 185638 95033
rect 185582 94959 185638 94968
rect 184388 86828 184440 86834
rect 184388 86770 184440 86776
rect 184296 81116 184348 81122
rect 184296 81058 184348 81064
rect 185688 79762 185716 135254
rect 185676 79756 185728 79762
rect 185676 79698 185728 79704
rect 180156 3460 180208 3466
rect 180156 3402 180208 3408
rect 186976 2242 187004 305662
rect 187056 229832 187108 229838
rect 187056 229774 187108 229780
rect 187068 33114 187096 229774
rect 187148 147688 187200 147694
rect 187148 147630 187200 147636
rect 187160 89350 187188 147630
rect 188356 91798 188384 387806
rect 206284 381540 206336 381546
rect 206284 381482 206336 381488
rect 202144 374672 202196 374678
rect 202144 374614 202196 374620
rect 198004 359508 198056 359514
rect 198004 359450 198056 359456
rect 191104 347132 191156 347138
rect 191104 347074 191156 347080
rect 189722 181384 189778 181393
rect 189722 181319 189778 181328
rect 188436 176724 188488 176730
rect 188436 176666 188488 176672
rect 188448 161430 188476 176666
rect 188436 161424 188488 161430
rect 188436 161366 188488 161372
rect 188528 113280 188580 113286
rect 188528 113222 188580 113228
rect 188436 109132 188488 109138
rect 188436 109074 188488 109080
rect 188344 91792 188396 91798
rect 188344 91734 188396 91740
rect 187148 89344 187200 89350
rect 187148 89286 187200 89292
rect 188448 78674 188476 109074
rect 188540 84114 188568 113222
rect 189736 96422 189764 181319
rect 189816 144968 189868 144974
rect 189816 144910 189868 144916
rect 189724 96416 189776 96422
rect 189724 96358 189776 96364
rect 189828 85270 189856 144910
rect 189816 85264 189868 85270
rect 189816 85206 189868 85212
rect 188528 84108 188580 84114
rect 188528 84050 188580 84056
rect 188436 78668 188488 78674
rect 188436 78610 188488 78616
rect 187056 33108 187108 33114
rect 187056 33050 187108 33056
rect 191116 7750 191144 347074
rect 196624 337476 196676 337482
rect 196624 337418 196676 337424
rect 195244 301572 195296 301578
rect 195244 301514 195296 301520
rect 192484 277500 192536 277506
rect 192484 277442 192536 277448
rect 192496 188494 192524 277442
rect 192484 188488 192536 188494
rect 192484 188430 192536 188436
rect 193862 177440 193918 177449
rect 193862 177375 193918 177384
rect 192576 136672 192628 136678
rect 192576 136614 192628 136620
rect 191196 131232 191248 131238
rect 191196 131174 191248 131180
rect 191208 92410 191236 131174
rect 192484 127016 192536 127022
rect 192484 126958 192536 126964
rect 191288 110560 191340 110566
rect 191288 110502 191340 110508
rect 191196 92404 191248 92410
rect 191196 92346 191248 92352
rect 191300 78538 191328 110502
rect 191288 78532 191340 78538
rect 191288 78474 191340 78480
rect 192496 75886 192524 126958
rect 192588 93974 192616 136614
rect 192576 93968 192628 93974
rect 192576 93910 192628 93916
rect 192484 75880 192536 75886
rect 192484 75822 192536 75828
rect 191104 7744 191156 7750
rect 191104 7686 191156 7692
rect 193876 5030 193904 177375
rect 193864 5024 193916 5030
rect 193864 4966 193916 4972
rect 195256 3466 195284 301514
rect 195428 142248 195480 142254
rect 195428 142190 195480 142196
rect 195336 119400 195388 119406
rect 195336 119342 195388 119348
rect 195348 20058 195376 119342
rect 195440 89622 195468 142190
rect 195428 89616 195480 89622
rect 195428 89558 195480 89564
rect 195336 20052 195388 20058
rect 195336 19994 195388 20000
rect 196636 17406 196664 337418
rect 196716 194132 196768 194138
rect 196716 194074 196768 194080
rect 196728 93537 196756 194074
rect 196808 153332 196860 153338
rect 196808 153274 196860 153280
rect 196714 93528 196770 93537
rect 196714 93463 196770 93472
rect 196716 89004 196768 89010
rect 196716 88946 196768 88952
rect 196624 17400 196676 17406
rect 196624 17342 196676 17348
rect 196728 3534 196756 88946
rect 196820 86766 196848 153274
rect 196808 86760 196860 86766
rect 196808 86702 196860 86708
rect 198016 13258 198044 359450
rect 198188 299600 198240 299606
rect 198188 299542 198240 299548
rect 198096 183116 198148 183122
rect 198096 183058 198148 183064
rect 198004 13252 198056 13258
rect 198004 13194 198056 13200
rect 198108 9178 198136 183058
rect 198200 181694 198228 299542
rect 199384 295656 199436 295662
rect 199384 295598 199436 295604
rect 198188 181688 198240 181694
rect 198188 181630 198240 181636
rect 199396 95130 199424 295598
rect 199476 180328 199528 180334
rect 199476 180270 199528 180276
rect 199384 95124 199436 95130
rect 199384 95066 199436 95072
rect 199488 11830 199516 180270
rect 200764 124296 200816 124302
rect 200764 124238 200816 124244
rect 200776 88262 200804 124238
rect 200856 100768 200908 100774
rect 200856 100710 200908 100716
rect 200764 88256 200816 88262
rect 200764 88198 200816 88204
rect 200868 77246 200896 100710
rect 200856 77240 200908 77246
rect 200856 77182 200908 77188
rect 202156 14618 202184 374614
rect 204904 351280 204956 351286
rect 204904 351222 204956 351228
rect 203524 301028 203576 301034
rect 203524 300970 203576 300976
rect 202236 296812 202288 296818
rect 202236 296754 202288 296760
rect 202248 175953 202276 296754
rect 203536 178974 203564 300970
rect 203524 178968 203576 178974
rect 203524 178910 203576 178916
rect 202234 175944 202290 175953
rect 202234 175879 202290 175888
rect 203616 135380 203668 135386
rect 203616 135322 203668 135328
rect 202236 123480 202288 123486
rect 202236 123422 202288 123428
rect 202144 14612 202196 14618
rect 202144 14554 202196 14560
rect 199476 11824 199528 11830
rect 199476 11766 199528 11772
rect 198096 9172 198148 9178
rect 198096 9114 198148 9120
rect 202248 3602 202276 123422
rect 203524 116612 203576 116618
rect 203524 116554 203576 116560
rect 203536 9110 203564 116554
rect 203628 92478 203656 135322
rect 203616 92472 203668 92478
rect 203616 92414 203668 92420
rect 204916 16046 204944 351222
rect 204996 278860 205048 278866
rect 204996 278802 205048 278808
rect 205008 180334 205036 278802
rect 204996 180328 205048 180334
rect 204996 180270 205048 180276
rect 204994 119368 205050 119377
rect 204994 119303 205050 119312
rect 204904 16040 204956 16046
rect 204904 15982 204956 15988
rect 203524 9104 203576 9110
rect 203524 9046 203576 9052
rect 205008 6390 205036 119303
rect 204996 6384 205048 6390
rect 204996 6326 205048 6332
rect 206296 6322 206324 381482
rect 209044 312588 209096 312594
rect 209044 312530 209096 312536
rect 207664 259480 207716 259486
rect 207664 259422 207716 259428
rect 206468 249824 206520 249830
rect 206468 249766 206520 249772
rect 206376 180260 206428 180266
rect 206376 180202 206428 180208
rect 206388 18766 206416 180202
rect 206480 177449 206508 249766
rect 207676 180266 207704 259422
rect 207664 180260 207716 180266
rect 207664 180202 207716 180208
rect 206466 177440 206522 177449
rect 206466 177375 206522 177384
rect 207664 117360 207716 117366
rect 207664 117302 207716 117308
rect 206468 103556 206520 103562
rect 206468 103498 206520 103504
rect 206480 93673 206508 103498
rect 206466 93664 206522 93673
rect 206466 93599 206522 93608
rect 207676 81394 207704 117302
rect 207664 81388 207716 81394
rect 207664 81330 207716 81336
rect 206376 18760 206428 18766
rect 206376 18702 206428 18708
rect 206284 6316 206336 6322
rect 206284 6258 206336 6264
rect 209056 3670 209084 312530
rect 213184 307148 213236 307154
rect 213184 307090 213236 307096
rect 211804 274712 211856 274718
rect 211804 274654 211856 274660
rect 210424 273284 210476 273290
rect 210424 273226 210476 273232
rect 209136 241596 209188 241602
rect 209136 241538 209188 241544
rect 209148 96626 209176 241538
rect 210436 176186 210464 273226
rect 211816 179042 211844 274654
rect 211804 179036 211856 179042
rect 211804 178978 211856 178984
rect 210516 178152 210568 178158
rect 210516 178094 210568 178100
rect 210424 176180 210476 176186
rect 210424 176122 210476 176128
rect 210528 150414 210556 178094
rect 211804 176112 211856 176118
rect 211804 176054 211856 176060
rect 210608 176044 210660 176050
rect 210608 175986 210660 175992
rect 210620 168298 210648 175986
rect 211816 169658 211844 176054
rect 211804 169652 211856 169658
rect 211804 169594 211856 169600
rect 210608 168292 210660 168298
rect 210608 168234 210660 168240
rect 211804 152448 211856 152454
rect 211804 152390 211856 152396
rect 210516 150408 210568 150414
rect 210516 150350 210568 150356
rect 209228 118788 209280 118794
rect 209228 118730 209280 118736
rect 209136 96620 209188 96626
rect 209136 96562 209188 96568
rect 209240 80034 209268 118730
rect 210424 117428 210476 117434
rect 210424 117370 210476 117376
rect 210436 82822 210464 117370
rect 210608 104984 210660 104990
rect 210608 104926 210660 104932
rect 210516 100836 210568 100842
rect 210516 100778 210568 100784
rect 210528 89690 210556 100778
rect 210620 94897 210648 104926
rect 210606 94888 210662 94897
rect 210606 94823 210662 94832
rect 210516 89684 210568 89690
rect 210516 89626 210568 89632
rect 211816 88126 211844 152390
rect 211896 102196 211948 102202
rect 211896 102138 211948 102144
rect 211908 89729 211936 102138
rect 211894 89720 211950 89729
rect 211894 89655 211950 89664
rect 211804 88120 211856 88126
rect 211804 88062 211856 88068
rect 210424 82816 210476 82822
rect 210424 82758 210476 82764
rect 209228 80028 209280 80034
rect 209228 79970 209280 79976
rect 213196 4962 213224 307090
rect 213276 270564 213328 270570
rect 213276 270506 213328 270512
rect 213288 181762 213316 270506
rect 213368 207800 213420 207806
rect 213368 207742 213420 207748
rect 213276 181756 213328 181762
rect 213276 181698 213328 181704
rect 213380 180402 213408 207742
rect 213460 184952 213512 184958
rect 213460 184894 213512 184900
rect 213368 180396 213420 180402
rect 213368 180338 213420 180344
rect 213276 175976 213328 175982
rect 213276 175918 213328 175924
rect 213288 166161 213316 175918
rect 213274 166152 213330 166161
rect 213274 166087 213330 166096
rect 213472 164801 213500 184894
rect 214576 178702 214604 394674
rect 215944 387116 215996 387122
rect 215944 387058 215996 387064
rect 214656 284368 214708 284374
rect 214656 284310 214708 284316
rect 214668 189786 214696 284310
rect 214656 189780 214708 189786
rect 214656 189722 214708 189728
rect 214748 189100 214800 189106
rect 214748 189042 214800 189048
rect 214656 186380 214708 186386
rect 214656 186322 214708 186328
rect 214564 178696 214616 178702
rect 214564 178638 214616 178644
rect 214104 178084 214156 178090
rect 214104 178026 214156 178032
rect 213828 176792 213880 176798
rect 213828 176734 213880 176740
rect 213840 175817 213868 176734
rect 213826 175808 213882 175817
rect 213826 175743 213882 175752
rect 214012 175228 214064 175234
rect 214012 175170 214064 175176
rect 213920 175160 213972 175166
rect 213918 175128 213920 175137
rect 213972 175128 213974 175137
rect 213918 175063 213974 175072
rect 214024 174729 214052 175170
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 213918 173768 213974 173777
rect 213918 173703 213974 173712
rect 214116 173369 214144 178026
rect 214564 176248 214616 176254
rect 214564 176190 214616 176196
rect 214102 173360 214158 173369
rect 214102 173295 214158 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172417 213960 172450
rect 214012 172440 214064 172446
rect 213918 172408 213974 172417
rect 214012 172382 214064 172388
rect 213918 172343 213974 172352
rect 214024 172009 214052 172382
rect 214010 172000 214066 172009
rect 214010 171935 214066 171944
rect 214012 171080 214064 171086
rect 214012 171022 214064 171028
rect 214024 170785 214052 171022
rect 214010 170776 214066 170785
rect 214010 170711 214066 170720
rect 213920 169720 213972 169726
rect 213920 169662 213972 169668
rect 214010 169688 214066 169697
rect 213932 169425 213960 169662
rect 214010 169623 214012 169632
rect 214064 169623 214066 169632
rect 214012 169594 214064 169600
rect 213918 169416 213974 169425
rect 213918 169351 213974 169360
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 214024 168065 214052 168234
rect 214010 168056 214066 168065
rect 214010 167991 214066 168000
rect 213918 166968 213974 166977
rect 213918 166903 213920 166912
rect 213972 166903 213974 166912
rect 213920 166874 213972 166880
rect 214012 166864 214064 166870
rect 214012 166806 214064 166812
rect 214024 166705 214052 166806
rect 214010 166696 214066 166705
rect 214010 166631 214066 166640
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 213458 164792 213514 164801
rect 213458 164727 213514 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163985 213960 164154
rect 213918 163976 213974 163985
rect 213918 163911 213974 163920
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214576 160857 214604 176190
rect 214668 161474 214696 186322
rect 214760 171134 214788 189042
rect 215114 171184 215170 171193
rect 214760 171106 215064 171134
rect 215114 171119 215170 171128
rect 214668 161446 214972 161474
rect 214562 160848 214618 160857
rect 214562 160783 214618 160792
rect 214104 160744 214156 160750
rect 214104 160686 214156 160692
rect 213920 160064 213972 160070
rect 213918 160032 213920 160041
rect 213972 160032 213974 160041
rect 213918 159967 213974 159976
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 214024 159497 214052 159938
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 214116 158681 214144 160686
rect 214102 158672 214158 158681
rect 214944 158658 214972 161446
rect 214102 158607 214158 158616
rect 214852 158630 214972 158658
rect 214012 157344 214064 157350
rect 213918 157312 213974 157321
rect 214012 157286 214064 157292
rect 213918 157247 213920 157256
rect 213972 157247 213974 157256
rect 213920 157218 213972 157224
rect 214024 156913 214052 157286
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 214852 155961 214880 158630
rect 215036 158137 215064 171106
rect 215128 171018 215156 171119
rect 215116 171012 215168 171018
rect 215116 170954 215168 170960
rect 215022 158128 215078 158137
rect 215022 158063 215078 158072
rect 214932 158024 214984 158030
rect 214932 157966 214984 157972
rect 214838 155952 214894 155961
rect 213920 155916 213972 155922
rect 214838 155887 214894 155896
rect 213920 155858 213972 155864
rect 213932 155553 213960 155858
rect 213918 155544 213974 155553
rect 213918 155479 213974 155488
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153368 213974 153377
rect 213918 153303 213920 153312
rect 213972 153303 213974 153312
rect 213920 153274 213972 153280
rect 214024 153270 214052 153847
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 213918 152688 213974 152697
rect 213918 152623 213974 152632
rect 213932 152454 213960 152623
rect 213920 152448 213972 152454
rect 213920 152390 213972 152396
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151842 213960 151943
rect 214654 151872 214710 151881
rect 213920 151836 213972 151842
rect 214654 151807 214710 151816
rect 213920 151778 213972 151784
rect 213918 150920 213974 150929
rect 213918 150855 213974 150864
rect 213932 150482 213960 150855
rect 214470 150784 214526 150793
rect 214470 150719 214526 150728
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 214024 150249 214052 150350
rect 214010 150240 214066 150249
rect 214010 150175 214066 150184
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 213918 146367 213974 146376
rect 213932 146334 213960 146367
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213920 144968 213972 144974
rect 213918 144936 213920 144945
rect 213972 144936 213974 144945
rect 213918 144871 213974 144880
rect 213918 143984 213974 143993
rect 213918 143919 213974 143928
rect 213932 143614 213960 143919
rect 213920 143608 213972 143614
rect 213274 143576 213330 143585
rect 213920 143550 213972 143556
rect 213274 143511 213330 143520
rect 213288 78606 213316 143511
rect 214024 142866 214052 146639
rect 214012 142860 214064 142866
rect 214012 142802 214064 142808
rect 214010 142760 214066 142769
rect 214010 142695 214066 142704
rect 213918 142352 213974 142361
rect 213918 142287 213974 142296
rect 213932 142254 213960 142287
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 142695
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 213918 140992 213974 141001
rect 213918 140927 213974 140936
rect 213932 140894 213960 140927
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141335
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 214484 140078 214512 150719
rect 214668 144226 214696 151807
rect 214944 149569 214972 157966
rect 214930 149560 214986 149569
rect 214930 149495 214986 149504
rect 214656 144220 214708 144226
rect 214656 144162 214708 144168
rect 214472 140072 214524 140078
rect 213918 140040 213974 140049
rect 214472 140014 214524 140020
rect 213918 139975 213974 139984
rect 213932 139466 213960 139975
rect 214010 139496 214066 139505
rect 213920 139460 213972 139466
rect 214010 139431 214066 139440
rect 213920 139402 213972 139408
rect 213918 138816 213974 138825
rect 213918 138751 213974 138760
rect 213932 138038 213960 138751
rect 214024 138718 214052 139431
rect 214012 138712 214064 138718
rect 214012 138654 214064 138660
rect 214654 138136 214710 138145
rect 214654 138071 214710 138080
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 137456 213974 137465
rect 213918 137391 213974 137400
rect 213932 136678 213960 137391
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 135688 214066 135697
rect 214010 135623 214066 135632
rect 213918 135416 213974 135425
rect 214024 135386 214052 135623
rect 213918 135351 213974 135360
rect 214012 135380 214064 135386
rect 213932 135318 213960 135351
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 214010 134328 214066 134337
rect 214010 134263 214066 134272
rect 213918 134056 213974 134065
rect 214024 134026 214052 134263
rect 213918 133991 213974 134000
rect 214012 134020 214064 134026
rect 213932 133958 213960 133991
rect 214012 133962 214064 133968
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214562 132560 214618 132569
rect 214562 132495 214618 132504
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 214024 131238 214052 131407
rect 214012 131232 214064 131238
rect 213918 131200 213974 131209
rect 214012 131174 214064 131180
rect 213918 131135 213920 131144
rect 213972 131135 213974 131144
rect 213920 131106 213972 131112
rect 213918 130112 213974 130121
rect 213918 130047 213974 130056
rect 213932 129810 213960 130047
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 213918 128480 213974 128489
rect 213918 128415 213974 128424
rect 213932 128382 213960 128415
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 127528 213974 127537
rect 213918 127463 213974 127472
rect 213932 127022 213960 127463
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 214024 125730 214052 126103
rect 213918 125695 213974 125704
rect 214012 125724 214064 125730
rect 213932 125662 213960 125695
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 214024 122942 214052 123519
rect 214012 122936 214064 122942
rect 213918 122904 213974 122913
rect 214012 122878 214064 122884
rect 213918 122839 213920 122848
rect 213972 122839 213974 122848
rect 213920 122810 213972 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 214024 121582 214052 122159
rect 214012 121576 214064 121582
rect 213918 121544 213974 121553
rect 214012 121518 214064 121524
rect 213918 121479 213920 121488
rect 213972 121479 213974 121488
rect 213920 121450 213972 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 214024 120222 214052 120799
rect 214012 120216 214064 120222
rect 213918 120184 213974 120193
rect 214012 120158 214064 120164
rect 213918 120119 213920 120128
rect 213972 120119 213974 120128
rect 213920 120090 213972 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213366 119096 213422 119105
rect 213366 119031 213422 119040
rect 213380 82754 213408 119031
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118862 213960 118895
rect 213920 118856 213972 118862
rect 213920 118798 213972 118804
rect 214024 118794 214052 119575
rect 214012 118788 214064 118794
rect 214012 118730 214064 118736
rect 213918 117600 213974 117609
rect 213918 117535 213974 117544
rect 213932 117366 213960 117535
rect 214012 117428 214064 117434
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 214024 117337 214052 117370
rect 213920 117302 213972 117308
rect 214010 117328 214066 117337
rect 214010 117263 214066 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 214024 116074 214052 116175
rect 214012 116068 214064 116074
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213918 115968 213920 115977
rect 213972 115968 213974 115977
rect 213918 115903 213974 115912
rect 213918 115016 213974 115025
rect 213918 114951 213974 114960
rect 213458 114608 213514 114617
rect 213932 114578 213960 114951
rect 213458 114543 213514 114552
rect 213920 114572 213972 114578
rect 213472 86970 213500 114543
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 213920 113280 213972 113286
rect 213918 113248 213920 113257
rect 213972 113248 213974 113257
rect 214024 113218 214052 113591
rect 213918 113183 213974 113192
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 214024 111926 214052 112231
rect 214012 111920 214064 111926
rect 213918 111888 213974 111897
rect 214012 111862 214064 111868
rect 213918 111823 213920 111832
rect 213972 111823 213974 111832
rect 213920 111794 213972 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 214024 110566 214052 110871
rect 214012 110560 214064 110566
rect 213918 110528 213974 110537
rect 214012 110502 214064 110508
rect 213918 110463 213920 110472
rect 213972 110463 213974 110472
rect 213920 110434 213972 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109168 213974 109177
rect 213918 109103 213920 109112
rect 213972 109103 213974 109112
rect 213920 109074 213972 109080
rect 214024 109070 214052 109647
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 214024 107778 214052 108287
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106584 213974 106593
rect 213918 106519 213974 106528
rect 213932 106350 213960 106519
rect 214024 106418 214052 106927
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 213918 105768 213974 105777
rect 213918 105703 213974 105712
rect 213932 104922 213960 105703
rect 214010 105224 214066 105233
rect 214010 105159 214066 105168
rect 214024 104990 214052 105159
rect 214012 104984 214064 104990
rect 214012 104926 214064 104932
rect 213920 104916 213972 104922
rect 213920 104858 213972 104864
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102504 213974 102513
rect 213918 102439 213974 102448
rect 213932 102202 213960 102439
rect 213920 102196 213972 102202
rect 213920 102138 213972 102144
rect 214010 101144 214066 101153
rect 214010 101079 214066 101088
rect 213918 100872 213974 100881
rect 214024 100842 214052 101079
rect 213918 100807 213974 100816
rect 214012 100836 214064 100842
rect 213932 100774 213960 100807
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 213918 99784 213974 99793
rect 213918 99719 213974 99728
rect 213932 99414 213960 99719
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 214024 98122 214052 98359
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 214576 93158 214604 132495
rect 214668 132494 214696 138071
rect 214668 132466 214788 132494
rect 214760 118017 214788 132466
rect 214746 118008 214802 118017
rect 214746 117943 214802 117952
rect 214654 103864 214710 103873
rect 214654 103799 214710 103808
rect 214564 93152 214616 93158
rect 214564 93094 214616 93100
rect 214668 91050 214696 103799
rect 214838 99512 214894 99521
rect 214838 99447 214894 99456
rect 214746 96656 214802 96665
rect 214746 96591 214802 96600
rect 214656 91044 214708 91050
rect 214656 90986 214708 90992
rect 213460 86964 213512 86970
rect 213460 86906 213512 86912
rect 214760 85474 214788 96591
rect 214852 90914 214880 99447
rect 214840 90908 214892 90914
rect 214840 90850 214892 90856
rect 214748 85468 214800 85474
rect 214748 85410 214800 85416
rect 213368 82748 213420 82754
rect 213368 82690 213420 82696
rect 213276 78600 213328 78606
rect 213276 78542 213328 78548
rect 213184 4956 213236 4962
rect 213184 4898 213236 4904
rect 209044 3664 209096 3670
rect 209044 3606 209096 3612
rect 202236 3596 202288 3602
rect 202236 3538 202288 3544
rect 215956 3534 215984 387058
rect 217232 345704 217284 345710
rect 217232 345646 217284 345652
rect 216036 313948 216088 313954
rect 216036 313890 216088 313896
rect 216048 3738 216076 313890
rect 216128 265056 216180 265062
rect 216128 264998 216180 265004
rect 216140 95062 216168 264998
rect 216218 97064 216274 97073
rect 216218 96999 216274 97008
rect 216128 95056 216180 95062
rect 216128 94998 216180 95004
rect 216232 85542 216260 96999
rect 216678 95840 216734 95849
rect 216678 95775 216734 95784
rect 216220 85536 216272 85542
rect 216220 85478 216272 85484
rect 216692 84182 216720 95775
rect 217244 93158 217272 345646
rect 218704 247104 218756 247110
rect 218704 247046 218756 247052
rect 218716 176118 218744 247046
rect 218796 199708 218848 199714
rect 218796 199650 218848 199656
rect 218808 177410 218836 199650
rect 220096 178770 220124 397530
rect 238022 392592 238078 392601
rect 238022 392527 238078 392536
rect 222936 372632 222988 372638
rect 222936 372574 222988 372580
rect 222844 302456 222896 302462
rect 222844 302398 222896 302404
rect 221464 281648 221516 281654
rect 221464 281590 221516 281596
rect 220176 205012 220228 205018
rect 220176 204954 220228 204960
rect 220084 178764 220136 178770
rect 220084 178706 220136 178712
rect 220188 177478 220216 204954
rect 221476 177546 221504 281590
rect 222856 178022 222884 302398
rect 222948 282198 222976 372574
rect 233884 355360 233936 355366
rect 233884 355302 233936 355308
rect 226984 307828 227036 307834
rect 226984 307770 227036 307776
rect 224224 299532 224276 299538
rect 224224 299474 224276 299480
rect 222936 282192 222988 282198
rect 222936 282134 222988 282140
rect 222844 178016 222896 178022
rect 222844 177958 222896 177964
rect 221464 177540 221516 177546
rect 221464 177482 221516 177488
rect 220176 177472 220228 177478
rect 220176 177414 220228 177420
rect 218796 177404 218848 177410
rect 218796 177346 218848 177352
rect 218704 176112 218756 176118
rect 218704 176054 218756 176060
rect 224236 175982 224264 299474
rect 225604 296744 225656 296750
rect 225604 296686 225656 296692
rect 224316 287088 224368 287094
rect 224316 287030 224368 287036
rect 224328 187066 224356 287030
rect 224316 187060 224368 187066
rect 224316 187002 224368 187008
rect 225616 176050 225644 296686
rect 226996 180470 227024 307770
rect 231124 302388 231176 302394
rect 231124 302330 231176 302336
rect 227076 298308 227128 298314
rect 227076 298250 227128 298256
rect 226984 180464 227036 180470
rect 226984 180406 227036 180412
rect 227088 177585 227116 298250
rect 227168 281580 227220 281586
rect 227168 281522 227220 281528
rect 227074 177576 227130 177585
rect 227074 177511 227130 177520
rect 227180 177342 227208 281522
rect 230480 236768 230532 236774
rect 230480 236710 230532 236716
rect 227720 183048 227772 183054
rect 227720 182990 227772 182996
rect 227168 177336 227220 177342
rect 227168 177278 227220 177284
rect 225604 176044 225656 176050
rect 225604 175986 225656 175992
rect 224224 175976 224276 175982
rect 224224 175918 224276 175924
rect 227732 175817 227760 182990
rect 229376 178016 229428 178022
rect 229376 177958 229428 177964
rect 229100 177540 229152 177546
rect 229100 177482 229152 177488
rect 227718 175808 227774 175817
rect 227718 175743 227774 175752
rect 229112 174729 229140 177482
rect 229192 176180 229244 176186
rect 229192 176122 229244 176128
rect 229098 174720 229154 174729
rect 229098 174655 229154 174664
rect 229204 172417 229232 176122
rect 229284 176112 229336 176118
rect 229284 176054 229336 176060
rect 229190 172408 229246 172417
rect 229190 172343 229246 172352
rect 229296 171465 229324 176054
rect 229282 171456 229338 171465
rect 229282 171391 229338 171400
rect 229388 168609 229416 177958
rect 229744 170468 229796 170474
rect 229744 170410 229796 170416
rect 229374 168600 229430 168609
rect 229374 168535 229430 168544
rect 229756 142089 229784 170410
rect 229836 170400 229888 170406
rect 229836 170342 229888 170348
rect 229848 151065 229876 170342
rect 230492 157729 230520 236710
rect 231136 216102 231164 302330
rect 233240 263628 233292 263634
rect 233240 263570 233292 263576
rect 231860 251864 231912 251870
rect 231860 251806 231912 251812
rect 231124 216096 231176 216102
rect 231124 216038 231176 216044
rect 230572 206372 230624 206378
rect 230572 206314 230624 206320
rect 230584 158681 230612 206314
rect 230664 196784 230716 196790
rect 230664 196726 230716 196732
rect 230676 171134 230704 196726
rect 231768 173868 231820 173874
rect 231768 173810 231820 173816
rect 231124 173800 231176 173806
rect 231780 173777 231808 173810
rect 231124 173742 231176 173748
rect 231766 173768 231822 173777
rect 231136 173369 231164 173742
rect 231492 173732 231544 173738
rect 231766 173703 231822 173712
rect 231492 173674 231544 173680
rect 231122 173360 231178 173369
rect 231122 173295 231178 173304
rect 231504 172825 231532 173674
rect 231490 172816 231546 172825
rect 231490 172751 231546 172760
rect 231768 172508 231820 172514
rect 231768 172450 231820 172456
rect 231780 171873 231808 172450
rect 231766 171864 231822 171873
rect 231766 171799 231822 171808
rect 230676 171106 230980 171134
rect 230756 169584 230808 169590
rect 230754 169552 230756 169561
rect 230808 169552 230810 169561
rect 230754 169487 230810 169496
rect 230570 158672 230626 158681
rect 230570 158607 230626 158616
rect 230478 157720 230534 157729
rect 230478 157655 230534 157664
rect 230952 156233 230980 171106
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231124 171012 231176 171018
rect 231124 170954 231176 170960
rect 231136 170513 231164 170954
rect 231492 170944 231544 170950
rect 231780 170921 231808 171022
rect 231492 170886 231544 170892
rect 231766 170912 231822 170921
rect 231122 170504 231178 170513
rect 231122 170439 231178 170448
rect 231504 169969 231532 170886
rect 231766 170847 231822 170856
rect 231490 169960 231546 169969
rect 231490 169895 231546 169904
rect 231492 169720 231544 169726
rect 231492 169662 231544 169668
rect 231504 169017 231532 169662
rect 231490 169008 231546 169017
rect 231490 168943 231546 168952
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231780 168065 231808 168302
rect 231766 168056 231822 168065
rect 231766 167991 231822 168000
rect 231766 167104 231822 167113
rect 231872 167090 231900 251806
rect 232044 241528 232096 241534
rect 232044 241470 232096 241476
rect 231952 227044 232004 227050
rect 231952 226986 232004 226992
rect 231822 167062 231900 167090
rect 231766 167039 231822 167048
rect 231676 167000 231728 167006
rect 231676 166942 231728 166948
rect 231688 166161 231716 166942
rect 231768 166932 231820 166938
rect 231768 166874 231820 166880
rect 231674 166152 231730 166161
rect 231674 166087 231730 166096
rect 231780 165753 231808 166874
rect 231766 165744 231822 165753
rect 231766 165679 231822 165688
rect 231124 165572 231176 165578
rect 231124 165514 231176 165520
rect 231136 164393 231164 165514
rect 231676 165504 231728 165510
rect 231676 165446 231728 165452
rect 231688 164801 231716 165446
rect 231768 165436 231820 165442
rect 231768 165378 231820 165384
rect 231780 165209 231808 165378
rect 231766 165200 231822 165209
rect 231766 165135 231822 165144
rect 231674 164792 231730 164801
rect 231674 164727 231730 164736
rect 231122 164384 231178 164393
rect 231122 164319 231178 164328
rect 231124 164212 231176 164218
rect 231124 164154 231176 164160
rect 231136 162897 231164 164154
rect 231768 164144 231820 164150
rect 231768 164086 231820 164092
rect 231676 164076 231728 164082
rect 231676 164018 231728 164024
rect 231688 163441 231716 164018
rect 231780 163849 231808 164086
rect 231766 163840 231822 163849
rect 231766 163775 231822 163784
rect 231674 163432 231730 163441
rect 231674 163367 231730 163376
rect 231122 162888 231178 162897
rect 231032 162852 231084 162858
rect 231122 162823 231178 162832
rect 231032 162794 231084 162800
rect 231044 161537 231072 162794
rect 231676 162716 231728 162722
rect 231676 162658 231728 162664
rect 231688 161945 231716 162658
rect 231768 162512 231820 162518
rect 231766 162480 231768 162489
rect 231820 162480 231822 162489
rect 231766 162415 231822 162424
rect 231674 161936 231730 161945
rect 231674 161871 231730 161880
rect 231030 161528 231086 161537
rect 231030 161463 231086 161472
rect 231676 161424 231728 161430
rect 231676 161366 231728 161372
rect 231688 160585 231716 161366
rect 231768 161356 231820 161362
rect 231768 161298 231820 161304
rect 231780 160993 231808 161298
rect 231766 160984 231822 160993
rect 231766 160919 231822 160928
rect 231674 160576 231730 160585
rect 231674 160511 231730 160520
rect 231768 160064 231820 160070
rect 231766 160032 231768 160041
rect 231820 160032 231822 160041
rect 231676 159996 231728 160002
rect 231766 159967 231822 159976
rect 231676 159938 231728 159944
rect 231688 159633 231716 159938
rect 231674 159624 231730 159633
rect 231674 159559 231730 159568
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 231688 159089 231716 159462
rect 231674 159080 231730 159089
rect 231674 159015 231730 159024
rect 231490 158808 231546 158817
rect 231490 158743 231546 158752
rect 230938 156224 230994 156233
rect 230938 156159 230994 156168
rect 230940 155916 230992 155922
rect 230940 155858 230992 155864
rect 230572 155848 230624 155854
rect 230570 155816 230572 155825
rect 230624 155816 230626 155825
rect 230570 155751 230626 155760
rect 230952 155281 230980 155858
rect 230938 155272 230994 155281
rect 230938 155207 230994 155216
rect 231400 154556 231452 154562
rect 231400 154498 231452 154504
rect 231124 154148 231176 154154
rect 231124 154090 231176 154096
rect 230756 153196 230808 153202
rect 230756 153138 230808 153144
rect 230768 152969 230796 153138
rect 230754 152960 230810 152969
rect 230754 152895 230810 152904
rect 229834 151056 229890 151065
rect 229834 150991 229890 151000
rect 230940 150408 230992 150414
rect 230940 150350 230992 150356
rect 230952 150113 230980 150350
rect 231032 150340 231084 150346
rect 231032 150282 231084 150288
rect 230938 150104 230994 150113
rect 230938 150039 230994 150048
rect 231044 149705 231072 150282
rect 231030 149696 231086 149705
rect 231030 149631 231086 149640
rect 230940 147620 230992 147626
rect 230940 147562 230992 147568
rect 230756 147552 230808 147558
rect 230756 147494 230808 147500
rect 230768 147257 230796 147494
rect 230754 147248 230810 147257
rect 230754 147183 230810 147192
rect 230952 146849 230980 147562
rect 230938 146840 230994 146849
rect 230938 146775 230994 146784
rect 230756 144220 230808 144226
rect 230756 144162 230808 144168
rect 230768 143993 230796 144162
rect 230754 143984 230810 143993
rect 230754 143919 230810 143928
rect 230480 143472 230532 143478
rect 230480 143414 230532 143420
rect 230492 142497 230520 143414
rect 230478 142488 230534 142497
rect 230478 142423 230534 142432
rect 229742 142080 229798 142089
rect 229742 142015 229798 142024
rect 230940 140616 230992 140622
rect 230940 140558 230992 140564
rect 230952 140185 230980 140558
rect 230938 140176 230994 140185
rect 230938 140111 230994 140120
rect 230020 139460 230072 139466
rect 230020 139402 230072 139408
rect 229928 136672 229980 136678
rect 229928 136614 229980 136620
rect 229744 135312 229796 135318
rect 229744 135254 229796 135260
rect 229098 96656 229154 96665
rect 229098 96591 229100 96600
rect 229152 96591 229154 96600
rect 229100 96562 229152 96568
rect 228364 95260 228416 95266
rect 228364 95202 228416 95208
rect 222844 94512 222896 94518
rect 222844 94454 222896 94460
rect 217232 93152 217284 93158
rect 217232 93094 217284 93100
rect 216680 84176 216732 84182
rect 216680 84118 216732 84124
rect 222856 18698 222884 94454
rect 228376 76566 228404 95202
rect 228364 76560 228416 76566
rect 228364 76502 228416 76508
rect 222844 18692 222896 18698
rect 222844 18634 222896 18640
rect 229756 4894 229784 135254
rect 229836 113212 229888 113218
rect 229836 113154 229888 113160
rect 229848 13122 229876 113154
rect 229940 50454 229968 136614
rect 230032 73914 230060 139402
rect 231032 138712 231084 138718
rect 231032 138654 231084 138660
rect 230756 134224 230808 134230
rect 230756 134166 230808 134172
rect 230768 134065 230796 134166
rect 230754 134056 230810 134065
rect 230754 133991 230810 134000
rect 231044 132569 231072 138654
rect 231030 132560 231086 132569
rect 231030 132495 231086 132504
rect 230756 132456 230808 132462
rect 230756 132398 230808 132404
rect 230768 132161 230796 132398
rect 230754 132152 230810 132161
rect 230754 132087 230810 132096
rect 230756 128308 230808 128314
rect 230756 128250 230808 128256
rect 230768 127945 230796 128250
rect 230754 127936 230810 127945
rect 230754 127871 230810 127880
rect 230664 124908 230716 124914
rect 230664 124850 230716 124856
rect 230676 118969 230704 124850
rect 230940 122800 230992 122806
rect 230940 122742 230992 122748
rect 230952 122233 230980 122742
rect 230938 122224 230994 122233
rect 230938 122159 230994 122168
rect 230662 118960 230718 118969
rect 230662 118895 230718 118904
rect 231136 117473 231164 154090
rect 231412 153921 231440 154498
rect 231398 153912 231454 153921
rect 231398 153847 231454 153856
rect 231308 153400 231360 153406
rect 231306 153368 231308 153377
rect 231360 153368 231362 153377
rect 231306 153303 231362 153312
rect 231216 149796 231268 149802
rect 231216 149738 231268 149744
rect 231122 117464 231178 117473
rect 231122 117399 231178 117408
rect 230664 117292 230716 117298
rect 230664 117234 230716 117240
rect 230676 117065 230704 117234
rect 231124 117156 231176 117162
rect 231124 117098 231176 117104
rect 230662 117056 230718 117065
rect 230662 116991 230718 117000
rect 230572 115252 230624 115258
rect 230572 115194 230624 115200
rect 230584 107953 230612 115194
rect 231136 114617 231164 117098
rect 231228 116113 231256 149738
rect 231308 149524 231360 149530
rect 231308 149466 231360 149472
rect 231320 149161 231348 149466
rect 231306 149152 231362 149161
rect 231306 149087 231362 149096
rect 231400 147008 231452 147014
rect 231400 146950 231452 146956
rect 231412 135425 231440 146950
rect 231504 146305 231532 158743
rect 231676 157344 231728 157350
rect 231676 157286 231728 157292
rect 231688 156777 231716 157286
rect 231768 157276 231820 157282
rect 231768 157218 231820 157224
rect 231780 157185 231808 157218
rect 231766 157176 231822 157185
rect 231766 157111 231822 157120
rect 231674 156768 231730 156777
rect 231674 156703 231730 156712
rect 231768 154352 231820 154358
rect 231766 154320 231768 154329
rect 231820 154320 231822 154329
rect 231766 154255 231822 154264
rect 231768 153128 231820 153134
rect 231768 153070 231820 153076
rect 231676 152720 231728 152726
rect 231676 152662 231728 152668
rect 231688 152561 231716 152662
rect 231674 152552 231730 152561
rect 231674 152487 231730 152496
rect 231780 152017 231808 153070
rect 231766 152008 231822 152017
rect 231766 151943 231822 151952
rect 231964 151814 231992 226986
rect 232056 166705 232084 241470
rect 232136 206440 232188 206446
rect 232136 206382 232188 206388
rect 232042 166696 232098 166705
rect 232042 166631 232098 166640
rect 232148 155854 232176 206382
rect 232504 167680 232556 167686
rect 232504 167622 232556 167628
rect 232136 155848 232188 155854
rect 232136 155790 232188 155796
rect 231872 151786 231992 151814
rect 231676 151768 231728 151774
rect 231676 151710 231728 151716
rect 231688 150657 231716 151710
rect 231768 151700 231820 151706
rect 231768 151642 231820 151648
rect 231780 151609 231808 151642
rect 231766 151600 231822 151609
rect 231766 151535 231822 151544
rect 231674 150648 231730 150657
rect 231674 150583 231730 150592
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148209 231808 148990
rect 231766 148200 231822 148209
rect 231766 148135 231822 148144
rect 231490 146296 231546 146305
rect 231490 146231 231546 146240
rect 231768 146260 231820 146266
rect 231768 146202 231820 146208
rect 231676 146192 231728 146198
rect 231676 146134 231728 146140
rect 231688 145353 231716 146134
rect 231780 145897 231808 146202
rect 231766 145888 231822 145897
rect 231766 145823 231822 145832
rect 231674 145344 231730 145353
rect 231674 145279 231730 145288
rect 231872 145058 231900 151786
rect 232516 147558 232544 167622
rect 233252 164218 233280 263570
rect 233896 257378 233924 355302
rect 234620 295452 234672 295458
rect 234620 295394 234672 295400
rect 233884 257372 233936 257378
rect 233884 257314 233936 257320
rect 233332 211812 233384 211818
rect 233332 211754 233384 211760
rect 233240 164212 233292 164218
rect 233240 164154 233292 164160
rect 233344 162858 233372 211754
rect 233424 209092 233476 209098
rect 233424 209034 233476 209040
rect 233436 165578 233464 209034
rect 233516 195424 233568 195430
rect 233516 195366 233568 195372
rect 233424 165572 233476 165578
rect 233424 165514 233476 165520
rect 233332 162852 233384 162858
rect 233332 162794 233384 162800
rect 232780 156188 232832 156194
rect 232780 156130 232832 156136
rect 232686 153232 232742 153241
rect 232686 153167 232742 153176
rect 232504 147552 232556 147558
rect 232504 147494 232556 147500
rect 231688 145030 231900 145058
rect 231688 144945 231716 145030
rect 231674 144936 231730 144945
rect 231674 144871 231730 144880
rect 231768 144900 231820 144906
rect 231768 144842 231820 144848
rect 231780 144401 231808 144842
rect 231766 144392 231822 144401
rect 231766 144327 231822 144336
rect 232700 144226 232728 153167
rect 232688 144220 232740 144226
rect 232688 144162 232740 144168
rect 232596 144152 232648 144158
rect 232596 144094 232648 144100
rect 231768 143540 231820 143546
rect 231768 143482 231820 143488
rect 231780 143449 231808 143482
rect 231766 143440 231822 143449
rect 231766 143375 231822 143384
rect 231492 140752 231544 140758
rect 231492 140694 231544 140700
rect 231766 140720 231822 140729
rect 231504 139777 231532 140694
rect 231766 140655 231768 140664
rect 231820 140655 231822 140664
rect 231768 140626 231820 140632
rect 231490 139768 231546 139777
rect 231490 139703 231546 139712
rect 231768 139392 231820 139398
rect 231768 139334 231820 139340
rect 231676 139256 231728 139262
rect 231674 139224 231676 139233
rect 231728 139224 231730 139233
rect 231674 139159 231730 139168
rect 231780 138825 231808 139334
rect 231766 138816 231822 138825
rect 231766 138751 231822 138760
rect 231492 137964 231544 137970
rect 231492 137906 231544 137912
rect 231504 136921 231532 137906
rect 231768 137896 231820 137902
rect 231768 137838 231820 137844
rect 231780 137329 231808 137838
rect 231766 137320 231822 137329
rect 231766 137255 231822 137264
rect 231490 136912 231546 136921
rect 231490 136847 231546 136856
rect 231768 136604 231820 136610
rect 231768 136546 231820 136552
rect 231676 136536 231728 136542
rect 231676 136478 231728 136484
rect 231688 135969 231716 136478
rect 231780 136377 231808 136546
rect 231766 136368 231822 136377
rect 231766 136303 231822 136312
rect 231674 135960 231730 135969
rect 231674 135895 231730 135904
rect 231582 135824 231638 135833
rect 231582 135759 231638 135768
rect 231398 135416 231454 135425
rect 231398 135351 231454 135360
rect 231306 133784 231362 133793
rect 231306 133719 231362 133728
rect 231320 125361 231348 133719
rect 231492 132388 231544 132394
rect 231492 132330 231544 132336
rect 231504 131617 231532 132330
rect 231490 131608 231546 131617
rect 231490 131543 231546 131552
rect 231400 131028 231452 131034
rect 231400 130970 231452 130976
rect 231412 129849 231440 130970
rect 231492 130960 231544 130966
rect 231492 130902 231544 130908
rect 231504 130257 231532 130902
rect 231490 130248 231546 130257
rect 231490 130183 231546 130192
rect 231398 129840 231454 129849
rect 231398 129775 231454 129784
rect 231596 126993 231624 135759
rect 231768 135244 231820 135250
rect 231768 135186 231820 135192
rect 231676 135176 231728 135182
rect 231676 135118 231728 135124
rect 231688 134473 231716 135118
rect 231780 135017 231808 135186
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231768 133884 231820 133890
rect 231768 133826 231820 133832
rect 231676 133816 231728 133822
rect 231676 133758 231728 133764
rect 231688 133113 231716 133758
rect 231780 133521 231808 133826
rect 231766 133512 231822 133521
rect 231766 133447 231822 133456
rect 231674 133104 231730 133113
rect 231674 133039 231730 133048
rect 231768 132320 231820 132326
rect 231768 132262 231820 132268
rect 231780 131209 231808 132262
rect 231766 131200 231822 131209
rect 231766 131135 231822 131144
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231676 129668 231728 129674
rect 231676 129610 231728 129616
rect 231688 128897 231716 129610
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231674 128888 231730 128897
rect 231674 128823 231730 128832
rect 231766 128344 231822 128353
rect 231766 128279 231822 128288
rect 231780 128246 231808 128279
rect 231768 128240 231820 128246
rect 231768 128182 231820 128188
rect 231676 128172 231728 128178
rect 231676 128114 231728 128120
rect 231688 127401 231716 128114
rect 231674 127392 231730 127401
rect 231674 127327 231730 127336
rect 231582 126984 231638 126993
rect 231582 126919 231638 126928
rect 231768 126948 231820 126954
rect 231768 126890 231820 126896
rect 231780 126449 231808 126890
rect 231766 126440 231822 126449
rect 231766 126375 231822 126384
rect 231584 125860 231636 125866
rect 231584 125802 231636 125808
rect 231492 125588 231544 125594
rect 231492 125530 231544 125536
rect 231306 125352 231362 125361
rect 231306 125287 231362 125296
rect 231504 124545 231532 125530
rect 231490 124536 231546 124545
rect 231490 124471 231546 124480
rect 231400 123480 231452 123486
rect 231400 123422 231452 123428
rect 231308 121372 231360 121378
rect 231308 121314 231360 121320
rect 231320 120737 231348 121314
rect 231306 120728 231362 120737
rect 231306 120663 231362 120672
rect 231308 120012 231360 120018
rect 231308 119954 231360 119960
rect 231320 119377 231348 119954
rect 231306 119368 231362 119377
rect 231306 119303 231362 119312
rect 231412 118810 231440 123422
rect 231596 123185 231624 125802
rect 231768 125520 231820 125526
rect 231768 125462 231820 125468
rect 231780 125089 231808 125462
rect 231766 125080 231822 125089
rect 231766 125015 231822 125024
rect 231768 124160 231820 124166
rect 231766 124128 231768 124137
rect 231820 124128 231822 124137
rect 231766 124063 231822 124072
rect 231582 123176 231638 123185
rect 231582 123111 231638 123120
rect 232504 122868 232556 122874
rect 232504 122810 232556 122816
rect 231768 122732 231820 122738
rect 231768 122674 231820 122680
rect 231492 122664 231544 122670
rect 231780 122641 231808 122674
rect 231492 122606 231544 122612
rect 231766 122632 231822 122641
rect 231504 121689 231532 122606
rect 231766 122567 231822 122576
rect 231490 121680 231546 121689
rect 231490 121615 231546 121624
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231492 121304 231544 121310
rect 231780 121281 231808 121382
rect 231492 121246 231544 121252
rect 231766 121272 231822 121281
rect 231504 120329 231532 121246
rect 231766 121207 231822 121216
rect 231490 120320 231546 120329
rect 231490 120255 231546 120264
rect 231768 120080 231820 120086
rect 231768 120022 231820 120028
rect 231780 119785 231808 120022
rect 231766 119776 231822 119785
rect 231766 119711 231822 119720
rect 231320 118782 231440 118810
rect 231214 116104 231270 116113
rect 231214 116039 231270 116048
rect 231216 115524 231268 115530
rect 231216 115466 231268 115472
rect 231228 115161 231256 115466
rect 231214 115152 231270 115161
rect 231214 115087 231270 115096
rect 231122 114608 231178 114617
rect 231122 114543 231178 114552
rect 231320 113665 231348 118782
rect 231400 118652 231452 118658
rect 231400 118594 231452 118600
rect 231412 118017 231440 118594
rect 231398 118008 231454 118017
rect 231398 117943 231454 117952
rect 231400 117836 231452 117842
rect 231400 117778 231452 117784
rect 231306 113656 231362 113665
rect 231306 113591 231362 113600
rect 231124 112464 231176 112470
rect 231124 112406 231176 112412
rect 230940 111172 230992 111178
rect 230940 111114 230992 111120
rect 230952 110809 230980 111114
rect 230938 110800 230994 110809
rect 230938 110735 230994 110744
rect 230570 107944 230626 107953
rect 230570 107879 230626 107888
rect 230756 106684 230808 106690
rect 230756 106626 230808 106632
rect 230768 106593 230796 106626
rect 230754 106584 230810 106593
rect 230754 106519 230810 106528
rect 230572 104848 230624 104854
rect 230572 104790 230624 104796
rect 230584 104281 230612 104790
rect 230570 104272 230626 104281
rect 230570 104207 230626 104216
rect 230480 104168 230532 104174
rect 230480 104110 230532 104116
rect 230492 102785 230520 104110
rect 231136 103329 231164 112406
rect 231412 104689 231440 117778
rect 231492 117224 231544 117230
rect 231492 117166 231544 117172
rect 231504 116521 231532 117166
rect 231490 116512 231546 116521
rect 231490 116447 231546 116456
rect 231768 114504 231820 114510
rect 231768 114446 231820 114452
rect 231492 114436 231544 114442
rect 231492 114378 231544 114384
rect 231504 113257 231532 114378
rect 231780 114209 231808 114446
rect 231766 114200 231822 114209
rect 231766 114135 231822 114144
rect 231490 113248 231546 113257
rect 231490 113183 231546 113192
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231676 112872 231728 112878
rect 231676 112814 231728 112820
rect 231688 112713 231716 112814
rect 231674 112704 231730 112713
rect 231674 112639 231730 112648
rect 231780 112305 231808 113086
rect 231766 112296 231822 112305
rect 231766 112231 231822 112240
rect 231768 111784 231820 111790
rect 231674 111752 231730 111761
rect 231768 111726 231820 111732
rect 231674 111687 231676 111696
rect 231728 111687 231730 111696
rect 231676 111658 231728 111664
rect 231780 111353 231808 111726
rect 231766 111344 231822 111353
rect 231766 111279 231822 111288
rect 231676 110424 231728 110430
rect 231676 110366 231728 110372
rect 231766 110392 231822 110401
rect 231688 109857 231716 110366
rect 231766 110327 231768 110336
rect 231820 110327 231822 110336
rect 231768 110298 231820 110304
rect 231674 109848 231730 109857
rect 231674 109783 231730 109792
rect 231676 109744 231728 109750
rect 231676 109686 231728 109692
rect 231688 109449 231716 109686
rect 231674 109440 231730 109449
rect 231674 109375 231730 109384
rect 231676 108996 231728 109002
rect 231676 108938 231728 108944
rect 231688 108497 231716 108938
rect 231768 108928 231820 108934
rect 231766 108896 231768 108905
rect 231820 108896 231822 108905
rect 231766 108831 231822 108840
rect 231674 108488 231730 108497
rect 231584 108452 231636 108458
rect 231674 108423 231730 108432
rect 231584 108394 231636 108400
rect 231492 107160 231544 107166
rect 231490 107128 231492 107137
rect 231544 107128 231546 107137
rect 231490 107063 231546 107072
rect 231492 106276 231544 106282
rect 231492 106218 231544 106224
rect 231504 105233 231532 106218
rect 231490 105224 231546 105233
rect 231490 105159 231546 105168
rect 231398 104680 231454 104689
rect 231398 104615 231454 104624
rect 231596 103737 231624 108394
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231780 107545 231808 107578
rect 231766 107536 231822 107545
rect 231766 107471 231822 107480
rect 231768 106208 231820 106214
rect 231768 106150 231820 106156
rect 231780 105641 231808 106150
rect 231766 105632 231822 105641
rect 231766 105567 231822 105576
rect 231582 103728 231638 103737
rect 231582 103663 231638 103672
rect 231122 103320 231178 103329
rect 231122 103255 231178 103264
rect 231584 102808 231636 102814
rect 230478 102776 230534 102785
rect 231584 102750 231636 102756
rect 230478 102711 230534 102720
rect 230940 102196 230992 102202
rect 230940 102138 230992 102144
rect 230572 102128 230624 102134
rect 230572 102070 230624 102076
rect 230584 100881 230612 102070
rect 230756 101992 230808 101998
rect 230756 101934 230808 101940
rect 230768 101425 230796 101934
rect 230754 101416 230810 101425
rect 230754 101351 230810 101360
rect 230570 100872 230626 100881
rect 230570 100807 230626 100816
rect 230952 98025 230980 102138
rect 231492 100700 231544 100706
rect 231492 100642 231544 100648
rect 231504 99929 231532 100642
rect 231490 99920 231546 99929
rect 231490 99855 231546 99864
rect 231492 98660 231544 98666
rect 231492 98602 231544 98608
rect 231504 98569 231532 98602
rect 231490 98560 231546 98569
rect 231490 98495 231546 98504
rect 230938 98016 230994 98025
rect 230938 97951 230994 97960
rect 231596 97617 231624 102750
rect 231676 101448 231728 101454
rect 231676 101390 231728 101396
rect 231688 100473 231716 101390
rect 231768 100632 231820 100638
rect 231768 100574 231820 100580
rect 231674 100464 231730 100473
rect 231674 100399 231730 100408
rect 231780 99521 231808 100574
rect 231766 99512 231822 99521
rect 231766 99447 231822 99456
rect 231768 99340 231820 99346
rect 231768 99282 231820 99288
rect 231780 99113 231808 99282
rect 231766 99104 231822 99113
rect 231766 99039 231822 99048
rect 231582 97608 231638 97617
rect 231582 97543 231638 97552
rect 231766 97064 231822 97073
rect 231766 96999 231822 97008
rect 231124 96688 231176 96694
rect 231124 96630 231176 96636
rect 230572 96620 230624 96626
rect 230572 96562 230624 96568
rect 230478 95704 230534 95713
rect 230478 95639 230534 95648
rect 230492 92546 230520 95639
rect 230584 93906 230612 96562
rect 230572 93900 230624 93906
rect 230572 93842 230624 93848
rect 230480 92540 230532 92546
rect 230480 92482 230532 92488
rect 230584 84194 230612 93842
rect 230492 84166 230612 84194
rect 230020 73908 230072 73914
rect 230020 73850 230072 73856
rect 229928 50448 229980 50454
rect 229928 50390 229980 50396
rect 230492 22778 230520 84166
rect 230480 22772 230532 22778
rect 230480 22714 230532 22720
rect 229836 13116 229888 13122
rect 229836 13058 229888 13064
rect 231136 8974 231164 96630
rect 231780 95946 231808 96999
rect 231768 95940 231820 95946
rect 231768 95882 231820 95888
rect 232516 14550 232544 122810
rect 232608 104854 232636 144094
rect 232792 143478 232820 156130
rect 233528 155922 233556 195366
rect 234068 163056 234120 163062
rect 234068 162998 234120 163004
rect 233884 162172 233936 162178
rect 233884 162114 233936 162120
rect 233516 155916 233568 155922
rect 233516 155858 233568 155864
rect 233896 153406 233924 162114
rect 233976 154624 234028 154630
rect 233976 154566 234028 154572
rect 233884 153400 233936 153406
rect 233884 153342 233936 153348
rect 233884 147688 233936 147694
rect 233884 147630 233936 147636
rect 232780 143472 232832 143478
rect 232780 143414 232832 143420
rect 232688 142860 232740 142866
rect 232688 142802 232740 142808
rect 232596 104848 232648 104854
rect 232596 104790 232648 104796
rect 232596 102264 232648 102270
rect 232596 102206 232648 102212
rect 232608 35290 232636 102206
rect 232700 101998 232728 142802
rect 232780 140820 232832 140826
rect 232780 140762 232832 140768
rect 232792 102202 232820 140762
rect 233896 107166 233924 147630
rect 233988 117162 234016 154566
rect 234080 125866 234108 162998
rect 234632 152726 234660 295394
rect 234712 289876 234764 289882
rect 234712 289818 234764 289824
rect 234724 159526 234752 289818
rect 237380 269204 237432 269210
rect 237380 269146 237432 269152
rect 236000 253972 236052 253978
rect 236000 253914 236052 253920
rect 234804 202224 234856 202230
rect 234804 202166 234856 202172
rect 234712 159520 234764 159526
rect 234712 159462 234764 159468
rect 234620 152720 234672 152726
rect 234620 152662 234672 152668
rect 234816 147626 234844 202166
rect 234896 199572 234948 199578
rect 234896 199514 234948 199520
rect 234908 150346 234936 199514
rect 235448 151972 235500 151978
rect 235448 151914 235500 151920
rect 234896 150340 234948 150346
rect 234896 150282 234948 150288
rect 234804 147620 234856 147626
rect 234804 147562 234856 147568
rect 234160 144968 234212 144974
rect 234160 144910 234212 144916
rect 234068 125860 234120 125866
rect 234068 125802 234120 125808
rect 233976 117156 234028 117162
rect 233976 117098 234028 117104
rect 234068 116000 234120 116006
rect 234068 115942 234120 115948
rect 233884 107160 233936 107166
rect 233884 107102 233936 107108
rect 233976 103556 234028 103562
rect 233976 103498 234028 103504
rect 232780 102196 232832 102202
rect 232780 102138 232832 102144
rect 232688 101992 232740 101998
rect 232688 101934 232740 101940
rect 233884 92540 233936 92546
rect 233884 92482 233936 92488
rect 232596 35284 232648 35290
rect 232596 35226 232648 35232
rect 232504 14544 232556 14550
rect 232504 14486 232556 14492
rect 231124 8968 231176 8974
rect 231124 8910 231176 8916
rect 229744 4888 229796 4894
rect 229744 4830 229796 4836
rect 216036 3732 216088 3738
rect 216036 3674 216088 3680
rect 196716 3528 196768 3534
rect 196716 3470 196768 3476
rect 215944 3528 215996 3534
rect 215944 3470 215996 3476
rect 195244 3460 195296 3466
rect 195244 3402 195296 3408
rect 233896 3398 233924 92482
rect 233988 32434 234016 103498
rect 234080 55894 234108 115942
rect 234172 108458 234200 144910
rect 235356 128376 235408 128382
rect 235356 128318 235408 128324
rect 235264 117360 235316 117366
rect 235264 117302 235316 117308
rect 234160 108452 234212 108458
rect 234160 108394 234212 108400
rect 234160 93900 234212 93906
rect 234160 93842 234212 93848
rect 234172 93770 234200 93842
rect 234160 93764 234212 93770
rect 234160 93706 234212 93712
rect 234068 55888 234120 55894
rect 234068 55830 234120 55836
rect 233976 32428 234028 32434
rect 233976 32370 234028 32376
rect 235276 6254 235304 117302
rect 235368 42158 235396 128318
rect 235460 111178 235488 151914
rect 236012 149530 236040 253914
rect 236092 194064 236144 194070
rect 236092 194006 236144 194012
rect 236000 149524 236052 149530
rect 236000 149466 236052 149472
rect 235540 147756 235592 147762
rect 235540 147698 235592 147704
rect 235448 111172 235500 111178
rect 235448 111114 235500 111120
rect 235552 106690 235580 147698
rect 235632 146328 235684 146334
rect 235632 146270 235684 146276
rect 235644 117842 235672 146270
rect 236104 139262 236132 194006
rect 236184 181620 236236 181626
rect 236184 181562 236236 181568
rect 236196 154358 236224 181562
rect 237392 175234 237420 269146
rect 237472 245676 237524 245682
rect 237472 245618 237524 245624
rect 236644 175228 236696 175234
rect 236644 175170 236696 175176
rect 237380 175228 237432 175234
rect 237380 175170 237432 175176
rect 236656 162518 236684 175170
rect 236644 162512 236696 162518
rect 236644 162454 236696 162460
rect 237380 157412 237432 157418
rect 237380 157354 237432 157360
rect 236184 154352 236236 154358
rect 236184 154294 236236 154300
rect 237392 154154 237420 157354
rect 237484 156194 237512 245618
rect 238036 178673 238064 392527
rect 258724 347812 258776 347818
rect 258724 347754 258776 347760
rect 251180 327752 251232 327758
rect 251180 327694 251232 327700
rect 240416 300960 240468 300966
rect 240416 300902 240468 300908
rect 239036 294092 239088 294098
rect 239036 294034 239088 294040
rect 238852 232552 238904 232558
rect 238852 232494 238904 232500
rect 238760 180328 238812 180334
rect 238760 180270 238812 180276
rect 238022 178664 238078 178673
rect 238022 178599 238078 178608
rect 237656 177472 237708 177478
rect 237656 177414 237708 177420
rect 237564 177404 237616 177410
rect 237564 177346 237616 177352
rect 237576 169726 237604 177346
rect 237564 169720 237616 169726
rect 237564 169662 237616 169668
rect 237668 169590 237696 177414
rect 238772 173738 238800 180270
rect 238760 173732 238812 173738
rect 238760 173674 238812 173680
rect 238116 172576 238168 172582
rect 238116 172518 238168 172524
rect 237656 169584 237708 169590
rect 237656 169526 237708 169532
rect 237472 156188 237524 156194
rect 237472 156130 237524 156136
rect 238024 155984 238076 155990
rect 238024 155926 238076 155932
rect 237380 154148 237432 154154
rect 237380 154090 237432 154096
rect 236828 150476 236880 150482
rect 236828 150418 236880 150424
rect 236736 139528 236788 139534
rect 236736 139470 236788 139476
rect 236092 139256 236144 139262
rect 236092 139198 236144 139204
rect 236644 136740 236696 136746
rect 236644 136682 236696 136688
rect 235632 117836 235684 117842
rect 235632 117778 235684 117784
rect 235540 106684 235592 106690
rect 235540 106626 235592 106632
rect 235356 42152 235408 42158
rect 235356 42094 235408 42100
rect 236656 22914 236684 136682
rect 236748 25566 236776 139470
rect 236840 109750 236868 150418
rect 236920 149728 236972 149734
rect 236920 149670 236972 149676
rect 236932 111722 236960 149670
rect 238036 115530 238064 155926
rect 238128 134230 238156 172518
rect 238758 168328 238814 168337
rect 238758 168263 238814 168272
rect 238300 165640 238352 165646
rect 238300 165582 238352 165588
rect 238208 153264 238260 153270
rect 238208 153206 238260 153212
rect 238116 134224 238168 134230
rect 238116 134166 238168 134172
rect 238116 125656 238168 125662
rect 238116 125598 238168 125604
rect 238024 115524 238076 115530
rect 238024 115466 238076 115472
rect 236920 111716 236972 111722
rect 236920 111658 236972 111664
rect 236828 109744 236880 109750
rect 236828 109686 236880 109692
rect 236920 102264 236972 102270
rect 236920 102206 236972 102212
rect 236828 96756 236880 96762
rect 236828 96698 236880 96704
rect 236840 36650 236868 96698
rect 236932 68338 236960 102206
rect 238024 98048 238076 98054
rect 238024 97990 238076 97996
rect 236920 68332 236972 68338
rect 236920 68274 236972 68280
rect 236828 36644 236880 36650
rect 236828 36586 236880 36592
rect 236736 25560 236788 25566
rect 236736 25502 236788 25508
rect 236644 22908 236696 22914
rect 236644 22850 236696 22856
rect 238036 10334 238064 97990
rect 238128 46306 238156 125598
rect 238220 112878 238248 153206
rect 238312 146169 238340 165582
rect 238772 161362 238800 168263
rect 238864 166938 238892 232494
rect 238944 178900 238996 178906
rect 238944 178842 238996 178848
rect 238956 168366 238984 178842
rect 239048 170474 239076 294034
rect 240232 200864 240284 200870
rect 240232 200806 240284 200812
rect 240140 181756 240192 181762
rect 240140 181698 240192 181704
rect 240152 172514 240180 181698
rect 240244 173806 240272 200806
rect 240324 178832 240376 178838
rect 240324 178774 240376 178780
rect 240232 173800 240284 173806
rect 240232 173742 240284 173748
rect 240140 172508 240192 172514
rect 240140 172450 240192 172456
rect 239036 170468 239088 170474
rect 239036 170410 239088 170416
rect 239680 169788 239732 169794
rect 239680 169730 239732 169736
rect 238944 168360 238996 168366
rect 238944 168302 238996 168308
rect 238852 166932 238904 166938
rect 238852 166874 238904 166880
rect 238760 161356 238812 161362
rect 238760 161298 238812 161304
rect 239588 156664 239640 156670
rect 239588 156606 239640 156612
rect 239404 153876 239456 153882
rect 239404 153818 239456 153824
rect 238298 146160 238354 146169
rect 238298 146095 238354 146104
rect 238392 119400 238444 119406
rect 238392 119342 238444 119348
rect 238208 112872 238260 112878
rect 238208 112814 238260 112820
rect 238208 110628 238260 110634
rect 238208 110570 238260 110576
rect 238220 51746 238248 110570
rect 238300 107908 238352 107914
rect 238300 107850 238352 107856
rect 238312 60110 238340 107850
rect 238404 98666 238432 119342
rect 239416 114442 239444 153818
rect 239496 129804 239548 129810
rect 239496 129746 239548 129752
rect 239404 114436 239456 114442
rect 239404 114378 239456 114384
rect 239404 111852 239456 111858
rect 239404 111794 239456 111800
rect 238392 98660 238444 98666
rect 238392 98602 238444 98608
rect 238300 60104 238352 60110
rect 238300 60046 238352 60052
rect 238208 51740 238260 51746
rect 238208 51682 238260 51688
rect 238116 46300 238168 46306
rect 238116 46242 238168 46248
rect 239416 18630 239444 111794
rect 239508 39438 239536 129746
rect 239600 117230 239628 156606
rect 239692 130966 239720 169730
rect 239772 168428 239824 168434
rect 239772 168370 239824 168376
rect 239680 130960 239732 130966
rect 239680 130902 239732 130908
rect 239784 129674 239812 168370
rect 240336 160002 240364 178774
rect 240428 164150 240456 300902
rect 248420 269136 248472 269142
rect 248420 269078 248472 269084
rect 242900 256760 242952 256766
rect 242900 256702 242952 256708
rect 241520 207664 241572 207670
rect 241520 207606 241572 207612
rect 241152 171148 241204 171154
rect 241152 171090 241204 171096
rect 240784 164280 240836 164286
rect 240784 164222 240836 164228
rect 240416 164144 240468 164150
rect 240416 164086 240468 164092
rect 240324 159996 240376 160002
rect 240324 159938 240376 159944
rect 239772 129668 239824 129674
rect 239772 129610 239824 129616
rect 240796 125526 240824 164222
rect 241060 161492 241112 161498
rect 241060 161434 241112 161440
rect 240968 154692 241020 154698
rect 240968 154634 241020 154640
rect 240876 138032 240928 138038
rect 240876 137974 240928 137980
rect 240784 125520 240836 125526
rect 240784 125462 240836 125468
rect 240784 121508 240836 121514
rect 240784 121450 240836 121456
rect 239588 117224 239640 117230
rect 239588 117166 239640 117172
rect 239496 39432 239548 39438
rect 239496 39374 239548 39380
rect 239404 18624 239456 18630
rect 239404 18566 239456 18572
rect 238024 10328 238076 10334
rect 238024 10270 238076 10276
rect 239312 7744 239364 7750
rect 239312 7686 239364 7692
rect 235264 6248 235316 6254
rect 235264 6190 235316 6196
rect 233884 3392 233936 3398
rect 233884 3334 233936 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 186964 2236 187016 2242
rect 186964 2178 187016 2184
rect 235828 480 235856 3334
rect 239324 480 239352 7686
rect 240506 3496 240562 3505
rect 240506 3431 240562 3440
rect 240520 480 240548 3431
rect 240796 2106 240824 121450
rect 240888 44946 240916 137974
rect 240980 114510 241008 154634
rect 241072 122670 241100 161434
rect 241164 138718 241192 171090
rect 241532 167006 241560 207606
rect 241612 188420 241664 188426
rect 241612 188362 241664 188368
rect 241624 170406 241652 188362
rect 241704 180396 241756 180402
rect 241704 180338 241756 180344
rect 241612 170400 241664 170406
rect 241612 170342 241664 170348
rect 241520 167000 241572 167006
rect 241520 166942 241572 166948
rect 241716 165510 241744 180338
rect 242532 173936 242584 173942
rect 242532 173878 242584 173884
rect 242440 168496 242492 168502
rect 242440 168438 242492 168444
rect 241704 165504 241756 165510
rect 241704 165446 241756 165452
rect 242164 163532 242216 163538
rect 242164 163474 242216 163480
rect 241152 138712 241204 138718
rect 241152 138654 241204 138660
rect 242176 124166 242204 163474
rect 242348 160132 242400 160138
rect 242348 160074 242400 160080
rect 242256 146940 242308 146946
rect 242256 146882 242308 146888
rect 242164 124160 242216 124166
rect 242164 124102 242216 124108
rect 241060 122664 241112 122670
rect 241060 122606 241112 122612
rect 240968 114504 241020 114510
rect 240968 114446 241020 114452
rect 240968 106480 241020 106486
rect 240968 106422 241020 106428
rect 240876 44940 240928 44946
rect 240876 44882 240928 44888
rect 240980 29714 241008 106422
rect 242268 106214 242296 146882
rect 242360 121310 242388 160074
rect 242452 131034 242480 168438
rect 242544 147014 242572 173878
rect 242532 147008 242584 147014
rect 242532 146950 242584 146956
rect 242912 143546 242940 256702
rect 244280 222896 244332 222902
rect 244280 222838 244332 222844
rect 242992 192568 243044 192574
rect 242992 192510 243044 192516
rect 243004 173874 243032 192510
rect 243084 178968 243136 178974
rect 243084 178910 243136 178916
rect 242992 173868 243044 173874
rect 242992 173810 243044 173816
rect 243096 167686 243124 178910
rect 243176 176044 243228 176050
rect 243176 175986 243228 175992
rect 243084 167680 243136 167686
rect 243084 167622 243136 167628
rect 243188 165442 243216 175986
rect 243728 173188 243780 173194
rect 243728 173130 243780 173136
rect 243636 167068 243688 167074
rect 243636 167010 243688 167016
rect 243176 165436 243228 165442
rect 243176 165378 243228 165384
rect 242900 143540 242952 143546
rect 242900 143482 242952 143488
rect 243544 135380 243596 135386
rect 243544 135322 243596 135328
rect 242440 131028 242492 131034
rect 242440 130970 242492 130976
rect 242348 121304 242400 121310
rect 242348 121246 242400 121252
rect 242440 120148 242492 120154
rect 242440 120090 242492 120096
rect 242348 113280 242400 113286
rect 242348 113222 242400 113228
rect 242256 106208 242308 106214
rect 242256 106150 242308 106156
rect 242164 104916 242216 104922
rect 242164 104858 242216 104864
rect 240968 29708 241020 29714
rect 240968 29650 241020 29656
rect 241520 17400 241572 17406
rect 241520 17342 241572 17348
rect 241532 16574 241560 17342
rect 241532 16546 241744 16574
rect 240784 2100 240836 2106
rect 240784 2042 240836 2048
rect 241716 480 241744 16546
rect 242176 4826 242204 104858
rect 242256 98116 242308 98122
rect 242256 98058 242308 98064
rect 242268 26926 242296 98058
rect 242360 49026 242388 113222
rect 242452 72486 242480 120090
rect 242440 72480 242492 72486
rect 242440 72422 242492 72428
rect 243556 65618 243584 135322
rect 243648 128178 243676 167010
rect 243740 136542 243768 173130
rect 244292 170950 244320 222838
rect 247040 218748 247092 218754
rect 247040 218690 247092 218696
rect 245660 216096 245712 216102
rect 245660 216038 245712 216044
rect 244372 193996 244424 194002
rect 244372 193938 244424 193944
rect 244280 170944 244332 170950
rect 244280 170886 244332 170892
rect 244384 162722 244412 193938
rect 244556 185768 244608 185774
rect 244556 185710 244608 185716
rect 244464 180192 244516 180198
rect 244464 180134 244516 180140
rect 244372 162716 244424 162722
rect 244372 162658 244424 162664
rect 244476 157282 244504 180134
rect 244568 164082 244596 185710
rect 245672 171086 245700 216038
rect 245844 182912 245896 182918
rect 245844 182854 245896 182860
rect 245752 179036 245804 179042
rect 245752 178978 245804 178984
rect 245660 171080 245712 171086
rect 245660 171022 245712 171028
rect 244924 169856 244976 169862
rect 244924 169798 244976 169804
rect 244556 164076 244608 164082
rect 244556 164018 244608 164024
rect 244464 157276 244516 157282
rect 244464 157218 244516 157224
rect 243820 145036 243872 145042
rect 243820 144978 243872 144984
rect 243728 136536 243780 136542
rect 243728 136478 243780 136484
rect 243636 128172 243688 128178
rect 243636 128114 243688 128120
rect 243636 114572 243688 114578
rect 243636 114514 243688 114520
rect 243544 65612 243596 65618
rect 243544 65554 243596 65560
rect 243648 54534 243676 114514
rect 243832 112470 243860 144978
rect 244936 132326 244964 169798
rect 245016 160200 245068 160206
rect 245016 160142 245068 160148
rect 244924 132320 244976 132326
rect 244924 132262 244976 132268
rect 244924 124228 244976 124234
rect 244924 124170 244976 124176
rect 243820 112464 243872 112470
rect 243820 112406 243872 112412
rect 243728 109064 243780 109070
rect 243728 109006 243780 109012
rect 243636 54528 243688 54534
rect 243636 54470 243688 54476
rect 243740 53174 243768 109006
rect 243728 53168 243780 53174
rect 243728 53110 243780 53116
rect 242348 49020 242400 49026
rect 242348 48962 242400 48968
rect 242256 26920 242308 26926
rect 242256 26862 242308 26868
rect 244936 7682 244964 124170
rect 245028 120018 245056 160142
rect 245108 157480 245160 157486
rect 245108 157422 245160 157428
rect 245016 120012 245068 120018
rect 245016 119954 245068 119960
rect 245120 117298 245148 157422
rect 245764 153134 245792 178978
rect 245856 171018 245884 182854
rect 246396 171216 246448 171222
rect 246396 171158 246448 171164
rect 245844 171012 245896 171018
rect 245844 170954 245896 170960
rect 246304 165708 246356 165714
rect 246304 165650 246356 165656
rect 245752 153128 245804 153134
rect 245752 153070 245804 153076
rect 245200 150544 245252 150550
rect 245200 150486 245252 150492
rect 245108 117292 245160 117298
rect 245108 117234 245160 117240
rect 245016 116068 245068 116074
rect 245016 116010 245068 116016
rect 245028 33794 245056 116010
rect 245212 108934 245240 150486
rect 246316 126954 246344 165650
rect 246408 132394 246436 171158
rect 246580 158772 246632 158778
rect 246580 158714 246632 158720
rect 246396 132388 246448 132394
rect 246396 132330 246448 132336
rect 246488 131164 246540 131170
rect 246488 131106 246540 131112
rect 246304 126948 246356 126954
rect 246304 126890 246356 126896
rect 246304 118856 246356 118862
rect 246304 118798 246356 118804
rect 245200 108928 245252 108934
rect 245200 108870 245252 108876
rect 245108 107772 245160 107778
rect 245108 107714 245160 107720
rect 245120 58750 245148 107714
rect 245108 58744 245160 58750
rect 245108 58686 245160 58692
rect 245016 33788 245068 33794
rect 245016 33730 245068 33736
rect 246316 13190 246344 118798
rect 246396 117428 246448 117434
rect 246396 117370 246448 117376
rect 246408 21486 246436 117370
rect 246500 61470 246528 131106
rect 246592 124914 246620 158714
rect 247052 146198 247080 218690
rect 247132 191140 247184 191146
rect 247132 191082 247184 191088
rect 247144 162178 247172 191082
rect 247224 177336 247276 177342
rect 247224 177278 247276 177284
rect 247132 162172 247184 162178
rect 247132 162114 247184 162120
rect 247236 160070 247264 177278
rect 247684 161560 247736 161566
rect 247684 161502 247736 161508
rect 247224 160064 247276 160070
rect 247224 160006 247276 160012
rect 247040 146192 247092 146198
rect 247040 146134 247092 146140
rect 246672 131776 246724 131782
rect 246672 131718 246724 131724
rect 246580 124908 246632 124914
rect 246580 124850 246632 124856
rect 246684 122738 246712 131718
rect 246672 122732 246724 122738
rect 246672 122674 246724 122680
rect 247696 121378 247724 161502
rect 247868 160268 247920 160274
rect 247868 160210 247920 160216
rect 247776 128444 247828 128450
rect 247776 128386 247828 128392
rect 247684 121372 247736 121378
rect 247684 121314 247736 121320
rect 247684 118788 247736 118794
rect 247684 118730 247736 118736
rect 246580 99408 246632 99414
rect 246580 99350 246632 99356
rect 246488 61464 246540 61470
rect 246488 61406 246540 61412
rect 246592 50386 246620 99350
rect 246580 50380 246632 50386
rect 246580 50322 246632 50328
rect 246396 21480 246448 21486
rect 246396 21422 246448 21428
rect 247696 15910 247724 118730
rect 247788 35222 247816 128386
rect 247880 120086 247908 160210
rect 248432 144906 248460 269078
rect 249800 185700 249852 185706
rect 249800 185642 249852 185648
rect 248604 184340 248656 184346
rect 248604 184282 248656 184288
rect 248512 180464 248564 180470
rect 248512 180406 248564 180412
rect 248420 144900 248472 144906
rect 248420 144842 248472 144848
rect 248524 140622 248552 180406
rect 248616 161430 248644 184282
rect 249064 164892 249116 164898
rect 249064 164834 249116 164840
rect 248604 161424 248656 161430
rect 248604 161366 248656 161372
rect 248512 140616 248564 140622
rect 248512 140558 248564 140564
rect 249076 128246 249104 164834
rect 249812 146266 249840 185642
rect 250536 167136 250588 167142
rect 250536 167078 250588 167084
rect 250444 156052 250496 156058
rect 250444 155994 250496 156000
rect 250456 149802 250484 155994
rect 250444 149796 250496 149802
rect 250444 149738 250496 149744
rect 249800 146260 249852 146266
rect 249800 146202 249852 146208
rect 249340 137284 249392 137290
rect 249340 137226 249392 137232
rect 249064 128240 249116 128246
rect 249064 128182 249116 128188
rect 249156 127016 249208 127022
rect 249156 126958 249208 126964
rect 249064 120216 249116 120222
rect 249064 120158 249116 120164
rect 247868 120080 247920 120086
rect 247868 120022 247920 120028
rect 247868 103624 247920 103630
rect 247868 103566 247920 103572
rect 247880 66910 247908 103566
rect 247868 66904 247920 66910
rect 247868 66846 247920 66852
rect 247776 35216 247828 35222
rect 247776 35158 247828 35164
rect 249076 17338 249104 120158
rect 249168 29646 249196 126958
rect 249248 106412 249300 106418
rect 249248 106354 249300 106360
rect 249260 62830 249288 106354
rect 249352 100638 249380 137226
rect 250548 128314 250576 167078
rect 250720 149116 250772 149122
rect 250720 149058 250772 149064
rect 250536 128308 250588 128314
rect 250536 128250 250588 128256
rect 250444 127084 250496 127090
rect 250444 127026 250496 127032
rect 249340 100632 249392 100638
rect 249340 100574 249392 100580
rect 249248 62824 249300 62830
rect 249248 62766 249300 62772
rect 249156 29640 249208 29646
rect 249156 29582 249208 29588
rect 250456 28286 250484 127026
rect 250628 113348 250680 113354
rect 250628 113290 250680 113296
rect 250536 107840 250588 107846
rect 250536 107782 250588 107788
rect 250548 33862 250576 107782
rect 250640 47598 250668 113290
rect 250732 109002 250760 149058
rect 250812 140888 250864 140894
rect 250812 140830 250864 140836
rect 250720 108996 250772 109002
rect 250720 108938 250772 108944
rect 250824 102814 250852 140830
rect 250812 102808 250864 102814
rect 250812 102750 250864 102756
rect 250720 100904 250772 100910
rect 250720 100846 250772 100852
rect 250628 47592 250680 47598
rect 250628 47534 250680 47540
rect 250732 42090 250760 100846
rect 250720 42084 250772 42090
rect 250720 42026 250772 42032
rect 250536 33856 250588 33862
rect 250536 33798 250588 33804
rect 250444 28280 250496 28286
rect 250444 28222 250496 28228
rect 249064 17332 249116 17338
rect 249064 17274 249116 17280
rect 247684 15904 247736 15910
rect 247684 15846 247736 15852
rect 246304 13184 246356 13190
rect 246304 13126 246356 13132
rect 244924 7676 244976 7682
rect 244924 7618 244976 7624
rect 244096 5024 244148 5030
rect 244096 4966 244148 4972
rect 242164 4820 242216 4826
rect 242164 4762 242216 4768
rect 242900 3732 242952 3738
rect 242900 3674 242952 3680
rect 242912 480 242940 3674
rect 244108 480 244136 4966
rect 247592 3664 247644 3670
rect 247592 3606 247644 3612
rect 245198 3496 245254 3505
rect 245198 3431 245254 3440
rect 246394 3496 246450 3505
rect 246394 3431 246450 3440
rect 245212 480 245240 3431
rect 246408 480 246436 3431
rect 247604 480 247632 3606
rect 248786 3496 248842 3505
rect 248786 3431 248842 3440
rect 249982 3496 250038 3505
rect 249982 3431 250038 3440
rect 248800 480 248828 3431
rect 249996 480 250024 3431
rect 251192 480 251220 327694
rect 253940 308440 253992 308446
rect 253940 308382 253992 308388
rect 252560 217320 252612 217326
rect 252560 217262 252612 217268
rect 251364 191276 251416 191282
rect 251364 191218 251416 191224
rect 251272 182980 251324 182986
rect 251272 182922 251324 182928
rect 251284 139398 251312 182922
rect 251376 151706 251404 191218
rect 251456 175976 251508 175982
rect 251456 175918 251508 175924
rect 251364 151700 251416 151706
rect 251364 151642 251416 151648
rect 251468 149054 251496 175918
rect 252572 154562 252600 217262
rect 252652 188352 252704 188358
rect 252652 188294 252704 188300
rect 252560 154556 252612 154562
rect 252560 154498 252612 154504
rect 252664 151774 252692 188294
rect 253480 165776 253532 165782
rect 253480 165718 253532 165724
rect 253388 161628 253440 161634
rect 253388 161570 253440 161576
rect 253204 151904 253256 151910
rect 253204 151846 253256 151852
rect 252652 151768 252704 151774
rect 252652 151710 252704 151716
rect 251456 149048 251508 149054
rect 251456 148990 251508 148996
rect 252100 142180 252152 142186
rect 252100 142122 252152 142128
rect 251272 139392 251324 139398
rect 251272 139334 251324 139340
rect 251916 138100 251968 138106
rect 251916 138042 251968 138048
rect 251824 124296 251876 124302
rect 251824 124238 251876 124244
rect 251836 2174 251864 124238
rect 251928 26994 251956 138042
rect 252112 101454 252140 142122
rect 253216 110362 253244 151846
rect 253296 125724 253348 125730
rect 253296 125666 253348 125672
rect 253204 110356 253256 110362
rect 253204 110298 253256 110304
rect 252100 101448 252152 101454
rect 252100 101390 252152 101396
rect 252008 100836 252060 100842
rect 252008 100778 252060 100784
rect 252020 40730 252048 100778
rect 253204 99476 253256 99482
rect 253204 99418 253256 99424
rect 252008 40724 252060 40730
rect 252008 40666 252060 40672
rect 251916 26988 251968 26994
rect 251916 26930 251968 26936
rect 253216 21418 253244 99418
rect 253308 57254 253336 125666
rect 253400 121446 253428 161570
rect 253492 126313 253520 165718
rect 253572 140072 253624 140078
rect 253572 140014 253624 140020
rect 253478 126304 253534 126313
rect 253478 126239 253534 126248
rect 253388 121440 253440 121446
rect 253388 121382 253440 121388
rect 253388 111920 253440 111926
rect 253388 111862 253440 111868
rect 253296 57248 253348 57254
rect 253296 57190 253348 57196
rect 253400 49094 253428 111862
rect 253480 104984 253532 104990
rect 253480 104926 253532 104932
rect 253492 65550 253520 104926
rect 253584 100706 253612 140014
rect 253572 100700 253624 100706
rect 253572 100642 253624 100648
rect 253480 65544 253532 65550
rect 253480 65486 253532 65492
rect 253388 49088 253440 49094
rect 253388 49030 253440 49036
rect 253204 21412 253256 21418
rect 253204 21354 253256 21360
rect 253952 16574 253980 308382
rect 256700 295520 256752 295526
rect 256700 295462 256752 295468
rect 255320 294160 255372 294166
rect 255320 294102 255372 294108
rect 254032 239556 254084 239562
rect 254032 239498 254084 239504
rect 254044 136610 254072 239498
rect 254584 174004 254636 174010
rect 254584 173946 254636 173952
rect 254032 136604 254084 136610
rect 254032 136546 254084 136552
rect 254596 135182 254624 173946
rect 255332 153202 255360 294102
rect 255964 211880 256016 211886
rect 255964 211822 256016 211828
rect 255976 177342 256004 211822
rect 255964 177336 256016 177342
rect 255964 177278 256016 177284
rect 256240 168564 256292 168570
rect 256240 168506 256292 168512
rect 255964 164348 256016 164354
rect 255964 164290 256016 164296
rect 255320 153196 255372 153202
rect 255320 153138 255372 153144
rect 254768 145104 254820 145110
rect 254768 145046 254820 145052
rect 254584 135176 254636 135182
rect 254584 135118 254636 135124
rect 254676 133952 254728 133958
rect 254676 133894 254728 133900
rect 254584 120284 254636 120290
rect 254584 120226 254636 120232
rect 253952 16546 254256 16574
rect 252374 3496 252430 3505
rect 252374 3431 252430 3440
rect 253478 3496 253534 3505
rect 253478 3431 253534 3440
rect 251824 2168 251876 2174
rect 251824 2110 251876 2116
rect 252388 480 252416 3431
rect 253492 480 253520 3431
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 254596 6186 254624 120226
rect 254688 69698 254716 133894
rect 254780 104174 254808 145046
rect 255976 125594 256004 164290
rect 256148 158024 256200 158030
rect 256148 157966 256200 157972
rect 256056 128512 256108 128518
rect 256056 128454 256108 128460
rect 255964 125588 256016 125594
rect 255964 125530 256016 125536
rect 255964 117496 256016 117502
rect 255964 117438 256016 117444
rect 254768 104168 254820 104174
rect 254768 104110 254820 104116
rect 254768 99544 254820 99550
rect 254768 99486 254820 99492
rect 254676 69692 254728 69698
rect 254676 69634 254728 69640
rect 254780 43450 254808 99486
rect 254768 43444 254820 43450
rect 254768 43386 254820 43392
rect 255976 17270 256004 117438
rect 256068 37942 256096 128454
rect 256160 118658 256188 157966
rect 256252 129742 256280 168506
rect 256712 137902 256740 295462
rect 256792 181688 256844 181694
rect 256792 181630 256844 181636
rect 256804 150414 256832 181630
rect 258080 180260 258132 180266
rect 258080 180202 258132 180208
rect 257344 171284 257396 171290
rect 257344 171226 257396 171232
rect 256792 150408 256844 150414
rect 256792 150350 256844 150356
rect 256700 137896 256752 137902
rect 256700 137838 256752 137844
rect 257356 132462 257384 171226
rect 258092 157350 258120 180202
rect 258736 177313 258764 347754
rect 262220 298240 262272 298246
rect 262220 298182 262272 298188
rect 261484 213308 261536 213314
rect 261484 213250 261536 213256
rect 258816 203652 258868 203658
rect 258816 203594 258868 203600
rect 258828 180198 258856 203594
rect 260840 193928 260892 193934
rect 260840 193870 260892 193876
rect 258816 180192 258868 180198
rect 258816 180134 258868 180140
rect 259458 180160 259514 180169
rect 259458 180095 259514 180104
rect 258722 177304 258778 177313
rect 258722 177239 258778 177248
rect 258908 169924 258960 169930
rect 258908 169866 258960 169872
rect 258724 162920 258776 162926
rect 258724 162862 258776 162868
rect 258080 157344 258132 157350
rect 258080 157286 258132 157292
rect 257528 148368 257580 148374
rect 257528 148310 257580 148316
rect 257344 132456 257396 132462
rect 257344 132398 257396 132404
rect 257436 129872 257488 129878
rect 257436 129814 257488 129820
rect 256240 129736 256292 129742
rect 256240 129678 256292 129684
rect 256240 125792 256292 125798
rect 256240 125734 256292 125740
rect 256148 118652 256200 118658
rect 256148 118594 256200 118600
rect 256148 110560 256200 110566
rect 256148 110502 256200 110508
rect 256160 47666 256188 110502
rect 256252 76634 256280 125734
rect 257344 121576 257396 121582
rect 257344 121518 257396 121524
rect 256240 76628 256292 76634
rect 256240 76570 256292 76576
rect 256148 47660 256200 47666
rect 256148 47602 256200 47608
rect 256056 37936 256108 37942
rect 256056 37878 256108 37884
rect 255964 17264 256016 17270
rect 255964 17206 256016 17212
rect 257356 10402 257384 121518
rect 257448 60042 257476 129814
rect 257540 107642 257568 148310
rect 258736 122806 258764 162862
rect 258816 153332 258868 153338
rect 258816 153274 258868 153280
rect 258724 122800 258776 122806
rect 258724 122742 258776 122748
rect 258828 113150 258856 153274
rect 258920 131102 258948 169866
rect 259092 149184 259144 149190
rect 259092 149126 259144 149132
rect 258908 131096 258960 131102
rect 258908 131038 258960 131044
rect 258908 121644 258960 121650
rect 258908 121586 258960 121592
rect 258816 113144 258868 113150
rect 258816 113086 258868 113092
rect 258724 111988 258776 111994
rect 258724 111930 258776 111936
rect 257620 109132 257672 109138
rect 257620 109074 257672 109080
rect 257528 107636 257580 107642
rect 257528 107578 257580 107584
rect 257528 102332 257580 102338
rect 257528 102274 257580 102280
rect 257436 60036 257488 60042
rect 257436 59978 257488 59984
rect 257540 39370 257568 102274
rect 257632 55962 257660 109074
rect 257620 55956 257672 55962
rect 257620 55898 257672 55904
rect 257528 39364 257580 39370
rect 257528 39306 257580 39312
rect 258736 15978 258764 111930
rect 258816 104032 258868 104038
rect 258816 103974 258868 103980
rect 258828 28354 258856 103974
rect 258920 46238 258948 121586
rect 259000 116136 259052 116142
rect 259000 116078 259052 116084
rect 258908 46232 258960 46238
rect 258908 46174 258960 46180
rect 259012 44878 259040 116078
rect 259104 115258 259132 149126
rect 259472 137970 259500 180095
rect 260472 150612 260524 150618
rect 260472 150554 260524 150560
rect 259460 137964 259512 137970
rect 259460 137906 259512 137912
rect 260196 135448 260248 135454
rect 260196 135390 260248 135396
rect 260104 123004 260156 123010
rect 260104 122946 260156 122952
rect 259092 115252 259144 115258
rect 259092 115194 259144 115200
rect 259000 44872 259052 44878
rect 259000 44814 259052 44820
rect 258816 28348 258868 28354
rect 258816 28290 258868 28296
rect 260116 19990 260144 122946
rect 260208 66978 260236 135390
rect 260288 114640 260340 114646
rect 260288 114582 260340 114588
rect 260196 66972 260248 66978
rect 260196 66914 260248 66920
rect 260300 53106 260328 114582
rect 260484 110430 260512 150554
rect 260852 140690 260880 193870
rect 261496 181762 261524 213250
rect 261484 181756 261536 181762
rect 261484 181698 261536 181704
rect 261482 174448 261538 174457
rect 261482 174383 261538 174392
rect 260840 140684 260892 140690
rect 260840 140626 260892 140632
rect 261496 135250 261524 174383
rect 261760 158840 261812 158846
rect 261760 158782 261812 158788
rect 261576 146396 261628 146402
rect 261576 146338 261628 146344
rect 261484 135244 261536 135250
rect 261484 135186 261536 135192
rect 261298 130792 261354 130801
rect 261298 130727 261354 130736
rect 261312 129878 261340 130727
rect 261300 129872 261352 129878
rect 261300 129814 261352 129820
rect 261484 124364 261536 124370
rect 261484 124306 261536 124312
rect 260472 110424 260524 110430
rect 260472 110366 260524 110372
rect 260380 109200 260432 109206
rect 260380 109142 260432 109148
rect 260392 54602 260420 109142
rect 261206 98968 261262 98977
rect 261206 98903 261262 98912
rect 261220 98122 261248 98903
rect 261208 98116 261260 98122
rect 261208 98058 261260 98064
rect 260380 54596 260432 54602
rect 260380 54538 260432 54544
rect 260288 53100 260340 53106
rect 260288 53042 260340 53048
rect 261496 32502 261524 124306
rect 261588 106282 261616 146338
rect 261668 134088 261720 134094
rect 261668 134030 261720 134036
rect 261576 106276 261628 106282
rect 261576 106218 261628 106224
rect 261574 100600 261630 100609
rect 261574 100535 261630 100544
rect 261588 38010 261616 100535
rect 261680 71126 261708 134030
rect 261772 133822 261800 158782
rect 262232 140758 262260 298182
rect 264256 181626 264284 400279
rect 269764 397520 269816 397526
rect 269764 397462 269816 397468
rect 267004 319524 267056 319530
rect 267004 319466 267056 319472
rect 266360 307080 266412 307086
rect 266360 307022 266412 307028
rect 265624 217388 265676 217394
rect 265624 217330 265676 217336
rect 264336 205080 264388 205086
rect 264336 205022 264388 205028
rect 264348 182782 264376 205022
rect 264336 182776 264388 182782
rect 264336 182718 264388 182724
rect 264244 181620 264296 181626
rect 264244 181562 264296 181568
rect 265636 177449 265664 217330
rect 265622 177440 265678 177449
rect 265622 177375 265678 177384
rect 264426 175808 264482 175817
rect 264426 175743 264482 175752
rect 264440 173942 264468 175743
rect 265714 174992 265770 175001
rect 265714 174927 265770 174936
rect 264428 173936 264480 173942
rect 264428 173878 264480 173884
rect 265728 173194 265756 174927
rect 265806 174176 265862 174185
rect 265806 174111 265862 174120
rect 265820 174010 265848 174111
rect 265808 174004 265860 174010
rect 265808 173946 265860 173952
rect 265898 173224 265954 173233
rect 265716 173188 265768 173194
rect 265898 173159 265954 173168
rect 265716 173130 265768 173136
rect 265530 172816 265586 172825
rect 265530 172751 265586 172760
rect 265544 172650 265572 172751
rect 262864 172644 262916 172650
rect 262864 172586 262916 172592
rect 265532 172644 265584 172650
rect 265532 172586 265584 172592
rect 262220 140752 262272 140758
rect 262220 140694 262272 140700
rect 262876 133890 262904 172586
rect 265912 172582 265940 173159
rect 265900 172576 265952 172582
rect 265714 172544 265770 172553
rect 265900 172518 265952 172524
rect 265714 172479 265770 172488
rect 265622 171592 265678 171601
rect 265622 171527 265678 171536
rect 265636 171290 265664 171527
rect 265624 171284 265676 171290
rect 265624 171226 265676 171232
rect 265438 170640 265494 170649
rect 265438 170575 265494 170584
rect 265254 170232 265310 170241
rect 265254 170167 265310 170176
rect 265268 169930 265296 170167
rect 265256 169924 265308 169930
rect 265256 169866 265308 169872
rect 265452 169862 265480 170575
rect 265440 169856 265492 169862
rect 265440 169798 265492 169804
rect 265622 169824 265678 169833
rect 265622 169759 265624 169768
rect 265676 169759 265678 169768
rect 265624 169730 265676 169736
rect 265346 169008 265402 169017
rect 265346 168943 265402 168952
rect 265360 168570 265388 168943
rect 265622 168600 265678 168609
rect 265348 168564 265400 168570
rect 265622 168535 265678 168544
rect 265348 168506 265400 168512
rect 265254 168464 265310 168473
rect 265636 168434 265664 168535
rect 265254 168399 265310 168408
rect 265624 168428 265676 168434
rect 264428 167068 264480 167074
rect 264428 167010 264480 167016
rect 264440 166841 264468 167010
rect 264426 166832 264482 166841
rect 264426 166767 264482 166776
rect 265268 164898 265296 168399
rect 265624 168370 265676 168376
rect 265346 167648 265402 167657
rect 265346 167583 265402 167592
rect 265360 167142 265388 167583
rect 265348 167136 265400 167142
rect 265348 167078 265400 167084
rect 265728 166994 265756 172479
rect 265898 172000 265954 172009
rect 265898 171935 265954 171944
rect 265808 171216 265860 171222
rect 265806 171184 265808 171193
rect 265860 171184 265862 171193
rect 265912 171154 265940 171935
rect 265806 171119 265862 171128
rect 265900 171148 265952 171154
rect 265900 171090 265952 171096
rect 265806 169416 265862 169425
rect 265806 169351 265862 169360
rect 265820 168502 265848 169351
rect 265808 168496 265860 168502
rect 265808 168438 265860 168444
rect 265636 166966 265756 166994
rect 265346 166016 265402 166025
rect 265346 165951 265402 165960
rect 265360 165646 265388 165951
rect 265348 165640 265400 165646
rect 265348 165582 265400 165588
rect 265346 165064 265402 165073
rect 265346 164999 265402 165008
rect 265256 164892 265308 164898
rect 265256 164834 265308 164840
rect 265162 164656 265218 164665
rect 265162 164591 265218 164600
rect 265176 164354 265204 164591
rect 265164 164348 265216 164354
rect 265164 164290 265216 164296
rect 265360 164286 265388 164999
rect 265348 164280 265400 164286
rect 265162 164248 265218 164257
rect 265348 164222 265400 164228
rect 265162 164183 265218 164192
rect 264242 163840 264298 163849
rect 264242 163775 264298 163784
rect 263140 154760 263192 154766
rect 263140 154702 263192 154708
rect 262956 143608 263008 143614
rect 262956 143550 263008 143556
rect 262968 141409 262996 143550
rect 262954 141400 263010 141409
rect 262954 141335 263010 141344
rect 262956 134020 263008 134026
rect 262956 133962 263008 133968
rect 262864 133884 262916 133890
rect 262864 133826 262916 133832
rect 261760 133816 261812 133822
rect 261760 133758 261812 133764
rect 262864 122936 262916 122942
rect 262864 122878 262916 122884
rect 261760 107704 261812 107710
rect 261760 107646 261812 107652
rect 261668 71120 261720 71126
rect 261668 71062 261720 71068
rect 261772 57322 261800 107646
rect 261760 57316 261812 57322
rect 261760 57258 261812 57264
rect 261576 38004 261628 38010
rect 261576 37946 261628 37952
rect 261484 32496 261536 32502
rect 261484 32438 261536 32444
rect 260104 19984 260156 19990
rect 260104 19926 260156 19932
rect 258724 15972 258776 15978
rect 258724 15914 258776 15920
rect 261760 13252 261812 13258
rect 261760 13194 261812 13200
rect 257344 10396 257396 10402
rect 257344 10338 257396 10344
rect 260656 6384 260708 6390
rect 260656 6326 260708 6332
rect 254584 6180 254636 6186
rect 254584 6122 254636 6128
rect 257066 4856 257122 4865
rect 257066 4791 257122 4800
rect 255870 3496 255926 3505
rect 255870 3431 255926 3440
rect 255884 480 255912 3431
rect 257080 480 257108 4791
rect 259458 3496 259514 3505
rect 259458 3431 259514 3440
rect 258262 3360 258318 3369
rect 258262 3295 258318 3304
rect 258276 480 258304 3295
rect 259472 480 259500 3431
rect 260668 480 260696 6326
rect 261772 480 261800 13194
rect 262876 9042 262904 122878
rect 262968 68406 262996 133962
rect 263048 132660 263100 132666
rect 263048 132602 263100 132608
rect 263060 75274 263088 132602
rect 263152 123486 263180 154702
rect 264256 133113 264284 163775
rect 265176 163538 265204 164183
rect 265164 163532 265216 163538
rect 265164 163474 265216 163480
rect 265636 163282 265664 166966
rect 265714 166424 265770 166433
rect 265714 166359 265770 166368
rect 265728 165714 265756 166359
rect 265808 165776 265860 165782
rect 265806 165744 265808 165753
rect 265860 165744 265862 165753
rect 265716 165708 265768 165714
rect 265806 165679 265862 165688
rect 265716 165650 265768 165656
rect 265806 163432 265862 163441
rect 265806 163367 265862 163376
rect 265452 163254 265664 163282
rect 264518 162480 264574 162489
rect 264518 162415 264574 162424
rect 264426 161936 264482 161945
rect 264426 161871 264482 161880
rect 264440 161634 264468 161871
rect 264428 161628 264480 161634
rect 264428 161570 264480 161576
rect 264532 161498 264560 162415
rect 264520 161492 264572 161498
rect 264520 161434 264572 161440
rect 265452 158846 265480 163254
rect 265820 163062 265848 163367
rect 265808 163056 265860 163062
rect 265530 163024 265586 163033
rect 265808 162998 265860 163004
rect 265530 162959 265586 162968
rect 265544 162926 265572 162959
rect 265532 162920 265584 162926
rect 265532 162862 265584 162868
rect 265530 161664 265586 161673
rect 265530 161599 265586 161608
rect 265544 161566 265572 161599
rect 265532 161560 265584 161566
rect 265532 161502 265584 161508
rect 265990 160848 266046 160857
rect 265990 160783 266046 160792
rect 265898 160440 265954 160449
rect 265898 160375 265954 160384
rect 265912 160274 265940 160375
rect 265900 160268 265952 160274
rect 265900 160210 265952 160216
rect 265808 160200 265860 160206
rect 265806 160168 265808 160177
rect 265860 160168 265862 160177
rect 266004 160138 266032 160783
rect 265806 160103 265862 160112
rect 265992 160132 266044 160138
rect 265992 160074 266044 160080
rect 265622 159896 265678 159905
rect 265622 159831 265678 159840
rect 265530 159488 265586 159497
rect 265530 159423 265586 159432
rect 265440 158840 265492 158846
rect 265440 158782 265492 158788
rect 265544 158778 265572 159423
rect 265532 158772 265584 158778
rect 265532 158714 265584 158720
rect 265070 157448 265126 157457
rect 265070 157383 265126 157392
rect 265084 156670 265112 157383
rect 265072 156664 265124 156670
rect 265072 156606 265124 156612
rect 265346 153912 265402 153921
rect 265346 153847 265402 153856
rect 265360 153270 265388 153847
rect 265348 153264 265400 153270
rect 265348 153206 265400 153212
rect 264334 152688 264390 152697
rect 264334 152623 264390 152632
rect 264242 133104 264298 133113
rect 264242 133039 264298 133048
rect 263140 123480 263192 123486
rect 263140 123422 263192 123428
rect 264242 119096 264298 119105
rect 264242 119031 264298 119040
rect 263140 105052 263192 105058
rect 263140 104994 263192 105000
rect 263048 75268 263100 75274
rect 263048 75210 263100 75216
rect 262956 68400 263008 68406
rect 262956 68342 263008 68348
rect 263152 64190 263180 104994
rect 263140 64184 263192 64190
rect 263140 64126 263192 64132
rect 262956 9172 263008 9178
rect 262956 9114 263008 9120
rect 262864 9036 262916 9042
rect 262864 8978 262916 8984
rect 262968 480 262996 9114
rect 264256 7614 264284 119031
rect 264348 111790 264376 152623
rect 265254 152144 265310 152153
rect 265254 152079 265310 152088
rect 265268 151978 265296 152079
rect 265256 151972 265308 151978
rect 265256 151914 265308 151920
rect 265438 150920 265494 150929
rect 265438 150855 265494 150864
rect 265452 150482 265480 150855
rect 265440 150476 265492 150482
rect 265440 150418 265492 150424
rect 265346 149696 265402 149705
rect 265346 149631 265402 149640
rect 265360 149190 265388 149631
rect 265348 149184 265400 149190
rect 265348 149126 265400 149132
rect 265438 149152 265494 149161
rect 265438 149087 265494 149096
rect 265452 148374 265480 149087
rect 265530 148744 265586 148753
rect 265530 148679 265586 148688
rect 265440 148368 265492 148374
rect 265440 148310 265492 148316
rect 265070 147928 265126 147937
rect 265070 147863 265126 147872
rect 265084 146946 265112 147863
rect 265544 147694 265572 148679
rect 265532 147688 265584 147694
rect 265532 147630 265584 147636
rect 265072 146940 265124 146946
rect 265072 146882 265124 146888
rect 265530 146704 265586 146713
rect 265530 146639 265586 146648
rect 265544 146334 265572 146639
rect 265532 146328 265584 146334
rect 265532 146270 265584 146276
rect 265438 146160 265494 146169
rect 265438 146095 265494 146104
rect 264978 143168 265034 143177
rect 264978 143103 265034 143112
rect 264992 140842 265020 143103
rect 265452 142905 265480 146095
rect 265530 144528 265586 144537
rect 265530 144463 265586 144472
rect 265544 143614 265572 144463
rect 265532 143608 265584 143614
rect 265532 143550 265584 143556
rect 265438 142896 265494 142905
rect 265438 142831 265494 142840
rect 265346 142760 265402 142769
rect 265346 142695 265402 142704
rect 265254 142216 265310 142225
rect 265360 142186 265388 142695
rect 265254 142151 265310 142160
rect 265348 142180 265400 142186
rect 264428 140820 264480 140826
rect 264428 140762 264480 140768
rect 264624 140814 265020 140842
rect 264440 140593 264468 140762
rect 264426 140584 264482 140593
rect 264426 140519 264482 140528
rect 264428 133952 264480 133958
rect 264428 133894 264480 133900
rect 264440 133793 264468 133894
rect 264426 133784 264482 133793
rect 264426 133719 264482 133728
rect 264426 130656 264482 130665
rect 264426 130591 264482 130600
rect 264440 129810 264468 130591
rect 264428 129804 264480 129810
rect 264428 129746 264480 129752
rect 264428 128512 264480 128518
rect 264428 128454 264480 128460
rect 264440 128217 264468 128454
rect 264426 128208 264482 128217
rect 264426 128143 264482 128152
rect 264428 127016 264480 127022
rect 264428 126958 264480 126964
rect 264440 126857 264468 126958
rect 264426 126848 264482 126857
rect 264426 126783 264482 126792
rect 264428 123004 264480 123010
rect 264428 122946 264480 122952
rect 264440 122641 264468 122946
rect 264426 122632 264482 122641
rect 264426 122567 264482 122576
rect 264428 121644 264480 121650
rect 264428 121586 264480 121592
rect 264440 121281 264468 121586
rect 264426 121272 264482 121281
rect 264426 121207 264482 121216
rect 264426 117328 264482 117337
rect 264426 117263 264482 117272
rect 264440 116006 264468 117263
rect 264428 116000 264480 116006
rect 264428 115942 264480 115948
rect 264336 111784 264388 111790
rect 264336 111726 264388 111732
rect 264426 111344 264482 111353
rect 264426 111279 264482 111288
rect 264334 101960 264390 101969
rect 264334 101895 264390 101904
rect 264348 14482 264376 101895
rect 264440 31074 264468 111279
rect 264520 107772 264572 107778
rect 264520 107714 264572 107720
rect 264532 107545 264560 107714
rect 264518 107536 264574 107545
rect 264518 107471 264574 107480
rect 264518 107128 264574 107137
rect 264518 107063 264574 107072
rect 264532 61402 264560 107063
rect 264624 102134 264652 140814
rect 265162 138136 265218 138145
rect 265162 138071 265164 138080
rect 265216 138071 265218 138080
rect 265164 138042 265216 138048
rect 265268 137290 265296 142151
rect 265348 142122 265400 142128
rect 265530 140992 265586 141001
rect 265530 140927 265586 140936
rect 265544 140894 265572 140927
rect 265532 140888 265584 140894
rect 265532 140830 265584 140836
rect 265636 138014 265664 159831
rect 265806 158808 265862 158817
rect 265806 158743 265862 158752
rect 265820 158030 265848 158743
rect 265990 158264 266046 158273
rect 265990 158199 266046 158208
rect 265808 158024 265860 158030
rect 265808 157966 265860 157972
rect 265806 157856 265862 157865
rect 265806 157791 265862 157800
rect 265820 157486 265848 157791
rect 265808 157480 265860 157486
rect 265808 157422 265860 157428
rect 266004 157418 266032 158199
rect 265992 157412 266044 157418
rect 265992 157354 266044 157360
rect 265898 156904 265954 156913
rect 265898 156839 265954 156848
rect 265806 156088 265862 156097
rect 265912 156058 265940 156839
rect 266082 156496 266138 156505
rect 266082 156431 266138 156440
rect 265806 156023 265862 156032
rect 265900 156052 265952 156058
rect 265820 155990 265848 156023
rect 265900 155994 265952 156000
rect 265808 155984 265860 155990
rect 265808 155926 265860 155932
rect 265714 155680 265770 155689
rect 265714 155615 265770 155624
rect 265728 154630 265756 155615
rect 265990 155272 266046 155281
rect 265990 155207 266046 155216
rect 265806 154864 265862 154873
rect 265806 154799 265862 154808
rect 265820 154766 265848 154799
rect 265808 154760 265860 154766
rect 265808 154702 265860 154708
rect 265898 154728 265954 154737
rect 266004 154698 266032 155207
rect 265898 154663 265954 154672
rect 265992 154692 266044 154698
rect 265716 154624 265768 154630
rect 265716 154566 265768 154572
rect 265912 153882 265940 154663
rect 265992 154634 266044 154640
rect 265900 153876 265952 153882
rect 265900 153818 265952 153824
rect 265806 153504 265862 153513
rect 265806 153439 265862 153448
rect 265820 153338 265848 153439
rect 265808 153332 265860 153338
rect 265808 153274 265860 153280
rect 265898 153232 265954 153241
rect 265898 153167 265954 153176
rect 265808 151904 265860 151910
rect 265806 151872 265808 151881
rect 265860 151872 265862 151881
rect 265806 151807 265862 151816
rect 265714 151328 265770 151337
rect 265714 151263 265770 151272
rect 265728 150618 265756 151263
rect 265716 150612 265768 150618
rect 265716 150554 265768 150560
rect 265808 150544 265860 150550
rect 265806 150512 265808 150521
rect 265860 150512 265862 150521
rect 265806 150447 265862 150456
rect 265806 150104 265862 150113
rect 265806 150039 265862 150048
rect 265820 149122 265848 150039
rect 265912 149734 265940 153167
rect 266096 152425 266124 156431
rect 266082 152416 266138 152425
rect 266082 152351 266138 152360
rect 265900 149728 265952 149734
rect 265900 149670 265952 149676
rect 265808 149116 265860 149122
rect 265808 149058 265860 149064
rect 265714 148336 265770 148345
rect 265714 148271 265770 148280
rect 265728 147762 265756 148271
rect 265716 147756 265768 147762
rect 265716 147698 265768 147704
rect 265898 147112 265954 147121
rect 265898 147047 265954 147056
rect 265912 146402 265940 147047
rect 265990 146568 266046 146577
rect 265990 146503 266046 146512
rect 265900 146396 265952 146402
rect 265900 146338 265952 146344
rect 265806 145752 265862 145761
rect 265806 145687 265862 145696
rect 265714 145344 265770 145353
rect 265714 145279 265770 145288
rect 265728 145042 265756 145279
rect 265716 145036 265768 145042
rect 265716 144978 265768 144984
rect 265820 144974 265848 145687
rect 265900 145104 265952 145110
rect 265900 145046 265952 145052
rect 265808 144968 265860 144974
rect 265912 144945 265940 145046
rect 265808 144910 265860 144916
rect 265898 144936 265954 144945
rect 265898 144871 265954 144880
rect 266004 144226 266032 146503
rect 265992 144220 266044 144226
rect 265992 144162 266044 144168
rect 265806 143576 265862 143585
rect 265806 143511 265862 143520
rect 265820 142866 265848 143511
rect 265808 142860 265860 142866
rect 265808 142802 265860 142808
rect 265806 142352 265862 142361
rect 265806 142287 265862 142296
rect 265820 140078 265848 142287
rect 265898 141400 265954 141409
rect 265898 141335 265954 141344
rect 265808 140072 265860 140078
rect 265808 140014 265860 140020
rect 265714 139768 265770 139777
rect 265714 139703 265770 139712
rect 265728 139466 265756 139703
rect 265808 139528 265860 139534
rect 265806 139496 265808 139505
rect 265860 139496 265862 139505
rect 265716 139460 265768 139466
rect 265806 139431 265862 139440
rect 265716 139402 265768 139408
rect 265806 138408 265862 138417
rect 265806 138343 265862 138352
rect 265820 138038 265848 138343
rect 265544 137986 265664 138014
rect 265808 138032 265860 138038
rect 265256 137284 265308 137290
rect 265256 137226 265308 137232
rect 265164 135448 265216 135454
rect 265164 135390 265216 135396
rect 265176 135289 265204 135390
rect 265162 135280 265218 135289
rect 265162 135215 265218 135224
rect 265254 134600 265310 134609
rect 265254 134535 265310 134544
rect 265268 134026 265296 134535
rect 265256 134020 265308 134026
rect 265256 133962 265308 133968
rect 265544 131782 265572 137986
rect 265808 137974 265860 137980
rect 265806 137592 265862 137601
rect 265806 137527 265862 137536
rect 265714 137184 265770 137193
rect 265714 137119 265770 137128
rect 265728 136746 265756 137119
rect 265716 136740 265768 136746
rect 265716 136682 265768 136688
rect 265820 136678 265848 137527
rect 265808 136672 265860 136678
rect 265808 136614 265860 136620
rect 265806 135416 265862 135425
rect 265806 135351 265808 135360
rect 265860 135351 265862 135360
rect 265808 135322 265860 135328
rect 265806 134192 265862 134201
rect 265806 134127 265862 134136
rect 265820 134094 265848 134127
rect 265808 134088 265860 134094
rect 265808 134030 265860 134036
rect 265622 132832 265678 132841
rect 265622 132767 265678 132776
rect 265636 132666 265664 132767
rect 265624 132660 265676 132666
rect 265624 132602 265676 132608
rect 265714 132016 265770 132025
rect 265714 131951 265770 131960
rect 265532 131776 265584 131782
rect 265532 131718 265584 131724
rect 265622 131200 265678 131209
rect 265728 131170 265756 131951
rect 265622 131135 265678 131144
rect 265716 131164 265768 131170
rect 265346 129024 265402 129033
rect 265346 128959 265402 128968
rect 265360 128382 265388 128959
rect 265348 128376 265400 128382
rect 265636 128354 265664 131135
rect 265716 131106 265768 131112
rect 265806 128616 265862 128625
rect 265806 128551 265862 128560
rect 265820 128450 265848 128551
rect 265808 128444 265860 128450
rect 265808 128386 265860 128392
rect 265348 128318 265400 128324
rect 265452 128326 265664 128354
rect 265346 127664 265402 127673
rect 265346 127599 265402 127608
rect 265360 127090 265388 127599
rect 265348 127084 265400 127090
rect 265348 127026 265400 127032
rect 265452 118694 265480 128326
rect 265806 126440 265862 126449
rect 265806 126375 265862 126384
rect 265622 126032 265678 126041
rect 265622 125967 265678 125976
rect 265636 125662 265664 125967
rect 265716 125792 265768 125798
rect 265716 125734 265768 125740
rect 265624 125656 265676 125662
rect 265728 125633 265756 125734
rect 265820 125730 265848 126375
rect 265808 125724 265860 125730
rect 265808 125666 265860 125672
rect 265624 125598 265676 125604
rect 265714 125624 265770 125633
rect 265714 125559 265770 125568
rect 265912 125202 265940 141335
rect 266082 136776 266138 136785
rect 266082 136711 266138 136720
rect 265990 136368 266046 136377
rect 265990 136303 266046 136312
rect 266004 135318 266032 136303
rect 265992 135312 266044 135318
rect 265992 135254 266044 135260
rect 265636 125174 265940 125202
rect 265532 124364 265584 124370
rect 265532 124306 265584 124312
rect 265544 124273 265572 124306
rect 265530 124264 265586 124273
rect 265530 124199 265586 124208
rect 265636 119626 265664 125174
rect 265806 125080 265862 125089
rect 265806 125015 265862 125024
rect 265820 124302 265848 125015
rect 265898 124672 265954 124681
rect 265898 124607 265954 124616
rect 265808 124296 265860 124302
rect 265808 124238 265860 124244
rect 265912 124234 265940 124607
rect 265900 124228 265952 124234
rect 265900 124170 265952 124176
rect 265898 123448 265954 123457
rect 265898 123383 265954 123392
rect 265806 123040 265862 123049
rect 265806 122975 265862 122984
rect 265820 122942 265848 122975
rect 265808 122936 265860 122942
rect 265808 122878 265860 122884
rect 265912 122874 265940 123383
rect 265900 122868 265952 122874
rect 265900 122810 265952 122816
rect 265898 122088 265954 122097
rect 265898 122023 265954 122032
rect 265806 121680 265862 121689
rect 265806 121615 265862 121624
rect 265820 121514 265848 121615
rect 265912 121582 265940 122023
rect 265900 121576 265952 121582
rect 265900 121518 265952 121524
rect 265808 121508 265860 121514
rect 265808 121450 265860 121456
rect 265990 120864 266046 120873
rect 265990 120799 266046 120808
rect 265898 120456 265954 120465
rect 265898 120391 265954 120400
rect 265808 120284 265860 120290
rect 265808 120226 265860 120232
rect 265820 120193 265848 120226
rect 265912 120222 265940 120391
rect 265900 120216 265952 120222
rect 265806 120184 265862 120193
rect 265900 120158 265952 120164
rect 266004 120154 266032 120799
rect 265806 120119 265862 120128
rect 265992 120148 266044 120154
rect 265992 120090 266044 120096
rect 265544 119598 265664 119626
rect 265544 119406 265572 119598
rect 265622 119504 265678 119513
rect 265622 119439 265678 119448
rect 265532 119400 265584 119406
rect 265532 119342 265584 119348
rect 265532 118856 265584 118862
rect 265530 118824 265532 118833
rect 265584 118824 265586 118833
rect 265636 118794 265664 119439
rect 265530 118759 265586 118768
rect 265624 118788 265676 118794
rect 265624 118730 265676 118736
rect 266096 118694 266124 136711
rect 265452 118666 265756 118694
rect 265162 118280 265218 118289
rect 265162 118215 265218 118224
rect 265176 117366 265204 118215
rect 265164 117360 265216 117366
rect 265164 117302 265216 117308
rect 265530 116920 265586 116929
rect 265530 116855 265586 116864
rect 265544 116142 265572 116855
rect 265622 116512 265678 116521
rect 265622 116447 265678 116456
rect 265532 116136 265584 116142
rect 265532 116078 265584 116084
rect 265636 116074 265664 116447
rect 265624 116068 265676 116074
rect 265624 116010 265676 116016
rect 265622 115288 265678 115297
rect 265622 115223 265678 115232
rect 265438 114880 265494 114889
rect 265438 114815 265494 114824
rect 265452 114646 265480 114815
rect 265440 114640 265492 114646
rect 265440 114582 265492 114588
rect 265636 114578 265664 115223
rect 265624 114572 265676 114578
rect 265624 114514 265676 114520
rect 265530 113928 265586 113937
rect 265530 113863 265586 113872
rect 265438 113520 265494 113529
rect 265438 113455 265494 113464
rect 265452 113286 265480 113455
rect 265544 113354 265572 113863
rect 265532 113348 265584 113354
rect 265532 113290 265584 113296
rect 265440 113280 265492 113286
rect 265440 113222 265492 113228
rect 265530 112704 265586 112713
rect 265530 112639 265586 112648
rect 265544 111858 265572 112639
rect 265622 112296 265678 112305
rect 265622 112231 265678 112240
rect 265636 111994 265664 112231
rect 265624 111988 265676 111994
rect 265624 111930 265676 111936
rect 265532 111852 265584 111858
rect 265532 111794 265584 111800
rect 265162 110936 265218 110945
rect 265162 110871 265218 110880
rect 265176 110566 265204 110871
rect 265164 110560 265216 110566
rect 265164 110502 265216 110508
rect 265530 110120 265586 110129
rect 265530 110055 265586 110064
rect 265544 109070 265572 110055
rect 265532 109064 265584 109070
rect 265532 109006 265584 109012
rect 265346 108352 265402 108361
rect 265346 108287 265402 108296
rect 265360 107710 265388 108287
rect 265348 107704 265400 107710
rect 265348 107646 265400 107652
rect 265254 105768 265310 105777
rect 265254 105703 265310 105712
rect 265268 105058 265296 105703
rect 265256 105052 265308 105058
rect 265256 104994 265308 105000
rect 265622 104952 265678 104961
rect 265622 104887 265624 104896
rect 265676 104887 265678 104896
rect 265624 104858 265676 104864
rect 265622 104544 265678 104553
rect 265622 104479 265678 104488
rect 265636 104038 265664 104479
rect 265624 104032 265676 104038
rect 265624 103974 265676 103980
rect 265530 103184 265586 103193
rect 265530 103119 265586 103128
rect 265346 102368 265402 102377
rect 265346 102303 265348 102312
rect 265400 102303 265402 102312
rect 265348 102274 265400 102280
rect 265544 102270 265572 103119
rect 265622 102776 265678 102785
rect 265622 102711 265678 102720
rect 265532 102264 265584 102270
rect 265532 102206 265584 102212
rect 265636 102202 265664 102711
rect 265624 102196 265676 102202
rect 265624 102138 265676 102144
rect 264612 102128 264664 102134
rect 264612 102070 264664 102076
rect 265162 99784 265218 99793
rect 265162 99719 265218 99728
rect 265176 99414 265204 99719
rect 265622 99512 265678 99521
rect 265622 99447 265624 99456
rect 265676 99447 265678 99456
rect 265624 99418 265676 99424
rect 265164 99408 265216 99414
rect 265164 99350 265216 99356
rect 264610 98832 264666 98841
rect 264610 98767 264666 98776
rect 264624 98054 264652 98767
rect 264612 98048 264664 98054
rect 264612 97990 264664 97996
rect 265622 97608 265678 97617
rect 265622 97543 265678 97552
rect 265346 97200 265402 97209
rect 265346 97135 265402 97144
rect 265360 96694 265388 97135
rect 265348 96688 265400 96694
rect 265348 96630 265400 96636
rect 265530 95704 265586 95713
rect 265530 95639 265586 95648
rect 265544 95266 265572 95639
rect 265532 95260 265584 95266
rect 265532 95202 265584 95208
rect 264520 61396 264572 61402
rect 264520 61338 264572 61344
rect 264428 31068 264480 31074
rect 264428 31010 264480 31016
rect 264336 14476 264388 14482
rect 264336 14418 264388 14424
rect 265636 11762 265664 97543
rect 265728 58682 265756 118666
rect 265820 118666 266124 118694
rect 265820 89010 265848 118666
rect 265990 117872 266046 117881
rect 265990 117807 266046 117816
rect 266004 117502 266032 117807
rect 265992 117496 266044 117502
rect 265898 117464 265954 117473
rect 265992 117438 266044 117444
rect 265898 117399 265900 117408
rect 265952 117399 265954 117408
rect 265900 117370 265952 117376
rect 266082 116104 266138 116113
rect 266082 116039 266138 116048
rect 265898 113248 265954 113257
rect 265898 113183 265900 113192
rect 265952 113183 265954 113192
rect 265900 113154 265952 113160
rect 265898 112160 265954 112169
rect 265898 112095 265954 112104
rect 265912 111926 265940 112095
rect 265900 111920 265952 111926
rect 265900 111862 265952 111868
rect 265900 110628 265952 110634
rect 265900 110570 265952 110576
rect 265912 110537 265940 110570
rect 265898 110528 265954 110537
rect 265898 110463 265954 110472
rect 265990 109712 266046 109721
rect 265990 109647 266046 109656
rect 266004 109206 266032 109647
rect 265992 109200 266044 109206
rect 265898 109168 265954 109177
rect 265992 109142 266044 109148
rect 265898 109103 265900 109112
rect 265952 109103 265954 109112
rect 265900 109074 265952 109080
rect 265990 108760 266046 108769
rect 265990 108695 266046 108704
rect 265898 107944 265954 107953
rect 265898 107879 265900 107888
rect 265952 107879 265954 107888
rect 265900 107850 265952 107856
rect 266004 107846 266032 108695
rect 265992 107840 266044 107846
rect 265992 107782 266044 107788
rect 265990 106720 266046 106729
rect 265990 106655 266046 106664
rect 265898 106584 265954 106593
rect 265898 106519 265954 106528
rect 265912 106486 265940 106519
rect 265900 106480 265952 106486
rect 265900 106422 265952 106428
rect 266004 106418 266032 106655
rect 265992 106412 266044 106418
rect 265992 106354 266044 106360
rect 265898 105360 265954 105369
rect 265898 105295 265954 105304
rect 265912 104990 265940 105295
rect 265900 104984 265952 104990
rect 265900 104926 265952 104932
rect 265990 104000 266046 104009
rect 265990 103935 266046 103944
rect 266004 103630 266032 103935
rect 265992 103624 266044 103630
rect 265898 103592 265954 103601
rect 265992 103566 266044 103572
rect 265898 103527 265900 103536
rect 265952 103527 265954 103536
rect 265900 103498 265952 103504
rect 265990 101552 266046 101561
rect 265990 101487 266046 101496
rect 265898 101008 265954 101017
rect 265898 100943 265954 100952
rect 265912 100910 265940 100943
rect 265900 100904 265952 100910
rect 265900 100846 265952 100852
rect 266004 100842 266032 101487
rect 265992 100836 266044 100842
rect 265992 100778 266044 100784
rect 265898 100192 265954 100201
rect 265898 100127 265954 100136
rect 265912 99550 265940 100127
rect 265900 99544 265952 99550
rect 265900 99486 265952 99492
rect 266096 99374 266124 116039
rect 265912 99346 266124 99374
rect 265808 89004 265860 89010
rect 265808 88946 265860 88952
rect 265912 83502 265940 99346
rect 265990 96792 266046 96801
rect 265990 96727 265992 96736
rect 266044 96727 266046 96736
rect 265992 96698 266044 96704
rect 265900 83496 265952 83502
rect 265900 83438 265952 83444
rect 265716 58676 265768 58682
rect 265716 58618 265768 58624
rect 266372 16574 266400 307022
rect 266372 16546 266584 16574
rect 265624 11756 265676 11762
rect 265624 11698 265676 11704
rect 264244 7608 264296 7614
rect 264244 7550 264296 7556
rect 264152 4956 264204 4962
rect 264152 4898 264204 4904
rect 264164 480 264192 4898
rect 265348 2236 265400 2242
rect 265348 2178 265400 2184
rect 265360 480 265388 2178
rect 266556 480 266584 16546
rect 267016 3670 267044 319466
rect 268384 224256 268436 224262
rect 268384 224198 268436 224204
rect 268396 177410 268424 224198
rect 269120 182776 269172 182782
rect 269120 182718 269172 182724
rect 269132 178809 269160 182718
rect 269776 181694 269804 397462
rect 317420 395344 317472 395350
rect 317420 395286 317472 395292
rect 313278 389192 313334 389201
rect 313278 389127 313334 389136
rect 306378 386472 306434 386481
rect 306378 386407 306434 386416
rect 303620 385688 303672 385694
rect 303620 385630 303672 385636
rect 300858 384568 300914 384577
rect 300858 384503 300914 384512
rect 273996 371272 274048 371278
rect 273996 371214 274048 371220
rect 271236 351212 271288 351218
rect 271236 351154 271288 351160
rect 271144 292664 271196 292670
rect 271144 292606 271196 292612
rect 269856 278792 269908 278798
rect 269856 278734 269908 278740
rect 269764 181688 269816 181694
rect 269764 181630 269816 181636
rect 269868 178838 269896 278734
rect 269948 204944 270000 204950
rect 269948 204886 270000 204892
rect 269856 178832 269908 178838
rect 269118 178800 269174 178809
rect 269856 178774 269908 178780
rect 269118 178735 269174 178744
rect 268384 177404 268436 177410
rect 268384 177346 268436 177352
rect 269960 175817 269988 204886
rect 271156 180266 271184 292606
rect 271248 279478 271276 351154
rect 272524 302320 272576 302326
rect 272524 302262 272576 302268
rect 271236 279472 271288 279478
rect 271236 279414 271288 279420
rect 271236 231124 271288 231130
rect 271236 231066 271288 231072
rect 271248 184346 271276 231066
rect 271236 184340 271288 184346
rect 271236 184282 271288 184288
rect 271144 180260 271196 180266
rect 271144 180202 271196 180208
rect 272536 179382 272564 302262
rect 273904 292596 273956 292602
rect 273904 292538 273956 292544
rect 272616 239488 272668 239494
rect 272616 239430 272668 239436
rect 272524 179376 272576 179382
rect 272524 179318 272576 179324
rect 272628 177546 272656 239430
rect 273916 180334 273944 292538
rect 274008 278050 274036 371214
rect 282184 342916 282236 342922
rect 282184 342858 282236 342864
rect 276664 337408 276716 337414
rect 276664 337350 276716 337356
rect 273996 278044 274048 278050
rect 273996 277986 274048 277992
rect 276676 261526 276704 337350
rect 280804 309188 280856 309194
rect 280804 309130 280856 309136
rect 278044 303680 278096 303686
rect 278044 303622 278096 303628
rect 276664 261520 276716 261526
rect 276664 261462 276716 261468
rect 276664 251252 276716 251258
rect 276664 251194 276716 251200
rect 275284 242956 275336 242962
rect 275284 242898 275336 242904
rect 273996 215960 274048 215966
rect 273996 215902 274048 215908
rect 273904 180328 273956 180334
rect 273904 180270 273956 180276
rect 272616 177540 272668 177546
rect 272616 177482 272668 177488
rect 274008 176050 274036 215902
rect 273996 176044 274048 176050
rect 273996 175986 274048 175992
rect 275296 175982 275324 242898
rect 275376 198008 275428 198014
rect 275376 197950 275428 197956
rect 275388 176186 275416 197950
rect 276676 177478 276704 251194
rect 276756 238060 276808 238066
rect 276756 238002 276808 238008
rect 276768 177682 276796 238002
rect 276848 233912 276900 233918
rect 276848 233854 276900 233860
rect 276756 177676 276808 177682
rect 276756 177618 276808 177624
rect 276664 177472 276716 177478
rect 276664 177414 276716 177420
rect 275376 176180 275428 176186
rect 275376 176122 275428 176128
rect 276860 176118 276888 233854
rect 276940 195288 276992 195294
rect 276940 195230 276992 195236
rect 276952 177614 276980 195230
rect 276940 177608 276992 177614
rect 276940 177550 276992 177556
rect 278056 176225 278084 303622
rect 278136 293276 278188 293282
rect 278136 293218 278188 293224
rect 278148 181830 278176 293218
rect 280160 266484 280212 266490
rect 280160 266426 280212 266432
rect 278136 181824 278188 181830
rect 278136 181766 278188 181772
rect 279332 179376 279384 179382
rect 279332 179318 279384 179324
rect 278780 178832 278832 178838
rect 278780 178774 278832 178780
rect 278792 177177 278820 178774
rect 278778 177168 278834 177177
rect 278778 177103 278834 177112
rect 278042 176216 278098 176225
rect 278042 176151 278098 176160
rect 276848 176112 276900 176118
rect 276848 176054 276900 176060
rect 275284 175976 275336 175982
rect 275284 175918 275336 175924
rect 269946 175808 270002 175817
rect 269946 175743 270002 175752
rect 267094 175400 267150 175409
rect 267094 175335 267150 175344
rect 267108 99346 267136 175335
rect 279344 173777 279372 179318
rect 279330 173768 279386 173777
rect 279330 173703 279386 173712
rect 280172 158545 280200 266426
rect 280816 199578 280844 309130
rect 282196 236774 282224 342858
rect 293960 333260 294012 333266
rect 293960 333202 294012 333208
rect 290464 291236 290516 291242
rect 290464 291178 290516 291184
rect 287336 288448 287388 288454
rect 287336 288390 287388 288396
rect 282920 282940 282972 282946
rect 282920 282882 282972 282888
rect 282276 252612 282328 252618
rect 282276 252554 282328 252560
rect 282184 236768 282236 236774
rect 282184 236710 282236 236716
rect 280804 199572 280856 199578
rect 280804 199514 280856 199520
rect 280252 191208 280304 191214
rect 280252 191150 280304 191156
rect 280158 158536 280214 158545
rect 280158 158471 280214 158480
rect 267186 123856 267242 123865
rect 267186 123791 267242 123800
rect 267096 99340 267148 99346
rect 267096 99282 267148 99288
rect 267200 94518 267228 123791
rect 280264 107817 280292 191150
rect 282288 185706 282316 252554
rect 282276 185700 282328 185706
rect 282276 185642 282328 185648
rect 281814 184240 281870 184249
rect 281540 184204 281592 184210
rect 281814 184175 281870 184184
rect 281540 184146 281592 184152
rect 280436 182844 280488 182850
rect 280436 182786 280488 182792
rect 280344 180124 280396 180130
rect 280344 180066 280396 180072
rect 280356 165481 280384 180066
rect 280448 169425 280476 182786
rect 280434 169416 280490 169425
rect 280434 169351 280490 169360
rect 280342 165472 280398 165481
rect 280342 165407 280398 165416
rect 281552 154737 281580 184146
rect 281632 176180 281684 176186
rect 281632 176122 281684 176128
rect 281644 170105 281672 176122
rect 281828 174049 281856 184175
rect 281814 174040 281870 174049
rect 281814 173975 281870 173984
rect 282090 172408 282146 172417
rect 282090 172343 282146 172352
rect 282104 171834 282132 172343
rect 282092 171828 282144 171834
rect 282092 171770 282144 171776
rect 282274 170912 282330 170921
rect 282274 170847 282330 170856
rect 281630 170096 281686 170105
rect 281630 170031 281686 170040
rect 282288 169930 282316 170847
rect 282276 169924 282328 169930
rect 282276 169866 282328 169872
rect 281724 169788 281776 169794
rect 281724 169730 281776 169736
rect 281736 167793 281764 169730
rect 282828 169720 282880 169726
rect 282828 169662 282880 169668
rect 282840 168609 282868 169662
rect 282826 168600 282882 168609
rect 282826 168535 282882 168544
rect 282460 168360 282512 168366
rect 282460 168302 282512 168308
rect 281722 167784 281778 167793
rect 281722 167719 281778 167728
rect 282472 167113 282500 168302
rect 282458 167104 282514 167113
rect 282458 167039 282514 167048
rect 282092 167000 282144 167006
rect 282092 166942 282144 166948
rect 282104 166297 282132 166942
rect 282644 166320 282696 166326
rect 282090 166288 282146 166297
rect 282644 166262 282696 166268
rect 282090 166223 282146 166232
rect 282092 165572 282144 165578
rect 282092 165514 282144 165520
rect 282104 164801 282132 165514
rect 282090 164792 282146 164801
rect 282090 164727 282146 164736
rect 282656 163985 282684 166262
rect 282828 164212 282880 164218
rect 282828 164154 282880 164160
rect 282642 163976 282698 163985
rect 282642 163911 282698 163920
rect 282840 163169 282868 164154
rect 282826 163160 282882 163169
rect 282826 163095 282882 163104
rect 282736 162920 282788 162926
rect 282736 162862 282788 162868
rect 282552 162852 282604 162858
rect 282552 162794 282604 162800
rect 282564 161673 282592 162794
rect 282550 161664 282606 161673
rect 282550 161599 282606 161608
rect 282368 161356 282420 161362
rect 282368 161298 282420 161304
rect 282380 160177 282408 161298
rect 282366 160168 282422 160177
rect 282366 160103 282422 160112
rect 282748 159361 282776 162862
rect 282828 162784 282880 162790
rect 282828 162726 282880 162732
rect 282840 162489 282868 162726
rect 282826 162480 282882 162489
rect 282826 162415 282882 162424
rect 282828 161424 282880 161430
rect 282828 161366 282880 161372
rect 282840 160857 282868 161366
rect 282826 160848 282882 160857
rect 282826 160783 282882 160792
rect 282734 159352 282790 159361
rect 282734 159287 282790 159296
rect 282276 158704 282328 158710
rect 282276 158646 282328 158652
rect 282288 157865 282316 158646
rect 282274 157856 282330 157865
rect 282274 157791 282330 157800
rect 282828 157344 282880 157350
rect 282828 157286 282880 157292
rect 282840 157049 282868 157286
rect 282826 157040 282882 157049
rect 282826 156975 282882 156984
rect 282828 155916 282880 155922
rect 282828 155858 282880 155864
rect 282840 155553 282868 155858
rect 282826 155544 282882 155553
rect 282826 155479 282882 155488
rect 281538 154728 281594 154737
rect 281538 154663 281594 154672
rect 281908 154216 281960 154222
rect 281908 154158 281960 154164
rect 281920 154057 281948 154158
rect 281906 154048 281962 154057
rect 281906 153983 281962 153992
rect 281724 153332 281776 153338
rect 281724 153274 281776 153280
rect 281736 153241 281764 153274
rect 281722 153232 281778 153241
rect 281722 153167 281778 153176
rect 282184 153196 282236 153202
rect 282184 153138 282236 153144
rect 282196 152425 282224 153138
rect 282182 152416 282238 152425
rect 282182 152351 282238 152360
rect 282828 151768 282880 151774
rect 282826 151736 282828 151745
rect 282880 151736 282882 151745
rect 282000 151700 282052 151706
rect 282826 151671 282882 151680
rect 282000 151642 282052 151648
rect 282012 150929 282040 151642
rect 281998 150920 282054 150929
rect 281998 150855 282054 150864
rect 282828 150408 282880 150414
rect 282828 150350 282880 150356
rect 282184 150340 282236 150346
rect 282184 150282 282236 150288
rect 282196 149433 282224 150282
rect 282840 150113 282868 150350
rect 282826 150104 282882 150113
rect 282826 150039 282882 150048
rect 282182 149424 282238 149433
rect 282182 149359 282238 149368
rect 282092 148980 282144 148986
rect 282092 148922 282144 148928
rect 282104 148617 282132 148922
rect 282090 148608 282146 148617
rect 282090 148543 282146 148552
rect 281724 147620 281776 147626
rect 281724 147562 281776 147568
rect 281736 147121 281764 147562
rect 281722 147112 281778 147121
rect 281722 147047 281778 147056
rect 282826 146296 282882 146305
rect 282826 146231 282828 146240
rect 282880 146231 282882 146240
rect 282828 146202 282880 146208
rect 282736 146192 282788 146198
rect 282736 146134 282788 146140
rect 282748 145489 282776 146134
rect 282734 145480 282790 145489
rect 282734 145415 282790 145424
rect 282828 144900 282880 144906
rect 282828 144842 282880 144848
rect 282840 144809 282868 144842
rect 282826 144800 282882 144809
rect 282826 144735 282882 144744
rect 282826 143984 282882 143993
rect 282826 143919 282882 143928
rect 282840 143750 282868 143919
rect 282828 143744 282880 143750
rect 282828 143686 282880 143692
rect 282092 143540 282144 143546
rect 282092 143482 282144 143488
rect 282104 143177 282132 143482
rect 282276 143472 282328 143478
rect 282276 143414 282328 143420
rect 282090 143168 282146 143177
rect 282090 143103 282146 143112
rect 282184 142996 282236 143002
rect 282184 142938 282236 142944
rect 281908 133884 281960 133890
rect 281908 133826 281960 133832
rect 281920 133249 281948 133826
rect 281906 133240 281962 133249
rect 281906 133175 281962 133184
rect 281724 130144 281776 130150
rect 281722 130112 281724 130121
rect 281776 130112 281778 130121
rect 281722 130047 281778 130056
rect 281908 127968 281960 127974
rect 281908 127910 281960 127916
rect 281920 127809 281948 127910
rect 281906 127800 281962 127809
rect 281906 127735 281962 127744
rect 282000 124024 282052 124030
rect 281998 123992 282000 124001
rect 282052 123992 282054 124001
rect 281998 123927 282054 123936
rect 282196 123185 282224 142938
rect 282288 142497 282316 143414
rect 282274 142488 282330 142497
rect 282274 142423 282330 142432
rect 282828 142112 282880 142118
rect 282828 142054 282880 142060
rect 282736 142044 282788 142050
rect 282736 141986 282788 141992
rect 282748 140865 282776 141986
rect 282840 141681 282868 142054
rect 282826 141672 282882 141681
rect 282826 141607 282882 141616
rect 282734 140856 282790 140865
rect 282734 140791 282790 140800
rect 282828 140752 282880 140758
rect 282828 140694 282880 140700
rect 282840 140185 282868 140694
rect 282826 140176 282882 140185
rect 282826 140111 282882 140120
rect 282828 139392 282880 139398
rect 282826 139360 282828 139369
rect 282880 139360 282882 139369
rect 282736 139324 282788 139330
rect 282826 139295 282882 139304
rect 282736 139266 282788 139272
rect 282748 138553 282776 139266
rect 282734 138544 282790 138553
rect 282734 138479 282790 138488
rect 282828 137964 282880 137970
rect 282828 137906 282880 137912
rect 282840 137873 282868 137906
rect 282826 137864 282882 137873
rect 282826 137799 282882 137808
rect 282736 136604 282788 136610
rect 282736 136546 282788 136552
rect 282748 135561 282776 136546
rect 282828 136536 282880 136542
rect 282828 136478 282880 136484
rect 282840 136377 282868 136478
rect 282826 136368 282882 136377
rect 282826 136303 282882 136312
rect 282734 135552 282790 135561
rect 282734 135487 282790 135496
rect 282736 135244 282788 135250
rect 282736 135186 282788 135192
rect 282748 134065 282776 135186
rect 282828 135176 282880 135182
rect 282828 135118 282880 135124
rect 282840 134745 282868 135118
rect 282826 134736 282882 134745
rect 282826 134671 282882 134680
rect 282734 134056 282790 134065
rect 282734 133991 282790 134000
rect 282932 132494 282960 282882
rect 284576 280220 284628 280226
rect 284576 280162 284628 280168
rect 284392 207732 284444 207738
rect 284392 207674 284444 207680
rect 283012 185632 283064 185638
rect 283012 185574 283064 185580
rect 283024 147801 283052 185574
rect 284300 177540 284352 177546
rect 284300 177482 284352 177488
rect 284312 169794 284340 177482
rect 284300 169788 284352 169794
rect 284300 169730 284352 169736
rect 283010 147792 283066 147801
rect 283010 147727 283066 147736
rect 282748 132466 282960 132494
rect 282748 132433 282776 132466
rect 282734 132424 282790 132433
rect 282734 132359 282790 132368
rect 282828 132388 282880 132394
rect 282828 132330 282880 132336
rect 282840 131753 282868 132330
rect 282826 131744 282882 131753
rect 282826 131679 282882 131688
rect 282274 130928 282330 130937
rect 282274 130863 282330 130872
rect 282288 130490 282316 130863
rect 282276 130484 282328 130490
rect 282276 130426 282328 130432
rect 282828 129260 282880 129266
rect 282828 129202 282880 129208
rect 282840 128625 282868 129202
rect 282826 128616 282882 128625
rect 282826 128551 282882 128560
rect 282828 126948 282880 126954
rect 282828 126890 282880 126896
rect 282840 126313 282868 126890
rect 282826 126304 282882 126313
rect 282826 126239 282882 126248
rect 282736 125588 282788 125594
rect 282736 125530 282788 125536
rect 282748 124817 282776 125530
rect 282828 125520 282880 125526
rect 282826 125488 282828 125497
rect 282880 125488 282882 125497
rect 282826 125423 282882 125432
rect 282734 124808 282790 124817
rect 282734 124743 282790 124752
rect 282182 123176 282238 123185
rect 282182 123111 282238 123120
rect 282092 122800 282144 122806
rect 282092 122742 282144 122748
rect 282104 122505 282132 122742
rect 282828 122732 282880 122738
rect 282828 122674 282880 122680
rect 282090 122496 282146 122505
rect 282090 122431 282146 122440
rect 282840 121689 282868 122674
rect 282826 121680 282882 121689
rect 282826 121615 282882 121624
rect 282736 121440 282788 121446
rect 282736 121382 282788 121388
rect 282748 120193 282776 121382
rect 282828 121372 282880 121378
rect 282828 121314 282880 121320
rect 282840 120873 282868 121314
rect 282826 120864 282882 120873
rect 282826 120799 282882 120808
rect 282734 120184 282790 120193
rect 282734 120119 282790 120128
rect 282828 120080 282880 120086
rect 282828 120022 282880 120028
rect 282840 119377 282868 120022
rect 282826 119368 282882 119377
rect 282826 119303 282882 119312
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 281908 118584 281960 118590
rect 281906 118552 281908 118561
rect 281960 118552 281962 118561
rect 281906 118487 281962 118496
rect 282840 117881 282868 118594
rect 284404 118590 284432 207674
rect 284484 184272 284536 184278
rect 284484 184214 284536 184220
rect 284496 153338 284524 184214
rect 284484 153332 284536 153338
rect 284484 153274 284536 153280
rect 284588 124030 284616 280162
rect 287152 273964 287204 273970
rect 287152 273906 287204 273912
rect 285680 262268 285732 262274
rect 285680 262210 285732 262216
rect 285692 143002 285720 262210
rect 285956 216028 286008 216034
rect 285956 215970 286008 215976
rect 285864 196716 285916 196722
rect 285864 196658 285916 196664
rect 285772 195356 285824 195362
rect 285772 195298 285824 195304
rect 285680 142996 285732 143002
rect 285680 142938 285732 142944
rect 285784 127974 285812 195298
rect 285876 130150 285904 196658
rect 285968 154222 285996 215970
rect 287060 177676 287112 177682
rect 287060 177618 287112 177624
rect 287072 171834 287100 177618
rect 287060 171828 287112 171834
rect 287060 171770 287112 171776
rect 285956 154216 286008 154222
rect 285956 154158 286008 154164
rect 287164 143750 287192 273906
rect 287244 220108 287296 220114
rect 287244 220050 287296 220056
rect 287152 143744 287204 143750
rect 287152 143686 287204 143692
rect 285864 130144 285916 130150
rect 285864 130086 285916 130092
rect 285772 127968 285824 127974
rect 285772 127910 285824 127916
rect 284576 124024 284628 124030
rect 284576 123966 284628 123972
rect 284392 118584 284444 118590
rect 284392 118526 284444 118532
rect 282826 117872 282882 117881
rect 282826 117807 282882 117816
rect 282184 117292 282236 117298
rect 282184 117234 282236 117240
rect 282196 116385 282224 117234
rect 282828 117224 282880 117230
rect 282828 117166 282880 117172
rect 282840 117065 282868 117166
rect 282826 117056 282882 117065
rect 282826 116991 282882 117000
rect 282182 116376 282238 116385
rect 282182 116311 282238 116320
rect 281724 115932 281776 115938
rect 281724 115874 281776 115880
rect 281736 114753 281764 115874
rect 282092 115864 282144 115870
rect 282092 115806 282144 115812
rect 282104 115569 282132 115806
rect 282090 115560 282146 115569
rect 282090 115495 282146 115504
rect 281722 114744 281778 114753
rect 281722 114679 281778 114688
rect 282276 114504 282328 114510
rect 282276 114446 282328 114452
rect 282288 114073 282316 114446
rect 282644 114436 282696 114442
rect 282644 114378 282696 114384
rect 282274 114064 282330 114073
rect 282274 113999 282330 114008
rect 282656 113257 282684 114378
rect 282642 113248 282698 113257
rect 282642 113183 282698 113192
rect 282092 113144 282144 113150
rect 282092 113086 282144 113092
rect 282104 112441 282132 113086
rect 282090 112432 282146 112441
rect 282090 112367 282146 112376
rect 282828 111784 282880 111790
rect 282828 111726 282880 111732
rect 282840 110945 282868 111726
rect 282826 110936 282882 110945
rect 282826 110871 282882 110880
rect 282828 110424 282880 110430
rect 282828 110366 282880 110372
rect 282840 109449 282868 110366
rect 282826 109440 282882 109449
rect 282826 109375 282882 109384
rect 282828 108996 282880 109002
rect 282828 108938 282880 108944
rect 282840 108633 282868 108938
rect 282826 108624 282882 108633
rect 282826 108559 282882 108568
rect 280250 107808 280306 107817
rect 280250 107743 280306 107752
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282840 105126 282868 105431
rect 287256 105126 287284 220050
rect 287348 140758 287376 288390
rect 288716 258120 288768 258126
rect 288716 258062 288768 258068
rect 288532 240168 288584 240174
rect 288532 240110 288584 240116
rect 288440 180328 288492 180334
rect 288440 180270 288492 180276
rect 288452 169930 288480 180270
rect 288440 169924 288492 169930
rect 288440 169866 288492 169872
rect 287336 140752 287388 140758
rect 287336 140694 287388 140700
rect 288544 129266 288572 240110
rect 288624 177608 288676 177614
rect 288624 177550 288676 177556
rect 288636 162926 288664 177550
rect 288624 162920 288676 162926
rect 288624 162862 288676 162868
rect 288728 130490 288756 258062
rect 289912 206304 289964 206310
rect 289912 206246 289964 206252
rect 289820 176112 289872 176118
rect 289820 176054 289872 176060
rect 289832 168366 289860 176054
rect 289820 168360 289872 168366
rect 289820 168302 289872 168308
rect 289924 165578 289952 206246
rect 290096 177336 290148 177342
rect 290096 177278 290148 177284
rect 290004 176044 290056 176050
rect 290004 175986 290056 175992
rect 289912 165572 289964 165578
rect 289912 165514 289964 165520
rect 290016 151706 290044 175986
rect 290004 151700 290056 151706
rect 290004 151642 290056 151648
rect 288716 130484 288768 130490
rect 288716 130426 288768 130432
rect 288532 129260 288584 129266
rect 288532 129202 288584 129208
rect 290108 125526 290136 177278
rect 290476 176050 290504 291178
rect 291844 260908 291896 260914
rect 291844 260850 291896 260856
rect 291200 199640 291252 199646
rect 291200 199582 291252 199588
rect 290464 176044 290516 176050
rect 290464 175986 290516 175992
rect 290096 125520 290148 125526
rect 290096 125462 290148 125468
rect 291212 110430 291240 199582
rect 291476 181552 291528 181558
rect 291476 181494 291528 181500
rect 291384 177472 291436 177478
rect 291290 177440 291346 177449
rect 291384 177414 291436 177420
rect 291290 177375 291346 177384
rect 291304 122738 291332 177375
rect 291396 150346 291424 177414
rect 291488 164218 291516 181494
rect 291856 177206 291884 260850
rect 292764 189780 292816 189786
rect 292764 189722 292816 189728
rect 292580 181756 292632 181762
rect 292580 181698 292632 181704
rect 291844 177200 291896 177206
rect 291844 177142 291896 177148
rect 291476 164212 291528 164218
rect 291476 164154 291528 164160
rect 291384 150340 291436 150346
rect 291384 150282 291436 150288
rect 291292 122732 291344 122738
rect 291292 122674 291344 122680
rect 292592 114442 292620 181698
rect 292672 177404 292724 177410
rect 292672 177346 292724 177352
rect 292684 136542 292712 177346
rect 292776 161362 292804 189722
rect 292856 176044 292908 176050
rect 292856 175986 292908 175992
rect 292868 162790 292896 175986
rect 292856 162784 292908 162790
rect 292856 162726 292908 162732
rect 292764 161356 292816 161362
rect 292764 161298 292816 161304
rect 292672 136536 292724 136542
rect 292672 136478 292724 136484
rect 292580 114436 292632 114442
rect 292580 114378 292632 114384
rect 291200 110424 291252 110430
rect 291200 110366 291252 110372
rect 282828 105120 282880 105126
rect 282828 105062 282880 105068
rect 287244 105120 287296 105126
rect 287244 105062 287296 105068
rect 281722 104816 281778 104825
rect 281722 104751 281778 104760
rect 280250 104000 280306 104009
rect 280250 103935 280306 103944
rect 280158 100872 280214 100881
rect 280158 100807 280214 100816
rect 279422 97336 279478 97345
rect 279422 97271 279478 97280
rect 279330 96656 279386 96665
rect 279330 96591 279386 96600
rect 268016 95940 268068 95946
rect 268016 95882 268068 95888
rect 267188 94512 267240 94518
rect 267188 94454 267240 94460
rect 268028 93838 268056 95882
rect 268016 93832 268068 93838
rect 268016 93774 268068 93780
rect 270972 93770 271000 96016
rect 276952 93838 276980 96016
rect 279344 95169 279372 96591
rect 279330 95160 279386 95169
rect 279330 95095 279386 95104
rect 279436 95062 279464 97271
rect 279424 95056 279476 95062
rect 279424 94998 279476 95004
rect 276940 93832 276992 93838
rect 276940 93774 276992 93780
rect 270960 93764 271012 93770
rect 270960 93706 271012 93712
rect 277400 93152 277452 93158
rect 277400 93094 277452 93100
rect 276020 91792 276072 91798
rect 276020 91734 276072 91740
rect 269120 73840 269172 73846
rect 269120 73782 269172 73788
rect 269132 16574 269160 73782
rect 273260 71052 273312 71058
rect 273260 70994 273312 71000
rect 271880 20052 271932 20058
rect 271880 19994 271932 20000
rect 271892 16574 271920 19994
rect 269132 16546 270080 16574
rect 271892 16546 272472 16574
rect 268384 14612 268436 14618
rect 268384 14554 268436 14560
rect 267004 3664 267056 3670
rect 267004 3606 267056 3612
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 267752 480 267780 3538
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 14554
rect 270052 480 270080 16546
rect 271236 9104 271288 9110
rect 271236 9046 271288 9052
rect 271248 480 271276 9046
rect 272444 480 272472 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 70994
rect 276032 3602 276060 91734
rect 277412 16574 277440 93094
rect 280172 86873 280200 100807
rect 280264 90982 280292 103935
rect 281630 102504 281686 102513
rect 281630 102439 281686 102448
rect 281538 100192 281594 100201
rect 281538 100127 281594 100136
rect 281552 95198 281580 100127
rect 281644 96422 281672 102439
rect 281632 96416 281684 96422
rect 281632 96358 281684 96364
rect 281540 95192 281592 95198
rect 281540 95134 281592 95140
rect 281736 95130 281764 104751
rect 281724 95124 281776 95130
rect 281724 95066 281776 95072
rect 280252 90976 280304 90982
rect 280252 90918 280304 90924
rect 280158 86864 280214 86873
rect 280158 86799 280214 86808
rect 287060 80708 287112 80714
rect 287060 80650 287112 80656
rect 281540 75200 281592 75206
rect 281540 75142 281592 75148
rect 280160 36576 280212 36582
rect 280160 36518 280212 36524
rect 280172 16574 280200 36518
rect 277412 16546 278360 16574
rect 280172 16546 280752 16574
rect 276112 16040 276164 16046
rect 276112 15982 276164 15988
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 15982
rect 276756 3596 276808 3602
rect 276756 3538 276808 3544
rect 274824 3460 274876 3466
rect 274824 3402 274876 3408
rect 276032 3454 276152 3482
rect 274836 480 274864 3402
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3538
rect 278332 480 278360 16546
rect 279514 3360 279570 3369
rect 279514 3295 279570 3304
rect 279528 480 279556 3295
rect 280724 480 280752 16546
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 354 281580 75142
rect 284392 22840 284444 22846
rect 284392 22782 284444 22788
rect 284404 6914 284432 22782
rect 285680 18760 285732 18766
rect 285680 18702 285732 18708
rect 285692 16574 285720 18702
rect 287072 16574 287100 80650
rect 293972 16574 294000 333202
rect 295340 267776 295392 267782
rect 295340 267718 295392 267724
rect 294052 198076 294104 198082
rect 294052 198018 294104 198024
rect 294064 135182 294092 198018
rect 294144 192500 294196 192506
rect 294144 192442 294196 192448
rect 294156 166326 294184 192442
rect 294236 175976 294288 175982
rect 294236 175918 294288 175924
rect 294144 166320 294196 166326
rect 294144 166262 294196 166268
rect 294248 162858 294276 175918
rect 294236 162852 294288 162858
rect 294236 162794 294288 162800
rect 294052 135176 294104 135182
rect 294052 135118 294104 135124
rect 295352 113150 295380 267718
rect 296720 257372 296772 257378
rect 296720 257314 296772 257320
rect 295432 214600 295484 214606
rect 295432 214542 295484 214548
rect 295444 167006 295472 214542
rect 295524 186992 295576 186998
rect 295524 186934 295576 186940
rect 295432 167000 295484 167006
rect 295432 166942 295484 166948
rect 295536 142050 295564 186934
rect 295616 177200 295668 177206
rect 295616 177142 295668 177148
rect 295524 142044 295576 142050
rect 295524 141986 295576 141992
rect 295628 137970 295656 177142
rect 295616 137964 295668 137970
rect 295616 137906 295668 137912
rect 295340 113144 295392 113150
rect 295340 113086 295392 113092
rect 296732 16574 296760 257314
rect 299480 239420 299532 239426
rect 299480 239362 299532 239368
rect 298098 225584 298154 225593
rect 298098 225519 298154 225528
rect 296904 199436 296956 199442
rect 296904 199378 296956 199384
rect 296812 180192 296864 180198
rect 296812 180134 296864 180140
rect 296824 118658 296852 180134
rect 296916 150414 296944 199378
rect 296996 193860 297048 193866
rect 296996 193802 297048 193808
rect 296904 150408 296956 150414
rect 296904 150350 296956 150356
rect 297008 146198 297036 193802
rect 296996 146192 297048 146198
rect 296996 146134 297048 146140
rect 296812 118652 296864 118658
rect 296812 118594 296864 118600
rect 298112 111790 298140 225519
rect 298190 196616 298246 196625
rect 298190 196551 298246 196560
rect 298204 144906 298232 196551
rect 298284 187060 298336 187066
rect 298284 187002 298336 187008
rect 298192 144900 298244 144906
rect 298192 144842 298244 144848
rect 298296 143478 298324 187002
rect 299388 178764 299440 178770
rect 299388 178706 299440 178712
rect 298744 178084 298796 178090
rect 298744 178026 298796 178032
rect 298284 143472 298336 143478
rect 298284 143414 298336 143420
rect 298756 115870 298784 178026
rect 299400 177970 299428 178706
rect 299492 178090 299520 239362
rect 299664 199504 299716 199510
rect 299664 199446 299716 199452
rect 299572 184340 299624 184346
rect 299572 184282 299624 184288
rect 299480 178084 299532 178090
rect 299480 178026 299532 178032
rect 299400 177942 299520 177970
rect 298744 115864 298796 115870
rect 298744 115806 298796 115812
rect 298100 111784 298152 111790
rect 298100 111726 298152 111732
rect 299492 16574 299520 177942
rect 299584 121378 299612 184282
rect 299676 151774 299704 199446
rect 299756 180260 299808 180266
rect 299756 180202 299808 180208
rect 299768 158710 299796 180202
rect 299756 158704 299808 158710
rect 299756 158646 299808 158652
rect 299664 151768 299716 151774
rect 299664 151710 299716 151716
rect 299572 121372 299624 121378
rect 299572 121314 299624 121320
rect 300872 16574 300900 384503
rect 302332 300892 302384 300898
rect 302332 300834 302384 300840
rect 302240 277432 302292 277438
rect 302240 277374 302292 277380
rect 300952 199572 301004 199578
rect 300952 199514 301004 199520
rect 300964 121446 300992 199514
rect 301044 181824 301096 181830
rect 301044 181766 301096 181772
rect 301056 157350 301084 181766
rect 301136 181484 301188 181490
rect 301136 181426 301188 181432
rect 301148 169726 301176 181426
rect 301136 169720 301188 169726
rect 301136 169662 301188 169668
rect 301044 157344 301096 157350
rect 301044 157286 301096 157292
rect 302252 126954 302280 277374
rect 302344 161430 302372 300834
rect 302424 210452 302476 210458
rect 302424 210394 302476 210400
rect 302332 161424 302384 161430
rect 302332 161366 302384 161372
rect 302240 126948 302292 126954
rect 302240 126890 302292 126896
rect 300952 121440 301004 121446
rect 300952 121382 301004 121388
rect 302436 115938 302464 210394
rect 302516 188488 302568 188494
rect 302516 188430 302568 188436
rect 302528 155922 302556 188430
rect 302516 155916 302568 155922
rect 302516 155858 302568 155864
rect 302424 115932 302476 115938
rect 302424 115874 302476 115880
rect 303632 16574 303660 385630
rect 303712 294024 303764 294030
rect 303712 293966 303764 293972
rect 303724 125594 303752 293966
rect 304998 292632 305054 292641
rect 304998 292567 305054 292576
rect 303804 229764 303856 229770
rect 303804 229706 303856 229712
rect 303712 125588 303764 125594
rect 303712 125530 303764 125536
rect 303816 114510 303844 229706
rect 303896 200796 303948 200802
rect 303896 200738 303948 200744
rect 303908 132394 303936 200738
rect 303896 132388 303948 132394
rect 303896 132330 303948 132336
rect 305012 122806 305040 292567
rect 305092 213240 305144 213246
rect 305092 213182 305144 213188
rect 305000 122800 305052 122806
rect 305000 122742 305052 122748
rect 305104 117230 305132 213182
rect 305184 202156 305236 202162
rect 305184 202098 305236 202104
rect 305196 147626 305224 202098
rect 305274 180024 305330 180033
rect 305274 179959 305330 179968
rect 305184 147620 305236 147626
rect 305184 147562 305236 147568
rect 305288 139330 305316 179959
rect 305276 139324 305328 139330
rect 305276 139266 305328 139272
rect 305092 117224 305144 117230
rect 305092 117166 305144 117172
rect 303804 114504 303856 114510
rect 303804 114446 303856 114452
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 299492 16546 299704 16574
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 284312 6886 284432 6914
rect 283104 6316 283156 6322
rect 283104 6258 283156 6264
rect 283116 480 283144 6258
rect 284312 480 284340 6886
rect 285404 3664 285456 3670
rect 285404 3606 285456 3612
rect 285416 480 285444 3606
rect 286612 480 286640 16546
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 292580 11824 292632 11830
rect 292580 11766 292632 11772
rect 290188 3528 290240 3534
rect 288990 3496 289046 3505
rect 290188 3470 290240 3476
rect 291382 3496 291438 3505
rect 288990 3431 289046 3440
rect 289004 480 289032 3431
rect 290200 480 290228 3470
rect 291382 3431 291438 3440
rect 291396 480 291424 3431
rect 292592 480 292620 11766
rect 293682 3496 293738 3505
rect 293682 3431 293738 3440
rect 293696 480 293724 3431
rect 294892 480 294920 16546
rect 296074 3496 296130 3505
rect 296074 3431 296130 3440
rect 296088 480 296116 3431
rect 297284 480 297312 16546
rect 298466 3904 298522 3913
rect 298466 3839 298522 3848
rect 298480 480 298508 3839
rect 299676 480 299704 16546
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 300780 480 300808 3431
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303158 3632 303214 3641
rect 303158 3567 303214 3576
rect 303172 480 303200 3567
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305550 3496 305606 3505
rect 305550 3431 305606 3440
rect 305564 480 305592 3431
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 386407
rect 309784 326392 309836 326398
rect 309784 326334 309836 326340
rect 309140 322244 309192 322250
rect 309140 322186 309192 322192
rect 307852 295384 307904 295390
rect 307852 295326 307904 295332
rect 306472 244316 306524 244322
rect 306472 244258 306524 244264
rect 306484 120086 306512 244258
rect 306564 236700 306616 236706
rect 306564 236642 306616 236648
rect 306576 143546 306604 236642
rect 306656 203584 306708 203590
rect 306656 203526 306708 203532
rect 306564 143540 306616 143546
rect 306564 143482 306616 143488
rect 306472 120080 306524 120086
rect 306472 120022 306524 120028
rect 306668 117298 306696 203526
rect 307760 181688 307812 181694
rect 307760 181630 307812 181636
rect 306656 117292 306708 117298
rect 306656 117234 306708 117240
rect 307772 882 307800 181630
rect 307864 139398 307892 295326
rect 307944 291848 307996 291854
rect 307944 291790 307996 291796
rect 307956 146266 307984 291790
rect 308036 185700 308088 185706
rect 308036 185642 308088 185648
rect 308048 153202 308076 185642
rect 308036 153196 308088 153202
rect 308036 153138 308088 153144
rect 307944 146260 307996 146266
rect 307944 146202 307996 146208
rect 307852 139392 307904 139398
rect 307852 139334 307904 139340
rect 309152 6914 309180 322186
rect 309232 302252 309284 302258
rect 309232 302194 309284 302200
rect 309244 136610 309272 302194
rect 309324 266416 309376 266422
rect 309324 266358 309376 266364
rect 309336 148986 309364 266358
rect 309324 148980 309376 148986
rect 309324 148922 309376 148928
rect 309232 136604 309284 136610
rect 309232 136546 309284 136552
rect 309796 16574 309824 326334
rect 311900 318164 311952 318170
rect 311900 318106 311952 318112
rect 310518 295352 310574 295361
rect 310518 295287 310574 295296
rect 310532 135250 310560 295287
rect 310704 264988 310756 264994
rect 310704 264930 310756 264936
rect 310612 248464 310664 248470
rect 310612 248406 310664 248412
rect 310520 135244 310572 135250
rect 310520 135186 310572 135192
rect 310624 109002 310652 248406
rect 310716 142118 310744 264930
rect 310704 142112 310756 142118
rect 310704 142054 310756 142060
rect 310612 108996 310664 109002
rect 310612 108938 310664 108944
rect 311912 16574 311940 318106
rect 313292 16574 313320 389127
rect 316038 366344 316094 366353
rect 316038 366279 316094 366288
rect 314660 349852 314712 349858
rect 314660 349794 314712 349800
rect 313372 233980 313424 233986
rect 313372 233922 313424 233928
rect 313384 133890 313412 233922
rect 313372 133884 313424 133890
rect 313372 133826 313424 133832
rect 309796 16546 309916 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309152 6886 309824 6914
rect 307942 3904 307998 3913
rect 307942 3839 307998 3848
rect 307760 876 307812 882
rect 307760 818 307812 824
rect 307956 480 307984 3839
rect 309048 876 309100 882
rect 309048 818 309100 824
rect 309060 480 309088 818
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 309888 3398 309916 16546
rect 309876 3392 309928 3398
rect 309876 3334 309928 3340
rect 311440 3392 311492 3398
rect 311440 3334 311492 3340
rect 311452 480 311480 3334
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 349794
rect 316052 3482 316080 366279
rect 316132 347064 316184 347070
rect 316132 347006 316184 347012
rect 316144 3602 316172 347006
rect 317432 16574 317460 395286
rect 349252 382968 349304 382974
rect 349252 382910 349304 382916
rect 318798 360904 318854 360913
rect 318798 360839 318854 360848
rect 318812 16574 318840 360839
rect 325700 356720 325752 356726
rect 325700 356662 325752 356668
rect 324412 354000 324464 354006
rect 324412 353942 324464 353948
rect 320180 316736 320232 316742
rect 320180 316678 320232 316684
rect 320192 16574 320220 316678
rect 322204 309800 322256 309806
rect 322204 309742 322256 309748
rect 321560 305652 321612 305658
rect 321560 305594 321612 305600
rect 321572 16574 321600 305594
rect 321652 244316 321704 244322
rect 321652 244258 321704 244264
rect 321664 242894 321692 244258
rect 321652 242888 321704 242894
rect 321652 242830 321704 242836
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316132 3596 316184 3602
rect 316132 3538 316184 3544
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 3538
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 322216 3058 322244 309742
rect 322938 300112 322994 300121
rect 322938 300047 322994 300056
rect 322204 3052 322256 3058
rect 322204 2994 322256 3000
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 300047
rect 324424 3534 324452 353942
rect 325712 16574 325740 356662
rect 331864 344344 331916 344350
rect 331864 344286 331916 344292
rect 328458 336016 328514 336025
rect 328458 335951 328514 335960
rect 327078 323640 327134 323649
rect 327078 323575 327134 323584
rect 327092 16574 327120 323575
rect 328472 16574 328500 335951
rect 331220 236768 331272 236774
rect 331220 236710 331272 236716
rect 329838 177304 329894 177313
rect 329838 177239 329894 177248
rect 329852 16574 329880 177239
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 324412 3052 324464 3058
rect 324412 2994 324464 3000
rect 324424 480 324452 2994
rect 325620 480 325648 3470
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 236710
rect 331876 3534 331904 344286
rect 338120 331900 338172 331906
rect 338120 331842 338172 331848
rect 336004 330540 336056 330546
rect 336004 330482 336056 330488
rect 333980 327140 334032 327146
rect 333980 327082 334032 327088
rect 332690 69592 332746 69601
rect 332690 69527 332746 69536
rect 332704 3670 332732 69527
rect 333992 16574 334020 327082
rect 335360 181620 335412 181626
rect 335360 181562 335412 181568
rect 335372 16574 335400 181562
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 3664 332744 3670
rect 332692 3606 332744 3612
rect 333888 3664 333940 3670
rect 333888 3606 333940 3612
rect 331864 3528 331916 3534
rect 331864 3470 331916 3476
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 332704 480 332732 3470
rect 333900 480 333928 3606
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335924 3482 335952 16546
rect 336016 3602 336044 330482
rect 336740 282192 336792 282198
rect 336740 282134 336792 282140
rect 336752 16574 336780 282134
rect 338132 16574 338160 331842
rect 342260 329112 342312 329118
rect 342260 329054 342312 329060
rect 339500 319456 339552 319462
rect 339500 319398 339552 319404
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 336004 3596 336056 3602
rect 336004 3538 336056 3544
rect 335924 3454 336320 3482
rect 336292 480 336320 3454
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 319398
rect 340878 283520 340934 283529
rect 340878 283455 340934 283464
rect 340892 3346 340920 283455
rect 340972 178696 341024 178702
rect 340972 178638 341024 178644
rect 340984 3534 341012 178638
rect 342272 16574 342300 329054
rect 345020 318096 345072 318102
rect 345020 318038 345072 318044
rect 343638 253192 343694 253201
rect 343638 253127 343694 253136
rect 343652 16574 343680 253127
rect 345032 16574 345060 318038
rect 346400 279472 346452 279478
rect 346400 279414 346452 279420
rect 346412 16574 346440 279414
rect 347780 278044 347832 278050
rect 347780 277986 347832 277992
rect 347792 16574 347820 277986
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 340892 3318 341012 3346
rect 340984 480 341012 3318
rect 342180 480 342208 3470
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349264 3534 349292 382910
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580354 365120 580410 365129
rect 580354 365055 580410 365064
rect 580264 365016 580316 365022
rect 580264 364958 580316 364964
rect 580276 351937 580304 364958
rect 580262 351928 580318 351937
rect 580262 351863 580318 351872
rect 580264 340944 580316 340950
rect 580264 340886 580316 340892
rect 352564 340196 352616 340202
rect 352564 340138 352616 340144
rect 350540 261520 350592 261526
rect 350540 261462 350592 261468
rect 350552 16574 350580 261462
rect 352576 193186 352604 340138
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 467104 287700 467156 287706
rect 467104 287642 467156 287648
rect 353944 260160 353996 260166
rect 353944 260102 353996 260108
rect 352564 193180 352616 193186
rect 352564 193122 352616 193128
rect 353956 167006 353984 260102
rect 358084 225004 358136 225010
rect 358084 224946 358136 224952
rect 353944 167000 353996 167006
rect 353944 166942 353996 166948
rect 358096 60722 358124 224946
rect 467116 126954 467144 287642
rect 468484 286340 468536 286346
rect 468484 286282 468536 286288
rect 468496 153202 468524 286282
rect 580276 272241 580304 340886
rect 580368 339454 580396 365055
rect 580356 339448 580408 339454
rect 580356 339390 580408 339396
rect 580354 325272 580410 325281
rect 580354 325207 580410 325216
rect 580368 315994 580396 325207
rect 580356 315988 580408 315994
rect 580356 315930 580408 315936
rect 582564 313336 582616 313342
rect 582564 313278 582616 313284
rect 582470 299568 582526 299577
rect 582470 299503 582526 299512
rect 580354 298752 580410 298761
rect 580354 298687 580410 298696
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 471244 269816 471296 269822
rect 471244 269758 471296 269764
rect 468484 153196 468536 153202
rect 468484 153138 468536 153144
rect 467104 126948 467156 126954
rect 467104 126890 467156 126896
rect 471256 100706 471284 269758
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580262 255912 580318 255921
rect 580262 255847 580318 255856
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580276 139369 580304 255847
rect 580368 246401 580396 298687
rect 582380 298172 582432 298178
rect 582380 298114 582432 298120
rect 580448 254584 580500 254590
rect 580448 254526 580500 254532
rect 580354 246392 580410 246401
rect 580354 246327 580410 246336
rect 580460 205737 580488 254526
rect 580540 247716 580592 247722
rect 580540 247658 580592 247664
rect 580552 232393 580580 247658
rect 580538 232384 580594 232393
rect 580538 232319 580594 232328
rect 580446 205728 580502 205737
rect 580446 205663 580502 205672
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 471244 100700 471296 100706
rect 471244 100642 471296 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 358084 60716 358136 60722
rect 358084 60658 358136 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 582392 19825 582420 298114
rect 582484 73001 582512 299503
rect 582576 219065 582604 313278
rect 582840 304292 582892 304298
rect 582840 304234 582892 304240
rect 582656 301504 582708 301510
rect 582656 301446 582708 301452
rect 582562 219056 582618 219065
rect 582562 218991 582618 219000
rect 582564 196648 582616 196654
rect 582564 196590 582616 196596
rect 582470 72992 582526 73001
rect 582470 72927 582526 72936
rect 582378 19816 582434 19825
rect 582378 19751 582434 19760
rect 350552 16546 351224 16574
rect 349252 3528 349304 3534
rect 349252 3470 349304 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 349264 480 349292 3334
rect 350460 480 350488 3470
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 582576 6633 582604 196590
rect 582668 112849 582696 301446
rect 582746 235240 582802 235249
rect 582746 235175 582802 235184
rect 582654 112840 582710 112849
rect 582654 112775 582710 112784
rect 582760 86193 582788 235175
rect 582852 179217 582880 304234
rect 582838 179208 582894 179217
rect 582838 179143 582894 179152
rect 582746 86184 582802 86193
rect 582746 86119 582802 86128
rect 582562 6624 582618 6633
rect 582562 6559 582618 6568
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3514 671200 3570 671256
rect 3514 658164 3570 658200
rect 3514 658144 3516 658164
rect 3516 658144 3568 658164
rect 3568 658144 3570 658164
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3238 579944 3294 580000
rect 3422 566888 3478 566944
rect 3146 553832 3202 553888
rect 3146 527856 3202 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3514 501744 3570 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 33046 474000 33102 474056
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3238 371320 3294 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3514 319232 3570 319288
rect 30286 375944 30342 376000
rect 3514 306176 3570 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 1398 24112 1454 24168
rect 3514 32408 3570 32464
rect 2870 25472 2926 25528
rect 3422 19352 3478 19408
rect 2962 6432 3018 6488
rect 13818 62736 13874 62792
rect 27618 51720 27674 51776
rect 19430 19896 19486 19952
rect 37094 439456 37150 439512
rect 38474 338000 38530 338056
rect 38658 40568 38714 40624
rect 42614 383152 42670 383208
rect 42798 30912 42854 30968
rect 48042 583752 48098 583808
rect 48962 433200 49018 433256
rect 48042 370504 48098 370560
rect 48042 340720 48098 340776
rect 49330 431840 49386 431896
rect 49330 430616 49386 430672
rect 49606 355272 49662 355328
rect 52090 494844 52092 494864
rect 52092 494844 52144 494864
rect 52144 494844 52146 494864
rect 52090 494808 52146 494844
rect 52090 492632 52146 492688
rect 49514 222808 49570 222864
rect 53286 491952 53342 492008
rect 53838 583888 53894 583944
rect 55862 584024 55918 584080
rect 56506 584024 56562 584080
rect 55034 583888 55090 583944
rect 53470 387504 53526 387560
rect 59082 538736 59138 538792
rect 56414 253816 56470 253872
rect 57794 186904 57850 186960
rect 61382 463528 61438 463584
rect 61382 462304 61438 462360
rect 60738 442856 60794 442912
rect 67638 581324 67694 581360
rect 67638 581304 67640 581324
rect 67640 581304 67692 581324
rect 67692 581304 67694 581324
rect 67914 580624 67970 580680
rect 67362 579128 67418 579184
rect 61382 337900 61384 337920
rect 61384 337900 61436 337920
rect 61436 337900 61438 337920
rect 61382 337864 61438 337900
rect 63222 467744 63278 467800
rect 62026 401648 62082 401704
rect 63314 447752 63370 447808
rect 64602 477400 64658 477456
rect 60922 253816 60978 253872
rect 63130 196696 63186 196752
rect 60646 93608 60702 93664
rect 62026 89664 62082 89720
rect 56598 73752 56654 73808
rect 53930 24792 53986 24848
rect 55126 24792 55182 24848
rect 53930 24112 53986 24168
rect 63498 355308 63500 355328
rect 63500 355308 63552 355328
rect 63552 355308 63554 355328
rect 63498 355272 63554 355308
rect 63498 72392 63554 72448
rect 64786 398792 64842 398848
rect 67178 568656 67234 568712
rect 66074 461352 66130 461408
rect 66074 460944 66130 461000
rect 65982 440292 66038 440328
rect 65982 440272 65984 440292
rect 65984 440272 66036 440292
rect 66036 440272 66038 440292
rect 67638 578448 67694 578504
rect 67638 577768 67694 577824
rect 67638 575728 67694 575784
rect 67730 575048 67786 575104
rect 67638 574368 67694 574424
rect 67730 573416 67786 573472
rect 67638 572756 67694 572792
rect 67638 572736 67640 572756
rect 67640 572736 67692 572756
rect 67692 572736 67694 572756
rect 68558 580624 68614 580680
rect 68650 571784 68706 571840
rect 68282 571648 68338 571704
rect 68466 571648 68522 571704
rect 67638 570016 67694 570072
rect 67638 568928 67694 568984
rect 67546 567568 67602 567624
rect 67362 480528 67418 480584
rect 67270 459448 67326 459504
rect 66994 451868 66996 451888
rect 66996 451868 67048 451888
rect 67048 451868 67050 451888
rect 66994 451832 67050 451868
rect 67638 567196 67640 567216
rect 67640 567196 67692 567216
rect 67692 567196 67694 567216
rect 67638 567160 67694 567196
rect 67638 564848 67694 564904
rect 67730 564476 67732 564496
rect 67732 564476 67784 564496
rect 67784 564476 67786 564496
rect 67730 564440 67786 564476
rect 67730 564168 67786 564224
rect 67638 563624 67694 563680
rect 67638 562980 67640 563000
rect 67640 562980 67692 563000
rect 67692 562980 67694 563000
rect 67638 562944 67694 562980
rect 67638 560360 67694 560416
rect 67638 559408 67694 559464
rect 68374 558864 68430 558920
rect 67638 557540 67640 557560
rect 67640 557540 67692 557560
rect 67692 557540 67694 557560
rect 67638 557504 67694 557540
rect 67730 556688 67786 556744
rect 67638 556180 67640 556200
rect 67640 556180 67692 556200
rect 67692 556180 67694 556200
rect 67638 556144 67694 556180
rect 67638 555328 67694 555384
rect 67730 554784 67786 554840
rect 67638 553444 67694 553480
rect 67638 553424 67640 553444
rect 67640 553424 67692 553444
rect 67692 553424 67694 553444
rect 67638 552084 67694 552120
rect 67638 552064 67640 552084
rect 67640 552064 67692 552084
rect 67692 552064 67694 552084
rect 67638 551248 67694 551304
rect 68282 550704 68338 550760
rect 67730 549888 67786 549944
rect 67638 549364 67694 549400
rect 67638 549344 67640 549364
rect 67640 549344 67692 549364
rect 67692 549344 67694 549364
rect 67638 548528 67694 548584
rect 67730 547168 67786 547224
rect 67638 546508 67694 546544
rect 67638 546488 67640 546508
rect 67640 546488 67692 546508
rect 67692 546488 67694 546508
rect 67730 544448 67786 544504
rect 67638 543788 67694 543824
rect 67638 543768 67640 543788
rect 67640 543768 67692 543788
rect 67692 543768 67694 543788
rect 67638 542544 67694 542600
rect 67638 541184 67694 541240
rect 67638 540096 67694 540152
rect 67730 488008 67786 488064
rect 67638 487872 67694 487928
rect 67638 485852 67694 485888
rect 67638 485832 67640 485852
rect 67640 485832 67692 485852
rect 67692 485832 67694 485852
rect 67638 485152 67694 485208
rect 67638 483656 67694 483712
rect 68098 482432 68154 482488
rect 67638 480140 67694 480176
rect 67638 480120 67640 480140
rect 67640 480120 67692 480140
rect 67692 480120 67694 480140
rect 67730 479848 67786 479904
rect 67730 477400 67786 477456
rect 67638 476312 67694 476368
rect 67730 476176 67786 476232
rect 67638 475632 67694 475688
rect 67638 474988 67640 475008
rect 67640 474988 67692 475008
rect 67692 474988 67694 475008
rect 67638 474952 67694 474988
rect 67638 474308 67640 474328
rect 67640 474308 67692 474328
rect 67692 474308 67694 474328
rect 67638 474272 67694 474308
rect 67638 472232 67694 472288
rect 67638 470872 67694 470928
rect 67730 470328 67786 470384
rect 67638 469648 67694 469704
rect 67638 468968 67694 469024
rect 67638 468172 67694 468208
rect 67638 468152 67640 468172
rect 67640 468152 67692 468172
rect 67692 468152 67694 468172
rect 67638 465568 67694 465624
rect 67638 465452 67694 465488
rect 67638 465432 67640 465452
rect 67640 465432 67692 465452
rect 67692 465432 67694 465452
rect 67638 464752 67694 464808
rect 67730 464208 67786 464264
rect 67638 462848 67694 462904
rect 67638 460672 67694 460728
rect 67730 460164 67732 460184
rect 67732 460164 67784 460184
rect 67784 460164 67786 460184
rect 67730 460128 67786 460164
rect 67638 458768 67694 458824
rect 68098 457952 68154 458008
rect 67638 457444 67640 457464
rect 67640 457444 67692 457464
rect 67692 457444 67694 457464
rect 67638 457408 67694 457444
rect 67638 455912 67694 455968
rect 67638 454552 67694 454608
rect 67730 453872 67786 453928
rect 67638 453192 67694 453248
rect 68834 576408 68890 576464
rect 68742 545808 68798 545864
rect 68742 484628 68798 484664
rect 68742 484608 68744 484628
rect 68744 484608 68796 484628
rect 68796 484608 68798 484628
rect 68558 481072 68614 481128
rect 68926 543224 68982 543280
rect 71778 583888 71834 583944
rect 69110 558864 69166 558920
rect 69110 553968 69166 554024
rect 68926 541728 68982 541784
rect 68374 476992 68430 477048
rect 68834 476992 68890 477048
rect 67730 451288 67786 451344
rect 67638 449948 67694 449984
rect 67638 449928 67640 449948
rect 67640 449928 67692 449948
rect 67692 449928 67694 449948
rect 67730 449268 67786 449304
rect 67730 449248 67732 449268
rect 67732 449248 67784 449268
rect 67784 449248 67786 449268
rect 68282 449248 68338 449304
rect 67638 449148 67640 449168
rect 67640 449148 67692 449168
rect 67692 449148 67694 449168
rect 67638 449112 67694 449148
rect 67638 447208 67694 447264
rect 67638 446392 67694 446448
rect 67730 445848 67786 445904
rect 67638 445052 67694 445088
rect 67638 445032 67640 445052
rect 67640 445032 67692 445052
rect 67692 445032 67694 445052
rect 67730 444216 67786 444272
rect 67638 443808 67694 443864
rect 67730 442856 67786 442912
rect 67638 442448 67694 442504
rect 67730 441632 67786 441688
rect 67730 441088 67786 441144
rect 67454 379888 67510 379944
rect 67638 440272 67694 440328
rect 67638 439456 67694 439512
rect 67730 382472 67786 382528
rect 67638 382064 67694 382120
rect 67638 380724 67694 380760
rect 67638 380704 67640 380724
rect 67640 380704 67692 380724
rect 67692 380704 67694 380724
rect 68006 380296 68062 380352
rect 67638 378256 67694 378312
rect 67638 377304 67694 377360
rect 67638 375128 67694 375184
rect 67730 374176 67786 374232
rect 67638 372408 67694 372464
rect 67638 371456 67694 371512
rect 67730 369164 67786 369200
rect 67730 369144 67732 369164
rect 67732 369144 67784 369164
rect 67784 369144 67786 369164
rect 67638 369008 67694 369064
rect 67638 367124 67694 367160
rect 67638 367104 67640 367124
rect 67640 367104 67692 367124
rect 67692 367104 67694 367124
rect 67638 366424 67694 366480
rect 67730 366288 67786 366344
rect 67638 363724 67694 363760
rect 67638 363704 67640 363724
rect 67640 363704 67692 363724
rect 67692 363704 67694 363724
rect 67730 363604 67732 363624
rect 67732 363604 67784 363624
rect 67784 363604 67786 363624
rect 67730 363568 67786 363604
rect 67638 362072 67694 362128
rect 67638 360984 67694 361040
rect 67638 359508 67694 359544
rect 67638 359488 67640 359508
rect 67640 359488 67692 359508
rect 67692 359488 67694 359508
rect 67730 358128 67786 358184
rect 67638 358028 67640 358048
rect 67640 358028 67692 358048
rect 67692 358028 67694 358048
rect 67638 357992 67694 358028
rect 67638 355544 67694 355600
rect 67730 355408 67786 355464
rect 67638 353776 67694 353832
rect 67638 352552 67694 352608
rect 67914 352416 67970 352472
rect 68926 468968 68982 469024
rect 68834 385736 68890 385792
rect 68742 383424 68798 383480
rect 74630 584296 74686 584352
rect 83186 586336 83242 586392
rect 84382 583888 84438 583944
rect 84474 583752 84530 583808
rect 91006 584024 91062 584080
rect 92846 582392 92902 582448
rect 97906 583752 97962 583808
rect 102598 581712 102654 581768
rect 69202 486512 69258 486568
rect 107106 583888 107162 583944
rect 106738 583752 106794 583808
rect 107106 578856 107162 578912
rect 106462 578040 106518 578096
rect 106370 574640 106426 574696
rect 106278 560360 106334 560416
rect 106186 552064 106242 552120
rect 105818 543768 105874 543824
rect 70398 532208 70454 532264
rect 69754 489912 69810 489968
rect 74538 531936 74594 531992
rect 76562 537512 76618 537568
rect 76470 532072 76526 532128
rect 77758 495488 77814 495544
rect 81622 537376 81678 537432
rect 80886 490456 80942 490512
rect 84842 490048 84898 490104
rect 89350 537376 89406 537432
rect 90638 494672 90694 494728
rect 92018 490592 92074 490648
rect 92846 491544 92902 491600
rect 97906 536016 97962 536072
rect 95146 490456 95202 490512
rect 97814 491408 97870 491464
rect 99378 536832 99434 536888
rect 99286 491272 99342 491328
rect 99286 489232 99342 489288
rect 69846 489096 69902 489152
rect 69294 482568 69350 482624
rect 69386 482432 69442 482488
rect 69202 457952 69258 458008
rect 69110 454008 69166 454064
rect 68926 372816 68982 372872
rect 68374 365064 68430 365120
rect 99470 476312 99526 476368
rect 99378 446528 99434 446584
rect 99286 442448 99342 442504
rect 69846 441224 69902 441280
rect 99286 441088 99342 441144
rect 71042 438912 71098 438968
rect 70674 437688 70730 437744
rect 79322 440680 79378 440736
rect 81438 440680 81494 440736
rect 71778 431840 71834 431896
rect 71042 387776 71098 387832
rect 74538 434560 74594 434616
rect 73526 387776 73582 387832
rect 77942 439456 77998 439512
rect 78678 437552 78734 437608
rect 76010 387640 76066 387696
rect 79690 438776 79746 438832
rect 79690 437552 79746 437608
rect 81898 437416 81954 437472
rect 84198 438912 84254 438968
rect 81530 391176 81586 391232
rect 84198 399608 84254 399664
rect 85118 399472 85174 399528
rect 85946 386416 86002 386472
rect 91282 438776 91338 438832
rect 90362 438640 90418 438696
rect 89626 435920 89682 435976
rect 92570 439048 92626 439104
rect 93674 404912 93730 404968
rect 93766 399472 93822 399528
rect 92478 397976 92534 398032
rect 91558 390632 91614 390688
rect 91926 390632 91982 390688
rect 95882 389136 95938 389192
rect 96526 389816 96582 389872
rect 96526 389136 96582 389192
rect 100114 489912 100170 489968
rect 100114 488280 100170 488336
rect 99746 443672 99802 443728
rect 102046 537920 102102 537976
rect 100942 536968 100998 537024
rect 102046 536968 102102 537024
rect 101862 489932 101918 489968
rect 101862 489912 101864 489932
rect 101864 489912 101916 489932
rect 101916 489912 101918 489932
rect 100666 476312 100722 476368
rect 100298 441088 100354 441144
rect 100850 451152 100906 451208
rect 100758 439728 100814 439784
rect 99194 392536 99250 392592
rect 98826 388320 98882 388376
rect 101954 478896 102010 478952
rect 103426 487872 103482 487928
rect 103334 487328 103390 487384
rect 103426 486648 103482 486704
rect 102322 485288 102378 485344
rect 102322 483792 102378 483848
rect 102322 482876 102324 482896
rect 102324 482876 102376 482896
rect 102376 482876 102378 482896
rect 102322 482840 102378 482876
rect 102414 482568 102470 482624
rect 102322 481516 102324 481536
rect 102324 481516 102376 481536
rect 102376 481516 102378 481536
rect 102322 481480 102378 481516
rect 102414 481208 102470 481264
rect 102322 479848 102378 479904
rect 103426 478080 103482 478136
rect 102414 477808 102470 477864
rect 102506 476992 102562 477048
rect 102322 476448 102378 476504
rect 102322 475632 102378 475688
rect 102414 475088 102470 475144
rect 102322 474272 102378 474328
rect 102506 474000 102562 474056
rect 102322 472912 102378 472968
rect 103426 472368 103482 472424
rect 102322 471688 102378 471744
rect 103426 471144 103482 471200
rect 102414 471008 102470 471064
rect 103426 470192 103482 470248
rect 102782 469648 102838 469704
rect 102322 468832 102378 468888
rect 102782 466928 102838 466984
rect 103426 466792 103482 466848
rect 102322 466112 102378 466168
rect 103426 465704 103482 465760
rect 103426 465432 103482 465488
rect 102414 464752 102470 464808
rect 102322 464208 102378 464264
rect 102322 463392 102378 463448
rect 102322 462032 102378 462088
rect 102322 461352 102378 461408
rect 102874 460128 102930 460184
rect 102322 459992 102378 460048
rect 102322 459312 102378 459368
rect 102414 458632 102470 458688
rect 102230 456048 102286 456104
rect 102230 454688 102286 454744
rect 102230 453872 102286 453928
rect 102230 453192 102286 453248
rect 102230 452548 102232 452568
rect 102232 452548 102284 452568
rect 102284 452548 102286 452568
rect 102230 452512 102286 452548
rect 102138 449268 102194 449304
rect 102138 449248 102140 449268
rect 102140 449248 102192 449268
rect 102192 449248 102194 449268
rect 102138 448468 102140 448488
rect 102140 448468 102192 448488
rect 102192 448468 102194 448488
rect 102138 448432 102194 448468
rect 102138 446256 102194 446312
rect 102046 441768 102102 441824
rect 102046 440136 102102 440192
rect 102046 438912 102102 438968
rect 100758 393352 100814 393408
rect 102414 456592 102470 456648
rect 102414 449112 102470 449168
rect 102414 447888 102470 447944
rect 102598 443672 102654 443728
rect 102874 442992 102930 443048
rect 103334 441768 103390 441824
rect 102874 441088 102930 441144
rect 103058 439728 103114 439784
rect 103518 458088 103574 458144
rect 103518 455368 103574 455424
rect 104806 538056 104862 538112
rect 104714 537784 104770 537840
rect 105542 536832 105598 536888
rect 104254 491544 104310 491600
rect 103518 450608 103574 450664
rect 104070 445712 104126 445768
rect 104070 445168 104126 445224
rect 104162 444352 104218 444408
rect 103518 444216 103574 444272
rect 103426 394032 103482 394088
rect 106094 540368 106150 540424
rect 109130 582392 109186 582448
rect 108946 580760 109002 580816
rect 108854 580080 108910 580136
rect 108854 579400 108910 579456
rect 108946 578720 109002 578776
rect 108210 577496 108266 577552
rect 108854 576680 108910 576736
rect 108946 576000 109002 576056
rect 108946 573996 108948 574016
rect 108948 573996 109000 574016
rect 109000 573996 109002 574016
rect 108946 573960 109002 573996
rect 107658 573280 107714 573336
rect 107842 573280 107898 573336
rect 108946 572736 109002 572792
rect 108946 571920 109002 571976
rect 107934 571376 107990 571432
rect 107750 563080 107806 563136
rect 107658 560380 107714 560416
rect 107658 560360 107660 560380
rect 107660 560360 107712 560380
rect 107712 560360 107714 560380
rect 107658 556280 107714 556336
rect 106922 551520 106978 551576
rect 107658 542680 107714 542736
rect 107566 540096 107622 540152
rect 106462 486512 106518 486568
rect 106094 456728 106150 456784
rect 107566 456048 107622 456104
rect 107842 548800 107898 548856
rect 108854 570560 108910 570616
rect 108946 570016 109002 570072
rect 108946 569200 109002 569256
rect 108946 567840 109002 567896
rect 108946 567196 108948 567216
rect 108948 567196 109000 567216
rect 109000 567196 109002 567216
rect 108946 567160 109002 567196
rect 108854 566480 108910 566536
rect 108946 565836 108948 565856
rect 108948 565836 109000 565856
rect 109000 565836 109002 565856
rect 108946 565800 109002 565836
rect 108946 565120 109002 565176
rect 108946 563780 109002 563816
rect 108946 563760 108948 563780
rect 108948 563760 109000 563780
rect 109000 563760 109002 563780
rect 108946 561040 109002 561096
rect 108854 559680 108910 559736
rect 108946 559000 109002 559056
rect 108578 558320 108634 558376
rect 108946 556960 109002 557016
rect 108946 554240 109002 554296
rect 108946 553560 109002 553616
rect 108946 552880 109002 552936
rect 108946 550840 109002 550896
rect 108854 550160 108910 550216
rect 108946 549480 109002 549536
rect 108946 547440 109002 547496
rect 108946 546080 109002 546136
rect 108946 545400 109002 545456
rect 108946 544720 109002 544776
rect 108946 543360 109002 543416
rect 108946 542000 109002 542056
rect 109222 555736 109278 555792
rect 109774 537920 109830 537976
rect 109130 488280 109186 488336
rect 109130 467880 109186 467936
rect 110326 490456 110382 490512
rect 111706 578196 111762 578232
rect 111706 578176 111708 578196
rect 111708 578176 111760 578196
rect 111760 578176 111762 578196
rect 111798 537784 111854 537840
rect 110418 393932 110420 393952
rect 110420 393932 110472 393952
rect 110472 393932 110474 393952
rect 110418 393896 110474 393932
rect 111982 466248 112038 466304
rect 112166 485052 112168 485072
rect 112168 485052 112220 485072
rect 112220 485052 112222 485072
rect 112166 485016 112222 485052
rect 113086 485016 113142 485072
rect 114466 488688 114522 488744
rect 113822 401240 113878 401296
rect 114650 459720 114706 459776
rect 116030 477400 116086 477456
rect 115938 475940 115940 475960
rect 115940 475940 115992 475960
rect 115992 475940 115994 475960
rect 115938 475904 115994 475940
rect 115202 458244 115258 458280
rect 115202 458224 115204 458244
rect 115204 458224 115256 458244
rect 115256 458224 115258 458244
rect 114926 389136 114982 389192
rect 69202 360848 69258 360904
rect 69110 356904 69166 356960
rect 69478 356904 69534 356960
rect 68742 352416 68798 352472
rect 67730 351464 67786 351520
rect 68282 351464 68338 351520
rect 67638 349832 67694 349888
rect 68006 349696 68062 349752
rect 68558 347112 68614 347168
rect 67638 346704 67694 346760
rect 67730 345616 67786 345672
rect 67730 344392 67786 344448
rect 67638 343712 67694 343768
rect 67638 341672 67694 341728
rect 67546 341536 67602 341592
rect 68650 334736 68706 334792
rect 68926 349696 68982 349752
rect 68834 348372 68836 348392
rect 68836 348372 68888 348392
rect 68888 348372 68890 348392
rect 68834 348336 68890 348372
rect 68742 333240 68798 333296
rect 66166 320728 66222 320784
rect 67638 291080 67694 291136
rect 68190 289448 68246 289504
rect 67638 288088 67694 288144
rect 66902 287408 66958 287464
rect 68282 286456 68338 286512
rect 67638 284416 67694 284472
rect 67730 283328 67786 283384
rect 67638 282104 67694 282160
rect 67638 280336 67694 280392
rect 67730 279928 67786 279984
rect 67638 279248 67694 279304
rect 67730 277752 67786 277808
rect 67638 277616 67694 277672
rect 67638 276392 67694 276448
rect 67822 275032 67878 275088
rect 67638 274896 67694 274952
rect 67730 274488 67786 274544
rect 67638 273536 67694 273592
rect 67638 272176 67694 272232
rect 67546 271904 67602 271960
rect 66074 227024 66130 227080
rect 67362 182824 67418 182880
rect 67638 270952 67694 271008
rect 67730 270816 67786 270872
rect 67730 269592 67786 269648
rect 67638 269456 67694 269512
rect 67638 268096 67694 268152
rect 67638 267416 67694 267472
rect 67730 267008 67786 267064
rect 67638 264968 67694 265024
rect 67638 264868 67640 264888
rect 67640 264868 67692 264888
rect 67692 264868 67694 264888
rect 67638 264832 67694 264868
rect 67730 263628 67786 263664
rect 67730 263608 67732 263628
rect 67732 263608 67784 263628
rect 67784 263608 67786 263628
rect 67638 263508 67640 263528
rect 67640 263508 67692 263528
rect 67692 263508 67694 263528
rect 67638 263472 67694 263508
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67638 261432 67694 261488
rect 67730 260908 67786 260944
rect 67730 260888 67732 260908
rect 67732 260888 67784 260908
rect 67784 260888 67786 260908
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 259528 67694 259584
rect 67730 258576 67786 258632
rect 67638 258188 67694 258224
rect 67638 258168 67640 258188
rect 67640 258168 67692 258188
rect 67692 258168 67694 258188
rect 67638 257896 67694 257952
rect 67638 256808 67694 256864
rect 67730 255332 67786 255368
rect 67730 255312 67732 255332
rect 67732 255312 67784 255332
rect 67784 255312 67786 255332
rect 67638 255212 67640 255232
rect 67640 255212 67692 255232
rect 67692 255212 67694 255232
rect 67638 255176 67694 255212
rect 67730 253972 67786 254008
rect 67730 253952 67732 253972
rect 67732 253952 67784 253972
rect 67784 253952 67786 253972
rect 67638 253852 67640 253872
rect 67640 253852 67692 253872
rect 67692 253852 67694 253872
rect 67638 253816 67694 253852
rect 67638 252612 67694 252648
rect 67638 252592 67640 252612
rect 67640 252592 67692 252612
rect 67692 252592 67694 252612
rect 67730 249872 67786 249928
rect 67638 249756 67694 249792
rect 67638 249736 67640 249756
rect 67640 249736 67692 249756
rect 67692 249736 67694 249756
rect 67638 247696 67694 247752
rect 67730 247152 67786 247208
rect 67638 246608 67694 246664
rect 67638 245248 67694 245304
rect 67638 244568 67694 244624
rect 115938 460128 115994 460184
rect 115938 459720 115994 459776
rect 117318 484336 117374 484392
rect 116122 384240 116178 384296
rect 116674 384240 116730 384296
rect 116122 383560 116178 383616
rect 116766 383596 116768 383616
rect 116768 383596 116820 383616
rect 116820 383596 116822 383616
rect 116766 383560 116822 383596
rect 116030 370232 116086 370288
rect 115938 353232 115994 353288
rect 115294 349152 115350 349208
rect 71134 339904 71190 339960
rect 71318 338000 71374 338056
rect 71318 337456 71374 337512
rect 72974 334600 73030 334656
rect 70030 298152 70086 298208
rect 69018 296792 69074 296848
rect 68742 293936 68798 293992
rect 68926 292712 68982 292768
rect 68834 290808 68890 290864
rect 68742 286048 68798 286104
rect 68650 285368 68706 285424
rect 71042 292304 71098 292360
rect 73158 302776 73214 302832
rect 75826 339360 75882 339416
rect 79046 339632 79102 339688
rect 76654 315288 76710 315344
rect 79046 337320 79102 337376
rect 78678 331744 78734 331800
rect 76562 295976 76618 296032
rect 84842 337456 84898 337512
rect 82082 322088 82138 322144
rect 89074 333920 89130 333976
rect 92386 306992 92442 307048
rect 90638 298288 90694 298344
rect 96526 331064 96582 331120
rect 95238 330656 95294 330712
rect 96526 330656 96582 330712
rect 94594 304136 94650 304192
rect 96526 300056 96582 300112
rect 95790 294072 95846 294128
rect 99010 292576 99066 292632
rect 111062 330384 111118 330440
rect 107566 296112 107622 296168
rect 111062 297336 111118 297392
rect 113178 300736 113234 300792
rect 114466 300736 114522 300792
rect 114466 299512 114522 299568
rect 115386 339496 115442 339552
rect 117502 461488 117558 461544
rect 117502 459584 117558 459640
rect 117318 385328 117374 385384
rect 117502 384920 117558 384976
rect 117318 382220 117374 382256
rect 117318 382200 117320 382220
rect 117320 382200 117372 382220
rect 117372 382200 117374 382220
rect 117318 380860 117374 380896
rect 117318 380840 117320 380860
rect 117320 380840 117372 380860
rect 117372 380840 117374 380860
rect 116674 359760 116730 359816
rect 115294 305632 115350 305688
rect 115846 295296 115902 295352
rect 115294 294208 115350 294264
rect 115754 294208 115810 294264
rect 114282 291896 114338 291952
rect 117502 373380 117558 373416
rect 117502 373360 117504 373380
rect 117504 373360 117556 373380
rect 117556 373360 117558 373380
rect 118238 384940 118294 384976
rect 118238 384920 118240 384940
rect 118240 384920 118292 384940
rect 118292 384920 118294 384940
rect 117686 379480 117742 379536
rect 118606 378820 118662 378856
rect 118606 378800 118608 378820
rect 118608 378800 118660 378820
rect 118660 378800 118662 378820
rect 118606 376760 118662 376816
rect 118606 376100 118662 376136
rect 119986 494944 120042 495000
rect 120170 488416 120226 488472
rect 118790 378120 118846 378176
rect 118606 376080 118608 376100
rect 118608 376080 118660 376100
rect 118660 376080 118662 376100
rect 118514 375400 118570 375456
rect 118606 374040 118662 374096
rect 118422 372680 118478 372736
rect 118606 371320 118662 371376
rect 118514 367920 118570 367976
rect 118606 367260 118662 367296
rect 118606 367240 118608 367260
rect 118608 367240 118660 367260
rect 118660 367240 118662 367260
rect 118606 365880 118662 365936
rect 118606 365200 118662 365256
rect 118606 364520 118662 364576
rect 117594 363568 117650 363624
rect 117962 362480 118018 362536
rect 118606 361800 118662 361856
rect 118606 361120 118662 361176
rect 118146 359080 118202 359136
rect 118606 358436 118608 358456
rect 118608 358436 118660 358456
rect 118660 358436 118662 358456
rect 118606 358400 118662 358436
rect 117686 357060 117742 357096
rect 117686 357040 117688 357060
rect 117688 357040 117740 357060
rect 117740 357040 117742 357060
rect 118606 355680 118662 355736
rect 118054 354320 118110 354376
rect 118606 353640 118662 353696
rect 117962 352960 118018 353016
rect 117410 351600 117466 351656
rect 117318 350920 117374 350976
rect 117778 348880 117834 348936
rect 117410 347520 117466 347576
rect 117778 340040 117834 340096
rect 118514 351600 118570 351656
rect 118422 350920 118478 350976
rect 118606 350240 118662 350296
rect 118606 348200 118662 348256
rect 118330 346160 118386 346216
rect 118606 345480 118662 345536
rect 118606 344800 118662 344856
rect 118146 343440 118202 343496
rect 118606 342760 118662 342816
rect 118606 342080 118662 342136
rect 118054 340720 118110 340776
rect 119342 377304 119398 377360
rect 118882 369960 118938 370016
rect 118974 368600 119030 368656
rect 119986 356088 120042 356144
rect 120354 442448 120410 442504
rect 120262 380976 120318 381032
rect 121642 463528 121698 463584
rect 121550 439320 121606 439376
rect 122102 439320 122158 439376
rect 123114 489912 123170 489968
rect 121918 388864 121974 388920
rect 120630 387776 120686 387832
rect 122102 387776 122158 387832
rect 122102 385192 122158 385248
rect 120446 337456 120502 337512
rect 118606 292848 118662 292904
rect 119802 289856 119858 289912
rect 69018 289720 69074 289776
rect 68926 284008 68982 284064
rect 68374 280472 68430 280528
rect 69110 268232 69166 268288
rect 68834 251776 68890 251832
rect 69018 245656 69074 245712
rect 67822 244160 67878 244216
rect 67730 243888 67786 243944
rect 67638 242528 67694 242584
rect 67638 241848 67694 241904
rect 67638 240488 67694 240544
rect 120170 292848 120226 292904
rect 120078 256400 120134 256456
rect 69294 255856 69350 255912
rect 120078 250960 120134 251016
rect 119986 240896 120042 240952
rect 75826 238584 75882 238640
rect 75918 228248 75974 228304
rect 74538 197920 74594 197976
rect 78678 192480 78734 192536
rect 77298 189624 77354 189680
rect 86222 238448 86278 238504
rect 84382 226888 84438 226944
rect 87050 208936 87106 208992
rect 91926 238448 91982 238504
rect 99470 213152 99526 213208
rect 103518 238720 103574 238776
rect 104806 238720 104862 238776
rect 67454 179968 67510 180024
rect 97722 177656 97778 177712
rect 99286 177656 99342 177712
rect 101954 177656 102010 177712
rect 110142 179424 110198 179480
rect 104806 177656 104862 177712
rect 110142 176976 110198 177032
rect 100666 176704 100722 176760
rect 102046 176704 102102 176760
rect 103334 176704 103390 176760
rect 105726 176704 105782 176760
rect 107014 176704 107070 176760
rect 108118 176724 108174 176760
rect 108118 176704 108120 176724
rect 108120 176704 108172 176724
rect 108172 176704 108174 176724
rect 122102 367648 122158 367704
rect 121642 314200 121698 314256
rect 121642 291760 121698 291816
rect 121642 290400 121698 290456
rect 121734 289040 121790 289096
rect 121826 288360 121882 288416
rect 121642 287680 121698 287736
rect 121642 287000 121698 287056
rect 121550 286320 121606 286376
rect 121734 285640 121790 285696
rect 121642 284960 121698 285016
rect 121550 284688 121606 284744
rect 121550 283600 121606 283656
rect 121550 282940 121606 282976
rect 121550 282920 121552 282940
rect 121552 282920 121604 282940
rect 121604 282920 121606 282940
rect 121642 282240 121698 282296
rect 121550 281580 121606 281616
rect 121550 281560 121552 281580
rect 121552 281560 121604 281580
rect 121604 281560 121606 281580
rect 121550 280880 121606 280936
rect 121642 279520 121698 279576
rect 121550 278860 121606 278896
rect 121550 278840 121552 278860
rect 121552 278840 121604 278860
rect 121604 278840 121606 278860
rect 121642 278160 121698 278216
rect 121550 277500 121606 277536
rect 121550 277480 121552 277500
rect 121552 277480 121604 277500
rect 121604 277480 121606 277500
rect 121550 276800 121606 276856
rect 121734 276120 121790 276176
rect 121550 274760 121606 274816
rect 121642 274080 121698 274136
rect 121826 275440 121882 275496
rect 121550 273400 121606 273456
rect 121642 272720 121698 272776
rect 121550 272040 121606 272096
rect 121550 271360 121606 271416
rect 121550 270000 121606 270056
rect 121642 269320 121698 269376
rect 121550 268640 121606 268696
rect 121550 267960 121606 268016
rect 121734 267280 121790 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121458 264560 121514 264616
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121550 261160 121606 261216
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 121550 259120 121606 259176
rect 121458 258440 121514 258496
rect 121550 257760 121606 257816
rect 120722 257080 120778 257136
rect 121458 255720 121514 255776
rect 121550 255040 121606 255096
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121734 261840 121790 261896
rect 121642 252320 121698 252376
rect 121458 251640 121514 251696
rect 121550 250280 121606 250336
rect 121458 249600 121514 249656
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 121458 246200 121514 246256
rect 121550 245520 121606 245576
rect 120170 244840 120226 244896
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121550 242120 121606 242176
rect 122286 375944 122342 376000
rect 122746 247560 122802 247616
rect 123022 388864 123078 388920
rect 124218 392536 124274 392592
rect 123850 369008 123906 369064
rect 122930 250960 122986 251016
rect 122102 241440 122158 241496
rect 121458 240760 121514 240816
rect 122378 240080 122434 240136
rect 124310 324284 124366 324320
rect 124310 324264 124312 324284
rect 124312 324264 124364 324284
rect 124364 324264 124366 324284
rect 127254 460128 127310 460184
rect 125782 332424 125838 332480
rect 129830 484336 129886 484392
rect 128450 338000 128506 338056
rect 127070 296112 127126 296168
rect 131118 485016 131174 485072
rect 129830 328380 129832 328400
rect 129832 328380 129884 328400
rect 129884 328380 129886 328400
rect 129830 328344 129886 328380
rect 129922 297336 129978 297392
rect 132498 477400 132554 477456
rect 129830 240896 129886 240952
rect 133142 329740 133144 329760
rect 133144 329740 133196 329760
rect 133196 329740 133198 329760
rect 133142 329704 133198 329740
rect 133786 329024 133842 329080
rect 135350 474000 135406 474056
rect 135442 457408 135498 457464
rect 133970 323720 134026 323776
rect 134614 385600 134670 385656
rect 348790 702480 348846 702536
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580262 630808 580318 630864
rect 580170 617480 580226 617536
rect 140870 341400 140926 341456
rect 138018 238584 138074 238640
rect 133878 226244 133880 226264
rect 133880 226244 133932 226264
rect 133932 226244 133934 226264
rect 133878 226208 133934 226244
rect 580170 590960 580226 591016
rect 579802 577632 579858 577688
rect 580170 564304 580226 564360
rect 580906 537784 580962 537840
rect 579802 524456 579858 524512
rect 580170 511264 580226 511320
rect 151818 471144 151874 471200
rect 149058 456048 149114 456104
rect 150438 457408 150494 457464
rect 580170 471416 580226 471472
rect 580354 484608 580410 484664
rect 580262 458088 580318 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 160742 401648 160798 401704
rect 153106 362208 153162 362264
rect 141422 190984 141478 191040
rect 114098 177656 114154 177712
rect 114466 177656 114522 177712
rect 118422 177656 118478 177712
rect 119986 177656 120042 177712
rect 122654 177656 122710 177712
rect 128266 177656 128322 177712
rect 129462 177656 129518 177712
rect 126794 176976 126850 177032
rect 133142 176976 133198 177032
rect 115846 176704 115902 176760
rect 123758 176704 123814 176760
rect 128174 176704 128230 176760
rect 130750 176704 130806 176760
rect 132406 176704 132462 176760
rect 134798 176704 134854 176760
rect 264242 400288 264298 400344
rect 164882 291896 164938 291952
rect 164882 181328 164938 181384
rect 160742 177384 160798 177440
rect 136086 176740 136088 176760
rect 136088 176740 136140 176760
rect 136140 176740 136142 176760
rect 136086 176704 136142 176740
rect 148230 176704 148286 176760
rect 116950 175480 117006 175536
rect 120814 175480 120870 175536
rect 124494 175480 124550 175536
rect 158902 175480 158958 175536
rect 110694 175344 110750 175400
rect 167550 171536 167606 171592
rect 169666 168408 169722 168464
rect 67454 129240 67510 129296
rect 66166 128016 66222 128072
rect 65522 125160 65578 125216
rect 66074 123528 66130 123584
rect 66074 122576 66130 122632
rect 67362 120808 67418 120864
rect 66166 94832 66222 94888
rect 66074 91024 66130 91080
rect 67546 126248 67602 126304
rect 67454 93744 67510 93800
rect 67638 102312 67694 102368
rect 67730 100680 67786 100736
rect 94962 94696 95018 94752
rect 104346 94696 104402 94752
rect 116674 94696 116730 94752
rect 120630 94696 120686 94752
rect 133142 94696 133198 94752
rect 151726 94696 151782 94752
rect 85670 93472 85726 93528
rect 107750 93472 107806 93528
rect 115846 93472 115902 93528
rect 122102 93472 122158 93528
rect 103426 93200 103482 93256
rect 110234 93200 110290 93256
rect 85118 92384 85174 92440
rect 88062 92384 88118 92440
rect 99286 92384 99342 92440
rect 100022 92384 100078 92440
rect 75826 91160 75882 91216
rect 86866 91160 86922 91216
rect 99102 91296 99158 91352
rect 89074 91160 89130 91216
rect 90638 91160 90694 91216
rect 91926 91160 91982 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97078 91160 97134 91216
rect 97906 91160 97962 91216
rect 97078 88168 97134 88224
rect 101862 91704 101918 91760
rect 99194 91160 99250 91216
rect 100574 91160 100630 91216
rect 101954 91296 102010 91352
rect 102046 91160 102102 91216
rect 103334 91160 103390 91216
rect 101954 84088 102010 84144
rect 105726 92404 105782 92440
rect 105726 92384 105728 92404
rect 105728 92384 105780 92404
rect 105780 92384 105782 92404
rect 106830 92384 106886 92440
rect 109682 92248 109738 92304
rect 104806 91160 104862 91216
rect 105726 91160 105782 91216
rect 102046 78512 102102 78568
rect 107106 91160 107162 91216
rect 108762 91160 108818 91216
rect 108762 86672 108818 86728
rect 114466 92420 114468 92440
rect 114468 92420 114520 92440
rect 114520 92420 114522 92440
rect 114466 92384 114522 92420
rect 120262 92384 120318 92440
rect 123206 92384 123262 92440
rect 124126 92384 124182 92440
rect 125414 92384 125470 92440
rect 112718 91568 112774 91624
rect 119526 91568 119582 91624
rect 110326 91160 110382 91216
rect 111062 91160 111118 91216
rect 111706 91160 111762 91216
rect 114466 91296 114522 91352
rect 115846 91296 115902 91352
rect 113086 91160 113142 91216
rect 114374 91160 114430 91216
rect 114374 83952 114430 84008
rect 115754 91160 115810 91216
rect 117226 91160 117282 91216
rect 118238 91160 118294 91216
rect 122838 91432 122894 91488
rect 119710 91160 119766 91216
rect 122286 91160 122342 91216
rect 134430 92384 134486 92440
rect 151542 92384 151598 92440
rect 152094 92384 152150 92440
rect 126886 91704 126942 91760
rect 126794 91296 126850 91352
rect 125506 91160 125562 91216
rect 126702 91160 126758 91216
rect 136270 91568 136326 91624
rect 128266 91160 128322 91216
rect 129462 91160 129518 91216
rect 130750 91160 130806 91216
rect 132406 91160 132462 91216
rect 132406 86536 132462 86592
rect 151726 91160 151782 91216
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 168194 110064 168250 110120
rect 167918 108704 167974 108760
rect 171782 187040 171838 187096
rect 115846 77152 115902 77208
rect 70398 24112 70454 24168
rect 92478 64096 92534 64152
rect 98642 43424 98698 43480
rect 117318 11600 117374 11656
rect 178682 294072 178738 294128
rect 178682 95104 178738 95160
rect 185582 296792 185638 296848
rect 181442 177248 181498 177304
rect 185582 94968 185638 95024
rect 189722 181328 189778 181384
rect 193862 177384 193918 177440
rect 196714 93472 196770 93528
rect 202234 175888 202290 175944
rect 204994 119312 205050 119368
rect 206466 177384 206522 177440
rect 206466 93608 206522 93664
rect 210606 94832 210662 94888
rect 211894 89664 211950 89720
rect 213274 166096 213330 166152
rect 213826 175752 213882 175808
rect 213918 175108 213920 175128
rect 213920 175108 213972 175128
rect 213972 175108 213974 175128
rect 213918 175072 213974 175108
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214102 173304 214158 173360
rect 213918 172352 213974 172408
rect 214010 171944 214066 172000
rect 214010 170720 214066 170776
rect 214010 169652 214066 169688
rect 214010 169632 214012 169652
rect 214012 169632 214064 169652
rect 214064 169632 214066 169652
rect 213918 169360 213974 169416
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 214010 168000 214066 168056
rect 213918 166932 213974 166968
rect 213918 166912 213920 166932
rect 213920 166912 213972 166932
rect 213972 166912 213974 166932
rect 214010 166640 214066 166696
rect 213918 165280 213974 165336
rect 213458 164736 213514 164792
rect 213918 163920 213974 163976
rect 213918 162560 213974 162616
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 215114 171128 215170 171184
rect 214562 160792 214618 160848
rect 213918 160012 213920 160032
rect 213920 160012 213972 160032
rect 213972 160012 213974 160032
rect 213918 159976 213974 160012
rect 214010 159432 214066 159488
rect 214102 158616 214158 158672
rect 213918 157276 213974 157312
rect 213918 157256 213920 157276
rect 213920 157256 213972 157276
rect 213972 157256 213974 157276
rect 214010 156848 214066 156904
rect 215022 158072 215078 158128
rect 214838 155896 214894 155952
rect 213918 155488 213974 155544
rect 214010 153856 214066 153912
rect 213918 153332 213974 153368
rect 213918 153312 213920 153332
rect 213920 153312 213972 153332
rect 213972 153312 213974 153332
rect 213918 152632 213974 152688
rect 213918 151952 213974 152008
rect 214654 151816 214710 151872
rect 213918 150864 213974 150920
rect 214470 150728 214526 150784
rect 214010 150184 214066 150240
rect 213918 148688 213974 148744
rect 213918 148008 213974 148064
rect 214010 146648 214066 146704
rect 213918 146376 213974 146432
rect 213918 144916 213920 144936
rect 213920 144916 213972 144936
rect 213972 144916 213974 144936
rect 213918 144880 213974 144916
rect 213918 143928 213974 143984
rect 213274 143520 213330 143576
rect 214010 142704 214066 142760
rect 213918 142296 213974 142352
rect 214010 141344 214066 141400
rect 213918 140936 213974 140992
rect 214930 149504 214986 149560
rect 213918 139984 213974 140040
rect 214010 139440 214066 139496
rect 213918 138760 213974 138816
rect 214654 138080 214710 138136
rect 213918 137400 213974 137456
rect 214010 135632 214066 135688
rect 213918 135360 213974 135416
rect 214010 134272 214066 134328
rect 213918 134000 213974 134056
rect 214562 132504 214618 132560
rect 214010 131416 214066 131472
rect 213918 131164 213974 131200
rect 213918 131144 213920 131164
rect 213920 131144 213972 131164
rect 213972 131144 213974 131164
rect 213918 130056 213974 130112
rect 213918 128424 213974 128480
rect 213918 127472 213974 127528
rect 214010 126112 214066 126168
rect 213918 125704 213974 125760
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 122868 213974 122904
rect 213918 122848 213920 122868
rect 213920 122848 213972 122868
rect 213972 122848 213974 122868
rect 214010 122168 214066 122224
rect 213918 121508 213974 121544
rect 213918 121488 213920 121508
rect 213920 121488 213972 121508
rect 213972 121488 213974 121508
rect 214010 120808 214066 120864
rect 213918 120148 213974 120184
rect 213918 120128 213920 120148
rect 213920 120128 213972 120148
rect 213972 120128 213974 120148
rect 214010 119584 214066 119640
rect 213366 119040 213422 119096
rect 213918 118904 213974 118960
rect 213918 117544 213974 117600
rect 214010 117272 214066 117328
rect 214010 116184 214066 116240
rect 213918 115948 213920 115968
rect 213920 115948 213972 115968
rect 213972 115948 213974 115968
rect 213918 115912 213974 115948
rect 213918 114960 213974 115016
rect 213458 114552 213514 114608
rect 214010 113600 214066 113656
rect 213918 113228 213920 113248
rect 213920 113228 213972 113248
rect 213972 113228 213974 113248
rect 213918 113192 213974 113228
rect 214010 112240 214066 112296
rect 213918 111852 213974 111888
rect 213918 111832 213920 111852
rect 213920 111832 213972 111852
rect 213972 111832 213974 111852
rect 214010 110880 214066 110936
rect 213918 110492 213974 110528
rect 213918 110472 213920 110492
rect 213920 110472 213972 110492
rect 213972 110472 213974 110492
rect 214010 109656 214066 109712
rect 213918 109132 213974 109168
rect 213918 109112 213920 109132
rect 213920 109112 213972 109132
rect 213972 109112 213974 109132
rect 214010 108296 214066 108352
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106528 213974 106584
rect 213918 105712 213974 105768
rect 214010 105168 214066 105224
rect 213918 103672 213974 103728
rect 213918 102448 213974 102504
rect 214010 101088 214066 101144
rect 213918 100816 213974 100872
rect 213918 99728 213974 99784
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 214746 117952 214802 118008
rect 214654 103808 214710 103864
rect 214838 99456 214894 99512
rect 214746 96600 214802 96656
rect 216218 97008 216274 97064
rect 216678 95784 216734 95840
rect 238022 392536 238078 392592
rect 227074 177520 227130 177576
rect 227718 175752 227774 175808
rect 229098 174664 229154 174720
rect 229190 172352 229246 172408
rect 229282 171400 229338 171456
rect 229374 168544 229430 168600
rect 231766 173712 231822 173768
rect 231122 173304 231178 173360
rect 231490 172760 231546 172816
rect 231766 171808 231822 171864
rect 230754 169532 230756 169552
rect 230756 169532 230808 169552
rect 230808 169532 230810 169552
rect 230754 169496 230810 169532
rect 230570 158616 230626 158672
rect 230478 157664 230534 157720
rect 231122 170448 231178 170504
rect 231766 170856 231822 170912
rect 231490 169904 231546 169960
rect 231490 168952 231546 169008
rect 231766 168000 231822 168056
rect 231766 167048 231822 167104
rect 231674 166096 231730 166152
rect 231766 165688 231822 165744
rect 231766 165144 231822 165200
rect 231674 164736 231730 164792
rect 231122 164328 231178 164384
rect 231766 163784 231822 163840
rect 231674 163376 231730 163432
rect 231122 162832 231178 162888
rect 231766 162460 231768 162480
rect 231768 162460 231820 162480
rect 231820 162460 231822 162480
rect 231766 162424 231822 162460
rect 231674 161880 231730 161936
rect 231030 161472 231086 161528
rect 231766 160928 231822 160984
rect 231674 160520 231730 160576
rect 231766 160012 231768 160032
rect 231768 160012 231820 160032
rect 231820 160012 231822 160032
rect 231766 159976 231822 160012
rect 231674 159568 231730 159624
rect 231674 159024 231730 159080
rect 231490 158752 231546 158808
rect 230938 156168 230994 156224
rect 230570 155796 230572 155816
rect 230572 155796 230624 155816
rect 230624 155796 230626 155816
rect 230570 155760 230626 155796
rect 230938 155216 230994 155272
rect 230754 152904 230810 152960
rect 229834 151000 229890 151056
rect 230938 150048 230994 150104
rect 231030 149640 231086 149696
rect 230754 147192 230810 147248
rect 230938 146784 230994 146840
rect 230754 143928 230810 143984
rect 230478 142432 230534 142488
rect 229742 142024 229798 142080
rect 230938 140120 230994 140176
rect 229098 96620 229154 96656
rect 229098 96600 229100 96620
rect 229100 96600 229152 96620
rect 229152 96600 229154 96620
rect 230754 134000 230810 134056
rect 231030 132504 231086 132560
rect 230754 132096 230810 132152
rect 230754 127880 230810 127936
rect 230938 122168 230994 122224
rect 230662 118904 230718 118960
rect 231398 153856 231454 153912
rect 231306 153348 231308 153368
rect 231308 153348 231360 153368
rect 231360 153348 231362 153368
rect 231306 153312 231362 153348
rect 231122 117408 231178 117464
rect 230662 117000 230718 117056
rect 231306 149096 231362 149152
rect 231766 157120 231822 157176
rect 231674 156712 231730 156768
rect 231766 154300 231768 154320
rect 231768 154300 231820 154320
rect 231820 154300 231822 154320
rect 231766 154264 231822 154300
rect 231674 152496 231730 152552
rect 231766 151952 231822 152008
rect 232042 166640 232098 166696
rect 231766 151544 231822 151600
rect 231674 150592 231730 150648
rect 231766 148144 231822 148200
rect 231490 146240 231546 146296
rect 231766 145832 231822 145888
rect 231674 145288 231730 145344
rect 232686 153176 232742 153232
rect 231674 144880 231730 144936
rect 231766 144336 231822 144392
rect 231766 143384 231822 143440
rect 231766 140684 231822 140720
rect 231766 140664 231768 140684
rect 231768 140664 231820 140684
rect 231820 140664 231822 140684
rect 231490 139712 231546 139768
rect 231674 139204 231676 139224
rect 231676 139204 231728 139224
rect 231728 139204 231730 139224
rect 231674 139168 231730 139204
rect 231766 138760 231822 138816
rect 231766 137264 231822 137320
rect 231490 136856 231546 136912
rect 231766 136312 231822 136368
rect 231674 135904 231730 135960
rect 231582 135768 231638 135824
rect 231398 135360 231454 135416
rect 231306 133728 231362 133784
rect 231490 131552 231546 131608
rect 231490 130192 231546 130248
rect 231398 129784 231454 129840
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231766 133456 231822 133512
rect 231674 133048 231730 133104
rect 231766 131144 231822 131200
rect 231766 130600 231822 130656
rect 231766 129240 231822 129296
rect 231674 128832 231730 128888
rect 231766 128288 231822 128344
rect 231674 127336 231730 127392
rect 231582 126928 231638 126984
rect 231766 126384 231822 126440
rect 231306 125296 231362 125352
rect 231490 124480 231546 124536
rect 231306 120672 231362 120728
rect 231306 119312 231362 119368
rect 231766 125024 231822 125080
rect 231766 124108 231768 124128
rect 231768 124108 231820 124128
rect 231820 124108 231822 124128
rect 231766 124072 231822 124108
rect 231582 123120 231638 123176
rect 231766 122576 231822 122632
rect 231490 121624 231546 121680
rect 231766 121216 231822 121272
rect 231490 120264 231546 120320
rect 231766 119720 231822 119776
rect 231214 116048 231270 116104
rect 231214 115096 231270 115152
rect 231122 114552 231178 114608
rect 231398 117952 231454 118008
rect 231306 113600 231362 113656
rect 230938 110744 230994 110800
rect 230570 107888 230626 107944
rect 230754 106528 230810 106584
rect 230570 104216 230626 104272
rect 231490 116456 231546 116512
rect 231766 114144 231822 114200
rect 231490 113192 231546 113248
rect 231674 112648 231730 112704
rect 231766 112240 231822 112296
rect 231674 111716 231730 111752
rect 231674 111696 231676 111716
rect 231676 111696 231728 111716
rect 231728 111696 231730 111716
rect 231766 111288 231822 111344
rect 231766 110356 231822 110392
rect 231766 110336 231768 110356
rect 231768 110336 231820 110356
rect 231820 110336 231822 110356
rect 231674 109792 231730 109848
rect 231674 109384 231730 109440
rect 231766 108876 231768 108896
rect 231768 108876 231820 108896
rect 231820 108876 231822 108896
rect 231766 108840 231822 108876
rect 231674 108432 231730 108488
rect 231490 107108 231492 107128
rect 231492 107108 231544 107128
rect 231544 107108 231546 107128
rect 231490 107072 231546 107108
rect 231490 105168 231546 105224
rect 231398 104624 231454 104680
rect 231766 107480 231822 107536
rect 231766 105576 231822 105632
rect 231582 103672 231638 103728
rect 231122 103264 231178 103320
rect 230478 102720 230534 102776
rect 230754 101360 230810 101416
rect 230570 100816 230626 100872
rect 231490 99864 231546 99920
rect 231490 98504 231546 98560
rect 230938 97960 230994 98016
rect 231674 100408 231730 100464
rect 231766 99456 231822 99512
rect 231766 99048 231822 99104
rect 231582 97552 231638 97608
rect 231766 97008 231822 97064
rect 230478 95648 230534 95704
rect 238022 178608 238078 178664
rect 238758 168272 238814 168328
rect 238298 146104 238354 146160
rect 240506 3440 240562 3496
rect 245198 3440 245254 3496
rect 246394 3440 246450 3496
rect 248786 3440 248842 3496
rect 249982 3440 250038 3496
rect 253478 126248 253534 126304
rect 252374 3440 252430 3496
rect 253478 3440 253534 3496
rect 259458 180104 259514 180160
rect 258722 177248 258778 177304
rect 261482 174392 261538 174448
rect 261298 130736 261354 130792
rect 261206 98912 261262 98968
rect 261574 100544 261630 100600
rect 265622 177384 265678 177440
rect 264426 175752 264482 175808
rect 265714 174936 265770 174992
rect 265806 174120 265862 174176
rect 265898 173168 265954 173224
rect 265530 172760 265586 172816
rect 265714 172488 265770 172544
rect 265622 171536 265678 171592
rect 265438 170584 265494 170640
rect 265254 170176 265310 170232
rect 265622 169788 265678 169824
rect 265622 169768 265624 169788
rect 265624 169768 265676 169788
rect 265676 169768 265678 169788
rect 265346 168952 265402 169008
rect 265622 168544 265678 168600
rect 265254 168408 265310 168464
rect 264426 166776 264482 166832
rect 265346 167592 265402 167648
rect 265898 171944 265954 172000
rect 265806 171164 265808 171184
rect 265808 171164 265860 171184
rect 265860 171164 265862 171184
rect 265806 171128 265862 171164
rect 265806 169360 265862 169416
rect 265346 165960 265402 166016
rect 265346 165008 265402 165064
rect 265162 164600 265218 164656
rect 265162 164192 265218 164248
rect 264242 163784 264298 163840
rect 262954 141344 263010 141400
rect 257066 4800 257122 4856
rect 255870 3440 255926 3496
rect 259458 3440 259514 3496
rect 258262 3304 258318 3360
rect 265714 166368 265770 166424
rect 265806 165724 265808 165744
rect 265808 165724 265860 165744
rect 265860 165724 265862 165744
rect 265806 165688 265862 165724
rect 265806 163376 265862 163432
rect 264518 162424 264574 162480
rect 264426 161880 264482 161936
rect 265530 162968 265586 163024
rect 265530 161608 265586 161664
rect 265990 160792 266046 160848
rect 265898 160384 265954 160440
rect 265806 160148 265808 160168
rect 265808 160148 265860 160168
rect 265860 160148 265862 160168
rect 265806 160112 265862 160148
rect 265622 159840 265678 159896
rect 265530 159432 265586 159488
rect 265070 157392 265126 157448
rect 265346 153856 265402 153912
rect 264334 152632 264390 152688
rect 264242 133048 264298 133104
rect 264242 119040 264298 119096
rect 265254 152088 265310 152144
rect 265438 150864 265494 150920
rect 265346 149640 265402 149696
rect 265438 149096 265494 149152
rect 265530 148688 265586 148744
rect 265070 147872 265126 147928
rect 265530 146648 265586 146704
rect 265438 146104 265494 146160
rect 264978 143112 265034 143168
rect 265530 144472 265586 144528
rect 265438 142840 265494 142896
rect 265346 142704 265402 142760
rect 265254 142160 265310 142216
rect 264426 140528 264482 140584
rect 264426 133728 264482 133784
rect 264426 130600 264482 130656
rect 264426 128152 264482 128208
rect 264426 126792 264482 126848
rect 264426 122576 264482 122632
rect 264426 121216 264482 121272
rect 264426 117272 264482 117328
rect 264426 111288 264482 111344
rect 264334 101904 264390 101960
rect 264518 107480 264574 107536
rect 264518 107072 264574 107128
rect 265162 138100 265218 138136
rect 265162 138080 265164 138100
rect 265164 138080 265216 138100
rect 265216 138080 265218 138100
rect 265530 140936 265586 140992
rect 265806 158752 265862 158808
rect 265990 158208 266046 158264
rect 265806 157800 265862 157856
rect 265898 156848 265954 156904
rect 265806 156032 265862 156088
rect 266082 156440 266138 156496
rect 265714 155624 265770 155680
rect 265990 155216 266046 155272
rect 265806 154808 265862 154864
rect 265898 154672 265954 154728
rect 265806 153448 265862 153504
rect 265898 153176 265954 153232
rect 265806 151852 265808 151872
rect 265808 151852 265860 151872
rect 265860 151852 265862 151872
rect 265806 151816 265862 151852
rect 265714 151272 265770 151328
rect 265806 150492 265808 150512
rect 265808 150492 265860 150512
rect 265860 150492 265862 150512
rect 265806 150456 265862 150492
rect 265806 150048 265862 150104
rect 266082 152360 266138 152416
rect 265714 148280 265770 148336
rect 265898 147056 265954 147112
rect 265990 146512 266046 146568
rect 265806 145696 265862 145752
rect 265714 145288 265770 145344
rect 265898 144880 265954 144936
rect 265806 143520 265862 143576
rect 265806 142296 265862 142352
rect 265898 141344 265954 141400
rect 265714 139712 265770 139768
rect 265806 139476 265808 139496
rect 265808 139476 265860 139496
rect 265860 139476 265862 139496
rect 265806 139440 265862 139476
rect 265806 138352 265862 138408
rect 265162 135224 265218 135280
rect 265254 134544 265310 134600
rect 265806 137536 265862 137592
rect 265714 137128 265770 137184
rect 265806 135380 265862 135416
rect 265806 135360 265808 135380
rect 265808 135360 265860 135380
rect 265860 135360 265862 135380
rect 265806 134136 265862 134192
rect 265622 132776 265678 132832
rect 265714 131960 265770 132016
rect 265622 131144 265678 131200
rect 265346 128968 265402 129024
rect 265806 128560 265862 128616
rect 265346 127608 265402 127664
rect 265806 126384 265862 126440
rect 265622 125976 265678 126032
rect 265714 125568 265770 125624
rect 266082 136720 266138 136776
rect 265990 136312 266046 136368
rect 265530 124208 265586 124264
rect 265806 125024 265862 125080
rect 265898 124616 265954 124672
rect 265898 123392 265954 123448
rect 265806 122984 265862 123040
rect 265898 122032 265954 122088
rect 265806 121624 265862 121680
rect 265990 120808 266046 120864
rect 265898 120400 265954 120456
rect 265806 120128 265862 120184
rect 265622 119448 265678 119504
rect 265530 118804 265532 118824
rect 265532 118804 265584 118824
rect 265584 118804 265586 118824
rect 265530 118768 265586 118804
rect 265162 118224 265218 118280
rect 265530 116864 265586 116920
rect 265622 116456 265678 116512
rect 265622 115232 265678 115288
rect 265438 114824 265494 114880
rect 265530 113872 265586 113928
rect 265438 113464 265494 113520
rect 265530 112648 265586 112704
rect 265622 112240 265678 112296
rect 265162 110880 265218 110936
rect 265530 110064 265586 110120
rect 265346 108296 265402 108352
rect 265254 105712 265310 105768
rect 265622 104916 265678 104952
rect 265622 104896 265624 104916
rect 265624 104896 265676 104916
rect 265676 104896 265678 104916
rect 265622 104488 265678 104544
rect 265530 103128 265586 103184
rect 265346 102332 265402 102368
rect 265346 102312 265348 102332
rect 265348 102312 265400 102332
rect 265400 102312 265402 102332
rect 265622 102720 265678 102776
rect 265162 99728 265218 99784
rect 265622 99476 265678 99512
rect 265622 99456 265624 99476
rect 265624 99456 265676 99476
rect 265676 99456 265678 99476
rect 264610 98776 264666 98832
rect 265622 97552 265678 97608
rect 265346 97144 265402 97200
rect 265530 95648 265586 95704
rect 265990 117816 266046 117872
rect 265898 117428 265954 117464
rect 265898 117408 265900 117428
rect 265900 117408 265952 117428
rect 265952 117408 265954 117428
rect 266082 116048 266138 116104
rect 265898 113212 265954 113248
rect 265898 113192 265900 113212
rect 265900 113192 265952 113212
rect 265952 113192 265954 113212
rect 265898 112104 265954 112160
rect 265898 110472 265954 110528
rect 265990 109656 266046 109712
rect 265898 109132 265954 109168
rect 265898 109112 265900 109132
rect 265900 109112 265952 109132
rect 265952 109112 265954 109132
rect 265990 108704 266046 108760
rect 265898 107908 265954 107944
rect 265898 107888 265900 107908
rect 265900 107888 265952 107908
rect 265952 107888 265954 107908
rect 265990 106664 266046 106720
rect 265898 106528 265954 106584
rect 265898 105304 265954 105360
rect 265990 103944 266046 104000
rect 265898 103556 265954 103592
rect 265898 103536 265900 103556
rect 265900 103536 265952 103556
rect 265952 103536 265954 103556
rect 265990 101496 266046 101552
rect 265898 100952 265954 101008
rect 265898 100136 265954 100192
rect 265990 96756 266046 96792
rect 265990 96736 265992 96756
rect 265992 96736 266044 96756
rect 266044 96736 266046 96756
rect 313278 389136 313334 389192
rect 306378 386416 306434 386472
rect 300858 384512 300914 384568
rect 269118 178744 269174 178800
rect 278778 177112 278834 177168
rect 278042 176160 278098 176216
rect 269946 175752 270002 175808
rect 267094 175344 267150 175400
rect 279330 173712 279386 173768
rect 280158 158480 280214 158536
rect 267186 123800 267242 123856
rect 281814 184184 281870 184240
rect 280434 169360 280490 169416
rect 280342 165416 280398 165472
rect 281814 173984 281870 174040
rect 282090 172352 282146 172408
rect 282274 170856 282330 170912
rect 281630 170040 281686 170096
rect 282826 168544 282882 168600
rect 281722 167728 281778 167784
rect 282458 167048 282514 167104
rect 282090 166232 282146 166288
rect 282090 164736 282146 164792
rect 282642 163920 282698 163976
rect 282826 163104 282882 163160
rect 282550 161608 282606 161664
rect 282366 160112 282422 160168
rect 282826 162424 282882 162480
rect 282826 160792 282882 160848
rect 282734 159296 282790 159352
rect 282274 157800 282330 157856
rect 282826 156984 282882 157040
rect 282826 155488 282882 155544
rect 281538 154672 281594 154728
rect 281906 153992 281962 154048
rect 281722 153176 281778 153232
rect 282182 152360 282238 152416
rect 282826 151716 282828 151736
rect 282828 151716 282880 151736
rect 282880 151716 282882 151736
rect 282826 151680 282882 151716
rect 281998 150864 282054 150920
rect 282826 150048 282882 150104
rect 282182 149368 282238 149424
rect 282090 148552 282146 148608
rect 281722 147056 281778 147112
rect 282826 146260 282882 146296
rect 282826 146240 282828 146260
rect 282828 146240 282880 146260
rect 282880 146240 282882 146260
rect 282734 145424 282790 145480
rect 282826 144744 282882 144800
rect 282826 143928 282882 143984
rect 282090 143112 282146 143168
rect 281906 133184 281962 133240
rect 281722 130092 281724 130112
rect 281724 130092 281776 130112
rect 281776 130092 281778 130112
rect 281722 130056 281778 130092
rect 281906 127744 281962 127800
rect 281998 123972 282000 123992
rect 282000 123972 282052 123992
rect 282052 123972 282054 123992
rect 281998 123936 282054 123972
rect 282274 142432 282330 142488
rect 282826 141616 282882 141672
rect 282734 140800 282790 140856
rect 282826 140120 282882 140176
rect 282826 139340 282828 139360
rect 282828 139340 282880 139360
rect 282880 139340 282882 139360
rect 282826 139304 282882 139340
rect 282734 138488 282790 138544
rect 282826 137808 282882 137864
rect 282826 136312 282882 136368
rect 282734 135496 282790 135552
rect 282826 134680 282882 134736
rect 282734 134000 282790 134056
rect 283010 147736 283066 147792
rect 282734 132368 282790 132424
rect 282826 131688 282882 131744
rect 282274 130872 282330 130928
rect 282826 128560 282882 128616
rect 282826 126248 282882 126304
rect 282826 125468 282828 125488
rect 282828 125468 282880 125488
rect 282880 125468 282882 125488
rect 282826 125432 282882 125468
rect 282734 124752 282790 124808
rect 282182 123120 282238 123176
rect 282090 122440 282146 122496
rect 282826 121624 282882 121680
rect 282826 120808 282882 120864
rect 282734 120128 282790 120184
rect 282826 119312 282882 119368
rect 281906 118532 281908 118552
rect 281908 118532 281960 118552
rect 281960 118532 281962 118552
rect 281906 118496 281962 118532
rect 282826 117816 282882 117872
rect 282826 117000 282882 117056
rect 282182 116320 282238 116376
rect 282090 115504 282146 115560
rect 281722 114688 281778 114744
rect 282274 114008 282330 114064
rect 282642 113192 282698 113248
rect 282090 112376 282146 112432
rect 282826 110880 282882 110936
rect 282826 109384 282882 109440
rect 282826 108568 282882 108624
rect 280250 107752 280306 107808
rect 282826 105440 282882 105496
rect 291290 177384 291346 177440
rect 281722 104760 281778 104816
rect 280250 103944 280306 104000
rect 280158 100816 280214 100872
rect 279422 97280 279478 97336
rect 279330 96600 279386 96656
rect 279330 95104 279386 95160
rect 281630 102448 281686 102504
rect 281538 100136 281594 100192
rect 280158 86808 280214 86864
rect 279514 3304 279570 3360
rect 298098 225528 298154 225584
rect 298190 196560 298246 196616
rect 304998 292576 305054 292632
rect 305274 179968 305330 180024
rect 288990 3440 289046 3496
rect 291382 3440 291438 3496
rect 293682 3440 293738 3496
rect 296074 3440 296130 3496
rect 298466 3848 298522 3904
rect 300766 3440 300822 3496
rect 303158 3576 303214 3632
rect 305550 3440 305606 3496
rect 310518 295296 310574 295352
rect 316038 366288 316094 366344
rect 307942 3848 307998 3904
rect 318798 360848 318854 360904
rect 322938 300056 322994 300112
rect 328458 335960 328514 336016
rect 327078 323584 327134 323640
rect 329838 177248 329894 177304
rect 332690 69536 332746 69592
rect 340878 283464 340934 283520
rect 343638 253136 343694 253192
rect 580170 378392 580226 378448
rect 580354 365064 580410 365120
rect 580262 351872 580318 351928
rect 579986 312024 580042 312080
rect 580354 325216 580410 325272
rect 582470 299512 582526 299568
rect 580354 298696 580410 298752
rect 580262 272176 580318 272232
rect 579802 258848 579858 258904
rect 580262 255856 580318 255912
rect 580170 245520 580226 245576
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580354 246336 580410 246392
rect 580538 232328 580594 232384
rect 580446 205672 580502 205728
rect 580262 139304 580318 139360
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 582562 219000 582618 219056
rect 582470 72936 582526 72992
rect 582378 19760 582434 19816
rect 582746 235184 582802 235240
rect 582654 112784 582710 112840
rect 582838 179152 582894 179208
rect 582746 86128 582802 86184
rect 582562 6568 582618 6624
<< metal3 >>
rect 111006 702476 111012 702540
rect 111076 702538 111082 702540
rect 348785 702538 348851 702541
rect 111076 702536 348851 702538
rect 111076 702480 348790 702536
rect 348846 702480 348851 702536
rect 111076 702478 348851 702480
rect 111076 702476 111082 702478
rect 348785 702475 348851 702478
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 57830 586332 57836 586396
rect 57900 586394 57906 586396
rect 83181 586394 83247 586397
rect 57900 586392 83247 586394
rect 57900 586336 83186 586392
rect 83242 586336 83247 586392
rect 57900 586334 83247 586336
rect 57900 586332 57906 586334
rect 83181 586331 83247 586334
rect 74625 584354 74691 584357
rect 64830 584352 74691 584354
rect 64830 584296 74630 584352
rect 74686 584296 74691 584352
rect 64830 584294 74691 584296
rect 55857 584082 55923 584085
rect 56501 584082 56567 584085
rect 64830 584082 64890 584294
rect 74625 584291 74691 584294
rect 55857 584080 64890 584082
rect 55857 584024 55862 584080
rect 55918 584024 56506 584080
rect 56562 584024 64890 584080
rect 55857 584022 64890 584024
rect 91001 584082 91067 584085
rect 115974 584082 115980 584084
rect 91001 584080 115980 584082
rect 91001 584024 91006 584080
rect 91062 584024 115980 584080
rect 91001 584022 115980 584024
rect 55857 584019 55923 584022
rect 56501 584019 56567 584022
rect 91001 584019 91067 584022
rect 115974 584020 115980 584022
rect 116044 584020 116050 584084
rect 53833 583946 53899 583949
rect 55029 583946 55095 583949
rect 71773 583946 71839 583949
rect 53833 583944 71839 583946
rect 53833 583888 53838 583944
rect 53894 583888 55034 583944
rect 55090 583888 71778 583944
rect 71834 583888 71839 583944
rect 53833 583886 71839 583888
rect 53833 583883 53899 583886
rect 55029 583883 55095 583886
rect 71773 583883 71839 583886
rect 84377 583946 84443 583949
rect 107101 583946 107167 583949
rect 84377 583944 107167 583946
rect 84377 583888 84382 583944
rect 84438 583888 107106 583944
rect 107162 583888 107167 583944
rect 84377 583886 107167 583888
rect 84377 583883 84443 583886
rect 107101 583883 107167 583886
rect 48037 583810 48103 583813
rect 84469 583810 84535 583813
rect 48037 583808 84535 583810
rect 48037 583752 48042 583808
rect 48098 583752 84474 583808
rect 84530 583752 84535 583808
rect 48037 583750 84535 583752
rect 48037 583747 48103 583750
rect 84469 583747 84535 583750
rect 97901 583810 97967 583813
rect 106733 583810 106799 583813
rect 97901 583808 106799 583810
rect 97901 583752 97906 583808
rect 97962 583752 106738 583808
rect 106794 583752 106799 583808
rect 97901 583750 106799 583752
rect 97901 583747 97967 583750
rect 106733 583747 106799 583750
rect 92841 582450 92907 582453
rect 109125 582450 109191 582453
rect 92841 582448 109191 582450
rect 92841 582392 92846 582448
rect 92902 582392 109130 582448
rect 109186 582392 109191 582448
rect 92841 582390 109191 582392
rect 92841 582387 92907 582390
rect 109125 582387 109191 582390
rect 102593 581770 102659 581773
rect 114502 581770 114508 581772
rect 102593 581768 114508 581770
rect 102593 581712 102598 581768
rect 102654 581712 114508 581768
rect 102593 581710 114508 581712
rect 102593 581707 102659 581710
rect 114502 581708 114508 581710
rect 114572 581708 114578 581772
rect 67633 581362 67699 581365
rect 70166 581362 70226 581468
rect 67633 581360 70226 581362
rect 67633 581304 67638 581360
rect 67694 581304 70226 581360
rect 67633 581302 70226 581304
rect 67633 581299 67699 581302
rect 108941 580818 109007 580821
rect 105892 580816 109007 580818
rect 67909 580682 67975 580685
rect 68553 580682 68619 580685
rect 70166 580682 70226 580788
rect 105892 580760 108946 580816
rect 109002 580760 109007 580816
rect 105892 580758 109007 580760
rect 108941 580755 109007 580758
rect 67909 580680 70226 580682
rect 67909 580624 67914 580680
rect 67970 580624 68558 580680
rect 68614 580624 70226 580680
rect 67909 580622 70226 580624
rect 67909 580619 67975 580622
rect 68553 580619 68619 580622
rect 108849 580138 108915 580141
rect 105892 580136 108915 580138
rect -960 580002 480 580092
rect 105892 580080 108854 580136
rect 108910 580080 108915 580136
rect 105892 580078 108915 580080
rect 108849 580075 108915 580078
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 108849 579458 108915 579461
rect 105892 579456 108915 579458
rect 67357 579186 67423 579189
rect 70166 579186 70226 579428
rect 105892 579400 108854 579456
rect 108910 579400 108915 579456
rect 105892 579398 108915 579400
rect 108849 579395 108915 579398
rect 67357 579184 70226 579186
rect 67357 579128 67362 579184
rect 67418 579128 70226 579184
rect 67357 579126 70226 579128
rect 67357 579123 67423 579126
rect 107101 578914 107167 578917
rect 118734 578914 118740 578916
rect 107101 578912 118740 578914
rect 107101 578856 107106 578912
rect 107162 578856 118740 578912
rect 107101 578854 118740 578856
rect 107101 578851 107167 578854
rect 118734 578852 118740 578854
rect 118804 578852 118810 578916
rect 108941 578778 109007 578781
rect 105892 578776 109007 578778
rect 67633 578506 67699 578509
rect 70166 578506 70226 578748
rect 105892 578720 108946 578776
rect 109002 578720 109007 578776
rect 105892 578718 109007 578720
rect 108941 578715 109007 578718
rect 67633 578504 70226 578506
rect 67633 578448 67638 578504
rect 67694 578448 70226 578504
rect 67633 578446 70226 578448
rect 67633 578443 67699 578446
rect 111701 578236 111767 578237
rect 111701 578232 111748 578236
rect 111812 578234 111818 578236
rect 111701 578176 111706 578232
rect 111701 578172 111748 578176
rect 111812 578174 111858 578234
rect 111812 578172 111818 578174
rect 111701 578171 111767 578172
rect 106457 578098 106523 578101
rect 105892 578096 106523 578098
rect 67633 577826 67699 577829
rect 70166 577826 70226 578068
rect 105892 578040 106462 578096
rect 106518 578040 106523 578096
rect 105892 578038 106523 578040
rect 106457 578035 106523 578038
rect 67633 577824 70226 577826
rect 67633 577768 67638 577824
rect 67694 577768 70226 577824
rect 67633 577766 70226 577768
rect 67633 577763 67699 577766
rect 579797 577690 579863 577693
rect 583520 577690 584960 577780
rect 579797 577688 584960 577690
rect 579797 577632 579802 577688
rect 579858 577632 584960 577688
rect 579797 577630 584960 577632
rect 579797 577627 579863 577630
rect 108205 577554 108271 577557
rect 105892 577552 108271 577554
rect 105892 577496 108210 577552
rect 108266 577496 108271 577552
rect 583520 577540 584960 577630
rect 105892 577494 108271 577496
rect 108205 577491 108271 577494
rect 66110 577084 66116 577148
rect 66180 577146 66186 577148
rect 70166 577146 70226 577388
rect 66180 577086 70226 577146
rect 66180 577084 66186 577086
rect 108849 576738 108915 576741
rect 105892 576736 108915 576738
rect 68829 576466 68895 576469
rect 70166 576466 70226 576708
rect 105892 576680 108854 576736
rect 108910 576680 108915 576736
rect 105892 576678 108915 576680
rect 108849 576675 108915 576678
rect 68829 576464 70226 576466
rect 68829 576408 68834 576464
rect 68890 576408 70226 576464
rect 68829 576406 70226 576408
rect 68829 576403 68895 576406
rect 108941 576058 109007 576061
rect 105892 576056 109007 576058
rect 67633 575786 67699 575789
rect 70166 575786 70226 576028
rect 105892 576000 108946 576056
rect 109002 576000 109007 576056
rect 105892 575998 109007 576000
rect 108941 575995 109007 575998
rect 67633 575784 70226 575786
rect 67633 575728 67638 575784
rect 67694 575728 70226 575784
rect 67633 575726 70226 575728
rect 67633 575723 67699 575726
rect 67725 575106 67791 575109
rect 70166 575106 70226 575348
rect 67725 575104 70226 575106
rect 67725 575048 67730 575104
rect 67786 575048 70226 575104
rect 67725 575046 70226 575048
rect 67725 575043 67791 575046
rect 106365 574698 106431 574701
rect 105892 574696 106431 574698
rect 67633 574426 67699 574429
rect 70166 574426 70226 574668
rect 105892 574640 106370 574696
rect 106426 574640 106431 574696
rect 105892 574638 106431 574640
rect 106365 574635 106431 574638
rect 67633 574424 70226 574426
rect 67633 574368 67638 574424
rect 67694 574368 70226 574424
rect 67633 574366 70226 574368
rect 67633 574363 67699 574366
rect 108941 574018 109007 574021
rect 105892 574016 109007 574018
rect 67725 573474 67791 573477
rect 70166 573474 70226 573988
rect 105892 573960 108946 574016
rect 109002 573960 109007 574016
rect 105892 573958 109007 573960
rect 108941 573955 109007 573958
rect 67725 573472 70226 573474
rect 67725 573416 67730 573472
rect 67786 573416 70226 573472
rect 67725 573414 70226 573416
rect 67725 573411 67791 573414
rect 107653 573338 107719 573341
rect 107837 573338 107903 573341
rect 105892 573336 107903 573338
rect 105892 573280 107658 573336
rect 107714 573280 107842 573336
rect 107898 573280 107903 573336
rect 105892 573278 107903 573280
rect 107653 573275 107719 573278
rect 107837 573275 107903 573278
rect 67633 572794 67699 572797
rect 69982 572794 70226 572828
rect 108941 572794 109007 572797
rect 67633 572792 70226 572794
rect 67633 572736 67638 572792
rect 67694 572768 70226 572792
rect 67694 572736 70042 572768
rect 70166 572764 70226 572768
rect 105892 572792 109007 572794
rect 67633 572734 70042 572736
rect 105892 572736 108946 572792
rect 109002 572736 109007 572792
rect 105892 572734 109007 572736
rect 67633 572731 67699 572734
rect 108941 572731 109007 572734
rect 108941 571978 109007 571981
rect 105892 571976 109007 571978
rect 66662 571780 66668 571844
rect 66732 571842 66738 571844
rect 68645 571842 68711 571845
rect 70166 571842 70226 571948
rect 105892 571920 108946 571976
rect 109002 571920 109007 571976
rect 105892 571918 109007 571920
rect 108941 571915 109007 571918
rect 66732 571840 70226 571842
rect 66732 571784 68650 571840
rect 68706 571784 70226 571840
rect 66732 571782 70226 571784
rect 66732 571780 66738 571782
rect 68645 571779 68711 571782
rect 68277 571706 68343 571709
rect 68461 571706 68527 571709
rect 68277 571704 70410 571706
rect 68277 571648 68282 571704
rect 68338 571648 68466 571704
rect 68522 571648 70410 571704
rect 68277 571646 70410 571648
rect 68277 571643 68343 571646
rect 68461 571643 68527 571646
rect 70350 571404 70410 571646
rect 107929 571434 107995 571437
rect 105892 571432 107995 571434
rect 105892 571376 107934 571432
rect 107990 571376 107995 571432
rect 105892 571374 107995 571376
rect 107929 571371 107995 571374
rect 108849 570618 108915 570621
rect 105892 570616 108915 570618
rect 68870 570284 68876 570348
rect 68940 570346 68946 570348
rect 70166 570346 70226 570588
rect 105892 570560 108854 570616
rect 108910 570560 108915 570616
rect 105892 570558 108915 570560
rect 108849 570555 108915 570558
rect 68940 570286 70226 570346
rect 68940 570284 68946 570286
rect 67633 570074 67699 570077
rect 108941 570074 109007 570077
rect 67633 570072 70042 570074
rect 67633 570016 67638 570072
rect 67694 570016 70042 570072
rect 67633 570014 70042 570016
rect 105892 570072 109007 570074
rect 105892 570016 108946 570072
rect 109002 570016 109007 570072
rect 105892 570014 109007 570016
rect 67633 570011 67699 570014
rect 69982 569802 70042 570014
rect 108941 570011 109007 570014
rect 70166 569802 70226 569908
rect 69982 569742 70226 569802
rect 108941 569258 109007 569261
rect 105892 569256 109007 569258
rect 67633 568986 67699 568989
rect 70166 568986 70226 569228
rect 105892 569200 108946 569256
rect 109002 569200 109007 569256
rect 105892 569198 109007 569200
rect 108941 569195 109007 569198
rect 67633 568984 70226 568986
rect 67633 568928 67638 568984
rect 67694 568928 70226 568984
rect 67633 568926 70226 568928
rect 67633 568923 67699 568926
rect 67173 568714 67239 568717
rect 67173 568712 70042 568714
rect 67173 568656 67178 568712
rect 67234 568680 70042 568712
rect 70166 568680 70226 568684
rect 67234 568656 70226 568680
rect 67173 568654 70226 568656
rect 67173 568651 67239 568654
rect 69982 568620 70226 568654
rect 108941 567898 109007 567901
rect 105892 567896 109007 567898
rect 67541 567626 67607 567629
rect 70166 567626 70226 567868
rect 105892 567840 108946 567896
rect 109002 567840 109007 567896
rect 105892 567838 109007 567840
rect 108941 567835 109007 567838
rect 67541 567624 70226 567626
rect 67541 567568 67546 567624
rect 67602 567568 70226 567624
rect 67541 567566 70226 567568
rect 67541 567563 67607 567566
rect 67633 567218 67699 567221
rect 108941 567218 109007 567221
rect 67633 567216 70042 567218
rect 67633 567160 67638 567216
rect 67694 567210 70042 567216
rect 105892 567216 109007 567218
rect 67694 567160 70226 567210
rect 67633 567158 70226 567160
rect 105892 567160 108946 567216
rect 109002 567160 109007 567216
rect 105892 567158 109007 567160
rect 67633 567155 67699 567158
rect 69982 567150 70226 567158
rect 108941 567155 109007 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 108849 566538 108915 566541
rect 105892 566536 108915 566538
rect 105892 566480 108854 566536
rect 108910 566480 108915 566536
rect 105892 566478 108915 566480
rect 108849 566475 108915 566478
rect 64638 565796 64644 565860
rect 64708 565858 64714 565860
rect 108941 565858 109007 565861
rect 64708 565798 70042 565858
rect 105892 565856 109007 565858
rect 64708 565796 64714 565798
rect 69982 565722 70042 565798
rect 70166 565722 70226 565828
rect 105892 565800 108946 565856
rect 109002 565800 109007 565856
rect 105892 565798 109007 565800
rect 108941 565795 109007 565798
rect 69982 565662 70226 565722
rect 108941 565178 109007 565181
rect 105892 565176 109007 565178
rect 67633 564906 67699 564909
rect 70166 564906 70226 565148
rect 105892 565120 108946 565176
rect 109002 565120 109007 565176
rect 105892 565118 109007 565120
rect 108941 565115 109007 565118
rect 67633 564904 70226 564906
rect 67633 564848 67638 564904
rect 67694 564848 70226 564904
rect 67633 564846 70226 564848
rect 67633 564843 67699 564846
rect 67725 564498 67791 564501
rect 106406 564498 106412 564500
rect 67725 564496 70042 564498
rect 67725 564440 67730 564496
rect 67786 564440 70042 564496
rect 67725 564438 70042 564440
rect 67725 564435 67791 564438
rect 69982 564362 70042 564438
rect 70166 564362 70226 564468
rect 105892 564438 106412 564498
rect 106406 564436 106412 564438
rect 106476 564436 106482 564500
rect 69982 564302 70226 564362
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 67725 564226 67791 564229
rect 67725 564224 70410 564226
rect 67725 564168 67730 564224
rect 67786 564168 70410 564224
rect 583520 564212 584960 564302
rect 67725 564166 70410 564168
rect 67725 564163 67791 564166
rect 70350 563924 70410 564166
rect 108941 563818 109007 563821
rect 105892 563816 109007 563818
rect 105892 563760 108946 563816
rect 109002 563760 109007 563816
rect 105892 563758 109007 563760
rect 108941 563755 109007 563758
rect 67633 563682 67699 563685
rect 67633 563680 70410 563682
rect 67633 563624 67638 563680
rect 67694 563624 70410 563680
rect 67633 563622 70410 563624
rect 67633 563619 67699 563622
rect 70350 563244 70410 563622
rect 107745 563138 107811 563141
rect 105892 563136 107811 563138
rect 105892 563080 107750 563136
rect 107806 563080 107811 563136
rect 105892 563078 107811 563080
rect 107745 563075 107811 563078
rect 67633 563002 67699 563005
rect 67633 563000 70226 563002
rect 67633 562944 67638 563000
rect 67694 562944 70226 563000
rect 67633 562942 70226 562944
rect 67633 562939 67699 562942
rect 70166 562564 70226 562942
rect 64830 562126 70410 562186
rect 61878 561852 61884 561916
rect 61948 561914 61954 561916
rect 64830 561914 64890 562126
rect 61948 561854 64890 561914
rect 70350 561884 70410 562126
rect 105494 561916 105554 562428
rect 61948 561852 61954 561854
rect 105486 561852 105492 561916
rect 105556 561852 105562 561916
rect 108941 561098 109007 561101
rect 105892 561096 109007 561098
rect 70166 560826 70226 561068
rect 105892 561040 108946 561096
rect 109002 561040 109007 561096
rect 105892 561038 109007 561040
rect 108941 561035 109007 561038
rect 64830 560766 70226 560826
rect 60590 560492 60596 560556
rect 60660 560554 60666 560556
rect 64830 560554 64890 560766
rect 60660 560494 64890 560554
rect 60660 560492 60666 560494
rect 67633 560418 67699 560421
rect 106273 560418 106339 560421
rect 107653 560418 107719 560421
rect 67633 560416 70042 560418
rect 67633 560360 67638 560416
rect 67694 560360 70042 560416
rect 105892 560416 107719 560418
rect 67633 560358 70042 560360
rect 67633 560355 67699 560358
rect 69982 560282 70042 560358
rect 70166 560282 70226 560388
rect 105892 560360 106278 560416
rect 106334 560360 107658 560416
rect 107714 560360 107719 560416
rect 105892 560358 107719 560360
rect 106273 560355 106339 560358
rect 107653 560355 107719 560358
rect 69982 560222 70226 560282
rect 108849 559738 108915 559741
rect 105892 559736 108915 559738
rect 105892 559680 108854 559736
rect 108910 559680 108915 559736
rect 105892 559678 108915 559680
rect 108849 559675 108915 559678
rect 67633 559466 67699 559469
rect 67633 559464 70410 559466
rect 67633 559408 67638 559464
rect 67694 559408 70410 559464
rect 67633 559406 70410 559408
rect 67633 559403 67699 559406
rect 70350 559164 70410 559406
rect 108941 559058 109007 559061
rect 105892 559056 109007 559058
rect 105892 559000 108946 559056
rect 109002 559000 109007 559056
rect 105892 558998 109007 559000
rect 108941 558995 109007 558998
rect 68369 558922 68435 558925
rect 69105 558922 69171 558925
rect 68369 558920 70226 558922
rect 68369 558864 68374 558920
rect 68430 558864 69110 558920
rect 69166 558864 70226 558920
rect 68369 558862 70226 558864
rect 68369 558859 68435 558862
rect 69105 558859 69171 558862
rect 70166 558484 70226 558862
rect 108573 558378 108639 558381
rect 105892 558376 108639 558378
rect 105892 558320 108578 558376
rect 108634 558320 108639 558376
rect 105892 558318 108639 558320
rect 108573 558315 108639 558318
rect 107694 557698 107700 557700
rect 67633 557562 67699 557565
rect 70166 557562 70226 557668
rect 105892 557638 107700 557698
rect 107694 557636 107700 557638
rect 107764 557636 107770 557700
rect 67633 557560 70226 557562
rect 67633 557504 67638 557560
rect 67694 557504 70226 557560
rect 67633 557502 70226 557504
rect 67633 557499 67699 557502
rect 108941 557018 109007 557021
rect 105892 557016 109007 557018
rect 67725 556746 67791 556749
rect 70166 556746 70226 556988
rect 105892 556960 108946 557016
rect 109002 556960 109007 557016
rect 105892 556958 109007 556960
rect 108941 556955 109007 556958
rect 67725 556744 70226 556746
rect 67725 556688 67730 556744
rect 67786 556688 70226 556744
rect 67725 556686 70226 556688
rect 67725 556683 67791 556686
rect 107653 556338 107719 556341
rect 105892 556336 107719 556338
rect 67633 556202 67699 556205
rect 70166 556202 70226 556308
rect 105892 556280 107658 556336
rect 107714 556280 107719 556336
rect 105892 556278 107719 556280
rect 107653 556275 107719 556278
rect 67633 556200 70226 556202
rect 67633 556144 67638 556200
rect 67694 556144 70226 556200
rect 67633 556142 70226 556144
rect 67633 556139 67699 556142
rect 109217 555794 109283 555797
rect 105892 555792 109283 555794
rect 105892 555736 109222 555792
rect 109278 555736 109283 555792
rect 105892 555734 109283 555736
rect 109217 555731 109283 555734
rect 67633 555386 67699 555389
rect 70166 555386 70226 555628
rect 67633 555384 70226 555386
rect 67633 555328 67638 555384
rect 67694 555328 70226 555384
rect 67633 555326 70226 555328
rect 67633 555323 67699 555326
rect 67725 554842 67791 554845
rect 70166 554842 70226 554948
rect 67725 554840 70226 554842
rect 67725 554784 67730 554840
rect 67786 554784 70226 554840
rect 67725 554782 70226 554784
rect 67725 554779 67791 554782
rect 108941 554298 109007 554301
rect 105892 554296 109007 554298
rect 69105 554026 69171 554029
rect 70166 554026 70226 554268
rect 105892 554240 108946 554296
rect 109002 554240 109007 554296
rect 105892 554238 109007 554240
rect 108941 554235 109007 554238
rect 69105 554024 70226 554026
rect -960 553890 480 553980
rect 69105 553968 69110 554024
rect 69166 553968 70226 554024
rect 69105 553966 70226 553968
rect 69105 553963 69171 553966
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 108941 553618 109007 553621
rect 105892 553616 109007 553618
rect 67633 553482 67699 553485
rect 70166 553482 70226 553588
rect 105892 553560 108946 553616
rect 109002 553560 109007 553616
rect 105892 553558 109007 553560
rect 108941 553555 109007 553558
rect 67633 553480 70226 553482
rect 67633 553424 67638 553480
rect 67694 553424 70226 553480
rect 67633 553422 70226 553424
rect 67633 553419 67699 553422
rect 108941 552938 109007 552941
rect 105892 552936 109007 552938
rect 105892 552880 108946 552936
rect 109002 552880 109007 552936
rect 105892 552878 109007 552880
rect 108941 552875 109007 552878
rect 67633 552122 67699 552125
rect 70166 552122 70226 552228
rect 67633 552120 70226 552122
rect 67633 552064 67638 552120
rect 67694 552064 70226 552120
rect 67633 552062 70226 552064
rect 105862 552122 105922 552228
rect 106181 552122 106247 552125
rect 105862 552120 106247 552122
rect 105862 552064 106186 552120
rect 106242 552064 106247 552120
rect 105862 552062 106247 552064
rect 67633 552059 67699 552062
rect 106181 552059 106247 552062
rect 106917 551578 106983 551581
rect 105892 551576 106983 551578
rect 67633 551306 67699 551309
rect 70166 551306 70226 551548
rect 105892 551520 106922 551576
rect 106978 551520 106983 551576
rect 105892 551518 106983 551520
rect 106917 551515 106983 551518
rect 67633 551304 70226 551306
rect 67633 551248 67638 551304
rect 67694 551248 70226 551304
rect 67633 551246 70226 551248
rect 67633 551243 67699 551246
rect 583520 551020 584960 551260
rect 108941 550898 109007 550901
rect 105892 550896 109007 550898
rect 68277 550762 68343 550765
rect 70166 550762 70226 550868
rect 105892 550840 108946 550896
rect 109002 550840 109007 550896
rect 105892 550838 109007 550840
rect 108941 550835 109007 550838
rect 68277 550760 70226 550762
rect 68277 550704 68282 550760
rect 68338 550704 70226 550760
rect 68277 550702 70226 550704
rect 68277 550699 68343 550702
rect 108849 550218 108915 550221
rect 105892 550216 108915 550218
rect 67725 549946 67791 549949
rect 70166 549946 70226 550188
rect 105892 550160 108854 550216
rect 108910 550160 108915 550216
rect 105892 550158 108915 550160
rect 108849 550155 108915 550158
rect 67725 549944 70226 549946
rect 67725 549888 67730 549944
rect 67786 549888 70226 549944
rect 67725 549886 70226 549888
rect 67725 549883 67791 549886
rect 108941 549538 109007 549541
rect 105892 549536 109007 549538
rect 67633 549402 67699 549405
rect 70166 549402 70226 549508
rect 105892 549480 108946 549536
rect 109002 549480 109007 549536
rect 105892 549478 109007 549480
rect 108941 549475 109007 549478
rect 67633 549400 70226 549402
rect 67633 549344 67638 549400
rect 67694 549344 70226 549400
rect 67633 549342 70226 549344
rect 67633 549339 67699 549342
rect 107837 548858 107903 548861
rect 105892 548856 107903 548858
rect 67633 548586 67699 548589
rect 70166 548586 70226 548828
rect 105892 548800 107842 548856
rect 107898 548800 107903 548856
rect 105892 548798 107903 548800
rect 107837 548795 107903 548798
rect 67633 548584 70226 548586
rect 67633 548528 67638 548584
rect 67694 548528 70226 548584
rect 67633 548526 70226 548528
rect 67633 548523 67699 548526
rect 62982 547980 62988 548044
rect 63052 548042 63058 548044
rect 70166 548042 70226 548148
rect 63052 547982 70226 548042
rect 63052 547980 63058 547982
rect 108941 547498 109007 547501
rect 105892 547496 109007 547498
rect 67725 547226 67791 547229
rect 70166 547226 70226 547468
rect 105892 547440 108946 547496
rect 109002 547440 109007 547496
rect 105892 547438 109007 547440
rect 108941 547435 109007 547438
rect 67725 547224 70226 547226
rect 67725 547168 67730 547224
rect 67786 547168 70226 547224
rect 67725 547166 70226 547168
rect 67725 547163 67791 547166
rect 107878 546818 107884 546820
rect 67633 546546 67699 546549
rect 70166 546546 70226 546788
rect 105892 546758 107884 546818
rect 107878 546756 107884 546758
rect 107948 546756 107954 546820
rect 67633 546544 70226 546546
rect 67633 546488 67638 546544
rect 67694 546488 70226 546544
rect 67633 546486 70226 546488
rect 67633 546483 67699 546486
rect 108941 546138 109007 546141
rect 105892 546136 109007 546138
rect 105892 546080 108946 546136
rect 109002 546080 109007 546136
rect 105892 546078 109007 546080
rect 108941 546075 109007 546078
rect 68737 545866 68803 545869
rect 68737 545864 70410 545866
rect 68737 545808 68742 545864
rect 68798 545808 70410 545864
rect 68737 545806 70410 545808
rect 68737 545803 68803 545806
rect 70350 545564 70410 545806
rect 108941 545458 109007 545461
rect 105892 545456 109007 545458
rect 105892 545400 108946 545456
rect 109002 545400 109007 545456
rect 105892 545398 109007 545400
rect 108941 545395 109007 545398
rect 108941 544778 109007 544781
rect 105892 544776 109007 544778
rect 67725 544506 67791 544509
rect 70166 544506 70226 544748
rect 105892 544720 108946 544776
rect 109002 544720 109007 544776
rect 105892 544718 109007 544720
rect 108941 544715 109007 544718
rect 67725 544504 70226 544506
rect 67725 544448 67730 544504
rect 67786 544448 70226 544504
rect 67725 544446 70226 544448
rect 67725 544443 67791 544446
rect 67633 543826 67699 543829
rect 70166 543826 70226 544068
rect 105862 543829 105922 544068
rect 67633 543824 70226 543826
rect 67633 543768 67638 543824
rect 67694 543768 70226 543824
rect 67633 543766 70226 543768
rect 105813 543824 105922 543829
rect 105813 543768 105818 543824
rect 105874 543768 105922 543824
rect 105813 543766 105922 543768
rect 67633 543763 67699 543766
rect 105813 543763 105879 543766
rect 108941 543418 109007 543421
rect 105892 543416 109007 543418
rect 68921 543282 68987 543285
rect 70166 543282 70226 543388
rect 105892 543360 108946 543416
rect 109002 543360 109007 543416
rect 105892 543358 109007 543360
rect 108941 543355 109007 543358
rect 68921 543280 70226 543282
rect 68921 543224 68926 543280
rect 68982 543224 70226 543280
rect 68921 543222 70226 543224
rect 68921 543219 68987 543222
rect 107653 542738 107719 542741
rect 105892 542736 107719 542738
rect 67633 542602 67699 542605
rect 70166 542602 70226 542708
rect 105892 542680 107658 542736
rect 107714 542680 107719 542736
rect 105892 542678 107719 542680
rect 107653 542675 107719 542678
rect 67633 542600 70226 542602
rect 67633 542544 67638 542600
rect 67694 542544 70226 542600
rect 67633 542542 70226 542544
rect 67633 542539 67699 542542
rect 108941 542058 109007 542061
rect 105892 542056 109007 542058
rect 68921 541786 68987 541789
rect 70166 541786 70226 542028
rect 105892 542000 108946 542056
rect 109002 542000 109007 542056
rect 105892 541998 109007 542000
rect 108941 541995 109007 541998
rect 68921 541784 70226 541786
rect 68921 541728 68926 541784
rect 68982 541728 70226 541784
rect 68921 541726 70226 541728
rect 68921 541723 68987 541726
rect 67633 541242 67699 541245
rect 70166 541242 70226 541348
rect 67633 541240 70226 541242
rect 67633 541184 67638 541240
rect 67694 541184 70226 541240
rect 67633 541182 70226 541184
rect 67633 541179 67699 541182
rect -960 540684 480 540924
rect 67633 540154 67699 540157
rect 70166 540154 70226 540668
rect 105862 540426 105922 540668
rect 106089 540426 106155 540429
rect 105862 540424 106155 540426
rect 105862 540368 106094 540424
rect 106150 540368 106155 540424
rect 105862 540366 106155 540368
rect 106089 540363 106155 540366
rect 107561 540154 107627 540157
rect 111006 540154 111012 540156
rect 67633 540152 70226 540154
rect 67633 540096 67638 540152
rect 67694 540096 70226 540152
rect 67633 540094 70226 540096
rect 105892 540152 111012 540154
rect 105892 540096 107566 540152
rect 107622 540096 111012 540152
rect 105892 540094 111012 540096
rect 67633 540091 67699 540094
rect 107561 540091 107627 540094
rect 111006 540092 111012 540094
rect 111076 540092 111082 540156
rect 59077 538794 59143 538797
rect 70342 538794 70348 538796
rect 59077 538792 70348 538794
rect 59077 538736 59082 538792
rect 59138 538736 70348 538792
rect 59077 538734 70348 538736
rect 59077 538731 59143 538734
rect 70342 538732 70348 538734
rect 70412 538732 70418 538796
rect 103646 538052 103652 538116
rect 103716 538114 103722 538116
rect 104801 538114 104867 538117
rect 103716 538112 104867 538114
rect 103716 538056 104806 538112
rect 104862 538056 104867 538112
rect 103716 538054 104867 538056
rect 103716 538052 103722 538054
rect 104801 538051 104867 538054
rect 102041 537978 102107 537981
rect 109769 537978 109835 537981
rect 102041 537976 109835 537978
rect 102041 537920 102046 537976
rect 102102 537920 109774 537976
rect 109830 537920 109835 537976
rect 102041 537918 109835 537920
rect 102041 537915 102107 537918
rect 109769 537915 109835 537918
rect 104709 537842 104775 537845
rect 111793 537842 111859 537845
rect 104709 537840 111859 537842
rect 104709 537784 104714 537840
rect 104770 537784 111798 537840
rect 111854 537784 111859 537840
rect 104709 537782 111859 537784
rect 104709 537779 104775 537782
rect 111793 537779 111859 537782
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect 57830 537508 57836 537572
rect 57900 537570 57906 537572
rect 76557 537570 76623 537573
rect 57900 537568 76623 537570
rect 57900 537512 76562 537568
rect 76618 537512 76623 537568
rect 57900 537510 76623 537512
rect 57900 537508 57906 537510
rect 76557 537507 76623 537510
rect 57830 537372 57836 537436
rect 57900 537434 57906 537436
rect 81617 537434 81683 537437
rect 57900 537432 81683 537434
rect 57900 537376 81622 537432
rect 81678 537376 81683 537432
rect 57900 537374 81683 537376
rect 57900 537372 57906 537374
rect 81617 537371 81683 537374
rect 89345 537434 89411 537437
rect 98494 537434 98500 537436
rect 89345 537432 98500 537434
rect 89345 537376 89350 537432
rect 89406 537376 98500 537432
rect 89345 537374 98500 537376
rect 89345 537371 89411 537374
rect 98494 537372 98500 537374
rect 98564 537372 98570 537436
rect 100937 537026 101003 537029
rect 102041 537026 102107 537029
rect 100937 537024 102107 537026
rect 100937 536968 100942 537024
rect 100998 536968 102046 537024
rect 102102 536968 102107 537024
rect 100937 536966 102107 536968
rect 100937 536963 101003 536966
rect 102041 536963 102107 536966
rect 99373 536890 99439 536893
rect 105537 536890 105603 536893
rect 99373 536888 105603 536890
rect 99373 536832 99378 536888
rect 99434 536832 105542 536888
rect 105598 536832 105603 536888
rect 99373 536830 105603 536832
rect 99373 536827 99439 536830
rect 105537 536827 105603 536830
rect 97901 536074 97967 536077
rect 114502 536074 114508 536076
rect 97901 536072 114508 536074
rect 97901 536016 97906 536072
rect 97962 536016 114508 536072
rect 97901 536014 114508 536016
rect 97901 536011 97967 536014
rect 114502 536012 114508 536014
rect 114572 536012 114578 536076
rect 53598 532204 53604 532268
rect 53668 532266 53674 532268
rect 70393 532266 70459 532269
rect 53668 532264 70459 532266
rect 53668 532208 70398 532264
rect 70454 532208 70459 532264
rect 53668 532206 70459 532208
rect 53668 532204 53674 532206
rect 70393 532203 70459 532206
rect 48078 532068 48084 532132
rect 48148 532130 48154 532132
rect 76465 532130 76531 532133
rect 48148 532128 76531 532130
rect 48148 532072 76470 532128
rect 76526 532072 76531 532128
rect 48148 532070 76531 532072
rect 48148 532068 48154 532070
rect 76465 532067 76531 532070
rect 44030 531932 44036 531996
rect 44100 531994 44106 531996
rect 74533 531994 74599 531997
rect 44100 531992 74599 531994
rect 44100 531936 74538 531992
rect 74594 531936 74599 531992
rect 44100 531934 74599 531936
rect 44100 531932 44106 531934
rect 74533 531931 74599 531934
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 583520 497844 584960 498084
rect 77753 495546 77819 495549
rect 118734 495546 118740 495548
rect 77753 495544 118740 495546
rect 77753 495488 77758 495544
rect 77814 495488 118740 495544
rect 77753 495486 118740 495488
rect 77753 495483 77819 495486
rect 118734 495484 118740 495486
rect 118804 495484 118810 495548
rect 118734 494940 118740 495004
rect 118804 495002 118810 495004
rect 119981 495002 120047 495005
rect 118804 495000 120047 495002
rect 118804 494944 119986 495000
rect 120042 494944 120047 495000
rect 118804 494942 120047 494944
rect 118804 494940 118810 494942
rect 119981 494939 120047 494942
rect 50838 494804 50844 494868
rect 50908 494866 50914 494868
rect 52085 494866 52151 494869
rect 50908 494864 52151 494866
rect 50908 494808 52090 494864
rect 52146 494808 52151 494864
rect 50908 494806 52151 494808
rect 50908 494804 50914 494806
rect 52085 494803 52151 494806
rect 90633 494730 90699 494733
rect 124438 494730 124444 494732
rect 90633 494728 124444 494730
rect 90633 494672 90638 494728
rect 90694 494672 124444 494728
rect 90633 494670 124444 494672
rect 90633 494667 90699 494670
rect 124438 494668 124444 494670
rect 124508 494668 124514 494732
rect 52085 492690 52151 492693
rect 52310 492690 52316 492692
rect 52085 492688 52316 492690
rect 52085 492632 52090 492688
rect 52146 492632 52316 492688
rect 52085 492630 52316 492632
rect 52085 492627 52151 492630
rect 52310 492628 52316 492630
rect 52380 492628 52386 492692
rect 53046 491948 53052 492012
rect 53116 492010 53122 492012
rect 53281 492010 53347 492013
rect 53116 492008 53347 492010
rect 53116 491952 53286 492008
rect 53342 491952 53347 492008
rect 53116 491950 53347 491952
rect 53116 491948 53122 491950
rect 53281 491947 53347 491950
rect 92841 491602 92907 491605
rect 104249 491602 104315 491605
rect 92841 491600 104315 491602
rect 92841 491544 92846 491600
rect 92902 491544 104254 491600
rect 104310 491544 104315 491600
rect 92841 491542 104315 491544
rect 92841 491539 92907 491542
rect 104249 491539 104315 491542
rect 97809 491466 97875 491469
rect 109534 491466 109540 491468
rect 97809 491464 109540 491466
rect 97809 491408 97814 491464
rect 97870 491408 109540 491464
rect 97809 491406 109540 491408
rect 97809 491403 97875 491406
rect 109534 491404 109540 491406
rect 109604 491404 109610 491468
rect 99281 491330 99347 491333
rect 111006 491330 111012 491332
rect 99281 491328 111012 491330
rect 99281 491272 99286 491328
rect 99342 491272 111012 491328
rect 99281 491270 111012 491272
rect 99281 491267 99347 491270
rect 111006 491268 111012 491270
rect 111076 491268 111082 491332
rect 92013 490650 92079 490653
rect 99414 490650 99420 490652
rect 92013 490648 99420 490650
rect 92013 490592 92018 490648
rect 92074 490592 99420 490648
rect 92013 490590 99420 490592
rect 92013 490587 92079 490590
rect 99414 490588 99420 490590
rect 99484 490588 99490 490652
rect 59118 490452 59124 490516
rect 59188 490514 59194 490516
rect 80881 490514 80947 490517
rect 59188 490512 80947 490514
rect 59188 490456 80886 490512
rect 80942 490456 80947 490512
rect 59188 490454 80947 490456
rect 59188 490452 59194 490454
rect 80881 490451 80947 490454
rect 95141 490514 95207 490517
rect 110321 490514 110387 490517
rect 95141 490512 110387 490514
rect 95141 490456 95146 490512
rect 95202 490456 110326 490512
rect 110382 490456 110387 490512
rect 95141 490454 110387 490456
rect 95141 490451 95207 490454
rect 110321 490451 110387 490454
rect 84837 490106 84903 490109
rect 115974 490106 115980 490108
rect 84837 490104 115980 490106
rect 84837 490048 84842 490104
rect 84898 490048 115980 490104
rect 84837 490046 115980 490048
rect 84837 490043 84903 490046
rect 115974 490044 115980 490046
rect 116044 490044 116050 490108
rect 69749 489970 69815 489973
rect 69749 489968 70226 489970
rect 69749 489912 69754 489968
rect 69810 489912 70226 489968
rect 69749 489910 70226 489912
rect 69749 489907 69815 489910
rect 70166 489804 70226 489910
rect 98494 489908 98500 489972
rect 98564 489970 98570 489972
rect 100109 489970 100175 489973
rect 98564 489968 100175 489970
rect 98564 489912 100114 489968
rect 100170 489912 100175 489968
rect 98564 489910 100175 489912
rect 98564 489908 98570 489910
rect 100109 489907 100175 489910
rect 101857 489970 101923 489973
rect 101990 489970 101996 489972
rect 101857 489968 101996 489970
rect 101857 489912 101862 489968
rect 101918 489912 101996 489968
rect 101857 489910 101996 489912
rect 101857 489907 101923 489910
rect 101990 489908 101996 489910
rect 102060 489908 102066 489972
rect 122782 489908 122788 489972
rect 122852 489970 122858 489972
rect 123109 489970 123175 489973
rect 122852 489968 123175 489970
rect 122852 489912 123114 489968
rect 123170 489912 123175 489968
rect 122852 489910 123175 489912
rect 122852 489908 122858 489910
rect 123109 489907 123175 489910
rect 99281 489290 99347 489293
rect 99281 489288 109050 489290
rect 99281 489232 99286 489288
rect 99342 489232 109050 489288
rect 99281 489230 109050 489232
rect 99281 489227 99347 489230
rect 55070 489092 55076 489156
rect 55140 489154 55146 489156
rect 69841 489154 69907 489157
rect 55140 489152 69907 489154
rect 55140 489096 69846 489152
rect 69902 489096 69907 489152
rect 55140 489094 69907 489096
rect 55140 489092 55146 489094
rect 69841 489091 69907 489094
rect -960 488596 480 488836
rect 99790 488610 99850 488988
rect 108990 488746 109050 489230
rect 114461 488746 114527 488749
rect 108990 488744 114527 488746
rect 108990 488688 114466 488744
rect 114522 488688 114527 488744
rect 108990 488686 114527 488688
rect 114461 488683 114527 488686
rect 99790 488550 115858 488610
rect 115798 488476 115858 488550
rect 115790 488474 115796 488476
rect 115668 488414 115796 488474
rect 115790 488412 115796 488414
rect 115860 488474 115866 488476
rect 120165 488474 120231 488477
rect 115860 488472 120231 488474
rect 115860 488416 120170 488472
rect 120226 488416 120231 488472
rect 115860 488414 120231 488416
rect 115860 488412 115866 488414
rect 120165 488411 120231 488414
rect 100109 488338 100175 488341
rect 109125 488338 109191 488341
rect 100109 488336 109191 488338
rect 67725 488066 67791 488069
rect 70166 488066 70226 488308
rect 67725 488064 70226 488066
rect 67725 488008 67730 488064
rect 67786 488008 70226 488064
rect 67725 488006 70226 488008
rect 67725 488003 67791 488006
rect 67633 487930 67699 487933
rect 99606 487930 99666 488308
rect 100109 488280 100114 488336
rect 100170 488280 109130 488336
rect 109186 488280 109191 488336
rect 100109 488278 109191 488280
rect 100109 488275 100175 488278
rect 109125 488275 109191 488278
rect 103421 487930 103487 487933
rect 67633 487928 70226 487930
rect 67633 487872 67638 487928
rect 67694 487872 70226 487928
rect 67633 487870 70226 487872
rect 99606 487928 103487 487930
rect 99606 487872 103426 487928
rect 103482 487872 103487 487928
rect 99606 487870 103487 487872
rect 67633 487867 67699 487870
rect 70166 487764 70226 487870
rect 103421 487867 103487 487870
rect 99606 487386 99666 487628
rect 103329 487386 103395 487389
rect 99606 487384 103395 487386
rect 99606 487328 103334 487384
rect 103390 487328 103395 487384
rect 99606 487326 103395 487328
rect 103329 487323 103395 487326
rect 69054 486508 69060 486572
rect 69124 486570 69130 486572
rect 69197 486570 69263 486573
rect 70166 486570 70226 486948
rect 99606 486706 99666 486948
rect 103421 486706 103487 486709
rect 99606 486704 103487 486706
rect 99606 486648 103426 486704
rect 103482 486648 103487 486704
rect 99606 486646 103487 486648
rect 103421 486643 103487 486646
rect 106457 486570 106523 486573
rect 69124 486568 70226 486570
rect 69124 486512 69202 486568
rect 69258 486512 70226 486568
rect 69124 486510 70226 486512
rect 99790 486568 109050 486570
rect 99790 486512 106462 486568
rect 106518 486512 109050 486568
rect 99790 486510 109050 486512
rect 69124 486508 69130 486510
rect 69197 486507 69263 486510
rect 99790 486404 99850 486510
rect 106457 486507 106523 486510
rect 108990 486434 109050 486510
rect 118918 486434 118924 486436
rect 108990 486374 118924 486434
rect 118918 486372 118924 486374
rect 118988 486372 118994 486436
rect 67633 485890 67699 485893
rect 70166 485890 70226 486268
rect 67633 485888 70226 485890
rect 67633 485832 67638 485888
rect 67694 485832 70226 485888
rect 67633 485830 70226 485832
rect 67633 485827 67699 485830
rect 67633 485210 67699 485213
rect 70166 485210 70226 485588
rect 99790 485346 99850 485588
rect 102317 485346 102383 485349
rect 99790 485344 102383 485346
rect 99790 485288 102322 485344
rect 102378 485288 102383 485344
rect 99790 485286 102383 485288
rect 102317 485283 102383 485286
rect 67633 485208 70226 485210
rect 67633 485152 67638 485208
rect 67694 485152 70226 485208
rect 67633 485150 70226 485152
rect 67633 485147 67699 485150
rect 111742 485012 111748 485076
rect 111812 485074 111818 485076
rect 112161 485074 112227 485077
rect 113081 485074 113147 485077
rect 111812 485072 113147 485074
rect 111812 485016 112166 485072
rect 112222 485016 113086 485072
rect 113142 485016 113147 485072
rect 111812 485014 113147 485016
rect 111812 485012 111818 485014
rect 112161 485011 112227 485014
rect 113081 485011 113147 485014
rect 115606 485012 115612 485076
rect 115676 485074 115682 485076
rect 131113 485074 131179 485077
rect 115676 485072 131179 485074
rect 115676 485016 131118 485072
rect 131174 485016 131179 485072
rect 115676 485014 131179 485016
rect 115676 485012 115682 485014
rect 131113 485011 131179 485014
rect 68737 484666 68803 484669
rect 70166 484666 70226 484908
rect 70342 484666 70348 484668
rect 68737 484664 70348 484666
rect 68737 484608 68742 484664
rect 68798 484608 70348 484664
rect 68737 484606 70348 484608
rect 68737 484603 68803 484606
rect 70342 484604 70348 484606
rect 70412 484604 70418 484668
rect 99790 484530 99850 484908
rect 580349 484666 580415 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 99790 484470 113098 484530
rect 583520 484516 584960 484606
rect 113038 484394 113098 484470
rect 117313 484394 117379 484397
rect 129825 484394 129891 484397
rect 113038 484392 129891 484394
rect 113038 484336 117318 484392
rect 117374 484336 129830 484392
rect 129886 484336 129891 484392
rect 113038 484334 129891 484336
rect 117313 484331 117379 484334
rect 129825 484331 129891 484334
rect 67633 483714 67699 483717
rect 70166 483714 70226 484228
rect 102317 483850 102383 483853
rect 67633 483712 70226 483714
rect 67633 483656 67638 483712
rect 67694 483656 70226 483712
rect 99790 483848 102383 483850
rect 99790 483792 102322 483848
rect 102378 483792 102383 483848
rect 99790 483790 102383 483792
rect 99790 483684 99850 483790
rect 102317 483787 102383 483790
rect 67633 483654 70226 483656
rect 67633 483651 67699 483654
rect 99790 483110 100034 483170
rect 99790 483004 99850 483110
rect 99974 482898 100034 483110
rect 102317 482898 102383 482901
rect 99974 482896 102383 482898
rect 68686 482564 68692 482628
rect 68756 482626 68762 482628
rect 69289 482626 69355 482629
rect 70350 482626 70410 482868
rect 99974 482840 102322 482896
rect 102378 482840 102383 482896
rect 99974 482838 102383 482840
rect 102317 482835 102383 482838
rect 102409 482626 102475 482629
rect 68756 482624 70410 482626
rect 68756 482568 69294 482624
rect 69350 482568 70410 482624
rect 68756 482566 70410 482568
rect 99790 482624 102475 482626
rect 99790 482568 102414 482624
rect 102470 482568 102475 482624
rect 99790 482566 102475 482568
rect 68756 482564 68762 482566
rect 69289 482563 69355 482566
rect 68093 482490 68159 482493
rect 69381 482490 69447 482493
rect 68093 482488 70226 482490
rect 68093 482432 68098 482488
rect 68154 482432 69386 482488
rect 69442 482432 70226 482488
rect 68093 482430 70226 482432
rect 68093 482427 68159 482430
rect 69381 482427 69447 482430
rect 70166 482324 70226 482430
rect 99790 482324 99850 482566
rect 102409 482563 102475 482566
rect 99790 481750 100034 481810
rect 99790 481644 99850 481750
rect 99974 481538 100034 481750
rect 102317 481538 102383 481541
rect 99974 481536 102383 481538
rect 68553 481130 68619 481133
rect 70166 481130 70226 481508
rect 99974 481480 102322 481536
rect 102378 481480 102383 481536
rect 99974 481478 102383 481480
rect 102317 481475 102383 481478
rect 102409 481266 102475 481269
rect 68553 481128 70226 481130
rect 68553 481072 68558 481128
rect 68614 481072 70226 481128
rect 68553 481070 70226 481072
rect 99790 481264 102475 481266
rect 99790 481208 102414 481264
rect 102470 481208 102475 481264
rect 99790 481206 102475 481208
rect 68553 481067 68619 481070
rect 99790 480964 99850 481206
rect 102409 481203 102475 481206
rect 65926 480524 65932 480588
rect 65996 480586 66002 480588
rect 67357 480586 67423 480589
rect 70350 480586 70410 480828
rect 65996 480584 70410 480586
rect 65996 480528 67362 480584
rect 67418 480528 70410 480584
rect 65996 480526 70410 480528
rect 65996 480524 66002 480526
rect 67357 480523 67423 480526
rect 69982 480210 70226 480270
rect 67633 480178 67699 480181
rect 69982 480178 70042 480210
rect 67633 480176 70042 480178
rect 67633 480120 67638 480176
rect 67694 480120 70042 480176
rect 70166 480148 70226 480210
rect 67633 480118 70042 480120
rect 67633 480115 67699 480118
rect 67725 479906 67791 479909
rect 99606 479906 99666 480148
rect 102317 479906 102383 479909
rect 67725 479904 70226 479906
rect 67725 479848 67730 479904
rect 67786 479848 70226 479904
rect 67725 479846 70226 479848
rect 99606 479904 102383 479906
rect 99606 479848 102322 479904
rect 102378 479848 102383 479904
rect 99606 479846 102383 479848
rect 67725 479843 67791 479846
rect 70166 479604 70226 479846
rect 102317 479843 102383 479846
rect 99790 478954 99850 479468
rect 101949 478954 102015 478957
rect 112294 478954 112300 478956
rect 99790 478952 112300 478954
rect 99790 478896 101954 478952
rect 102010 478896 112300 478952
rect 99790 478894 112300 478896
rect 101949 478891 102015 478894
rect 112294 478892 112300 478894
rect 112364 478892 112370 478956
rect 66110 478484 66116 478548
rect 66180 478546 66186 478548
rect 70350 478546 70410 478788
rect 66180 478486 70410 478546
rect 66180 478484 66186 478486
rect 103421 478138 103487 478141
rect 106406 478138 106412 478140
rect 103421 478136 106412 478138
rect 99790 477866 99850 478108
rect 103421 478080 103426 478136
rect 103482 478080 106412 478136
rect 103421 478078 106412 478080
rect 103421 478075 103487 478078
rect 106406 478076 106412 478078
rect 106476 478076 106482 478140
rect 102409 477866 102475 477869
rect 99790 477864 102475 477866
rect 99790 477808 102414 477864
rect 102470 477808 102475 477864
rect 99790 477806 102475 477808
rect 102409 477803 102475 477806
rect 61694 477396 61700 477460
rect 61764 477458 61770 477460
rect 64597 477458 64663 477461
rect 67725 477458 67791 477461
rect 61764 477456 67791 477458
rect 61764 477400 64602 477456
rect 64658 477400 67730 477456
rect 67786 477400 67791 477456
rect 116025 477458 116091 477461
rect 117078 477458 117084 477460
rect 116025 477456 117084 477458
rect 61764 477398 67791 477400
rect 61764 477396 61770 477398
rect 64597 477395 64663 477398
rect 67725 477395 67791 477398
rect 68369 477050 68435 477053
rect 68829 477050 68895 477053
rect 70166 477050 70226 477428
rect 68369 477048 70226 477050
rect 68369 476992 68374 477048
rect 68430 476992 68834 477048
rect 68890 476992 70226 477048
rect 68369 476990 70226 476992
rect 99790 477050 99850 477428
rect 116025 477400 116030 477456
rect 116086 477400 117084 477456
rect 116025 477398 117084 477400
rect 116025 477395 116091 477398
rect 117078 477396 117084 477398
rect 117148 477458 117154 477460
rect 132493 477458 132559 477461
rect 117148 477456 132559 477458
rect 117148 477400 132498 477456
rect 132554 477400 132559 477456
rect 117148 477398 132559 477400
rect 117148 477396 117154 477398
rect 132493 477395 132559 477398
rect 102501 477050 102567 477053
rect 99790 477048 102567 477050
rect 99790 476992 102506 477048
rect 102562 476992 102567 477048
rect 99790 476990 102567 476992
rect 68369 476987 68435 476990
rect 68829 476987 68895 476990
rect 102501 476987 102567 476990
rect 67633 476370 67699 476373
rect 70534 476370 70594 476748
rect 99790 476506 99850 476748
rect 102317 476506 102383 476509
rect 99790 476504 102383 476506
rect 99790 476448 102322 476504
rect 102378 476448 102383 476504
rect 99790 476446 102383 476448
rect 102317 476443 102383 476446
rect 67633 476368 70594 476370
rect 67633 476312 67638 476368
rect 67694 476312 70594 476368
rect 67633 476310 70594 476312
rect 99465 476370 99531 476373
rect 100661 476370 100727 476373
rect 99465 476368 100727 476370
rect 99465 476312 99470 476368
rect 99526 476312 100666 476368
rect 100722 476312 100727 476368
rect 99465 476310 100727 476312
rect 67633 476307 67699 476310
rect 99465 476307 99531 476310
rect 67725 476234 67791 476237
rect 67725 476232 70042 476234
rect 67725 476176 67730 476232
rect 67786 476176 70042 476232
rect 99790 476204 99850 476310
rect 100661 476307 100727 476310
rect 67725 476174 70042 476176
rect 67725 476171 67791 476174
rect 69982 476130 70042 476174
rect 69982 476070 70226 476130
rect 70166 476068 70226 476070
rect 115933 475962 115999 475965
rect 118734 475962 118740 475964
rect 115933 475960 118740 475962
rect 115933 475904 115938 475960
rect 115994 475904 118740 475960
rect 115933 475902 118740 475904
rect 115933 475899 115999 475902
rect 118734 475900 118740 475902
rect 118804 475900 118810 475964
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 67633 475690 67699 475693
rect 102317 475690 102383 475693
rect 67633 475688 70226 475690
rect 67633 475632 67638 475688
rect 67694 475632 70226 475688
rect 67633 475630 70226 475632
rect 67633 475627 67699 475630
rect 70166 475524 70226 475630
rect 99790 475688 102383 475690
rect 99790 475632 102322 475688
rect 102378 475632 102383 475688
rect 99790 475630 102383 475632
rect 99790 475524 99850 475630
rect 102317 475627 102383 475630
rect 102409 475146 102475 475149
rect 99790 475144 102475 475146
rect 99790 475088 102414 475144
rect 102470 475088 102475 475144
rect 99790 475086 102475 475088
rect 67633 475010 67699 475013
rect 67633 475008 70226 475010
rect 67633 474952 67638 475008
rect 67694 474952 70226 475008
rect 67633 474950 70226 474952
rect 67633 474947 67699 474950
rect 70166 474844 70226 474950
rect 99790 474844 99850 475086
rect 102409 475083 102475 475086
rect 67633 474330 67699 474333
rect 102317 474330 102383 474333
rect 67633 474328 70226 474330
rect 67633 474272 67638 474328
rect 67694 474272 70226 474328
rect 67633 474270 70226 474272
rect 67633 474267 67699 474270
rect 70166 474164 70226 474270
rect 99790 474328 102383 474330
rect 99790 474272 102322 474328
rect 102378 474272 102383 474328
rect 99790 474270 102383 474272
rect 99790 474164 99850 474270
rect 102317 474267 102383 474270
rect 33041 474058 33107 474061
rect 66662 474058 66668 474060
rect 33041 474056 66668 474058
rect 33041 474000 33046 474056
rect 33102 474000 66668 474056
rect 33041 473998 66668 474000
rect 33041 473995 33107 473998
rect 66662 473996 66668 473998
rect 66732 473996 66738 474060
rect 102501 474058 102567 474061
rect 117998 474058 118004 474060
rect 102501 474056 118004 474058
rect 102501 474000 102506 474056
rect 102562 474000 118004 474056
rect 102501 473998 118004 474000
rect 102501 473995 102567 473998
rect 117998 473996 118004 473998
rect 118068 474058 118074 474060
rect 135345 474058 135411 474061
rect 118068 474056 135411 474058
rect 118068 474000 135350 474056
rect 135406 474000 135411 474056
rect 118068 473998 135411 474000
rect 118068 473996 118074 473998
rect 135345 473995 135411 473998
rect 66662 473724 66668 473788
rect 66732 473786 66738 473788
rect 66732 473726 70226 473786
rect 66732 473724 66738 473726
rect 70166 473484 70226 473726
rect 102317 472970 102383 472973
rect 99790 472968 102383 472970
rect 99790 472912 102322 472968
rect 102378 472912 102383 472968
rect 99790 472910 102383 472912
rect 99790 472804 99850 472910
rect 102317 472907 102383 472910
rect 103421 472426 103487 472429
rect 99790 472424 103487 472426
rect 99790 472368 103426 472424
rect 103482 472368 103487 472424
rect 99790 472366 103487 472368
rect 67633 472290 67699 472293
rect 67633 472288 70226 472290
rect 67633 472232 67638 472288
rect 67694 472232 70226 472288
rect 67633 472230 70226 472232
rect 67633 472227 67699 472230
rect 70166 472124 70226 472230
rect 99790 472124 99850 472366
rect 103421 472363 103487 472366
rect 102317 471746 102383 471749
rect 99790 471744 102383 471746
rect 99790 471688 102322 471744
rect 102378 471688 102383 471744
rect 99790 471686 102383 471688
rect 99790 471444 99850 471686
rect 102317 471683 102383 471686
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 68870 471004 68876 471068
rect 68940 471066 68946 471068
rect 70350 471066 70410 471308
rect 103421 471202 103487 471205
rect 104934 471202 104940 471204
rect 103421 471200 104940 471202
rect 103421 471144 103426 471200
rect 103482 471144 104940 471200
rect 103421 471142 104940 471144
rect 103421 471139 103487 471142
rect 104934 471140 104940 471142
rect 105004 471202 105010 471204
rect 151813 471202 151879 471205
rect 105004 471200 151879 471202
rect 105004 471144 151818 471200
rect 151874 471144 151879 471200
rect 105004 471142 151879 471144
rect 105004 471140 105010 471142
rect 151813 471139 151879 471142
rect 102409 471066 102475 471069
rect 68940 471006 70410 471066
rect 99790 471064 102475 471066
rect 99790 471008 102414 471064
rect 102470 471008 102475 471064
rect 99790 471006 102475 471008
rect 68940 471004 68946 471006
rect 67633 470930 67699 470933
rect 67633 470928 70226 470930
rect 67633 470872 67638 470928
rect 67694 470872 70226 470928
rect 67633 470870 70226 470872
rect 67633 470867 67699 470870
rect 70166 470764 70226 470870
rect 99790 470764 99850 471006
rect 102409 471003 102475 471006
rect 67725 470386 67791 470389
rect 67725 470384 70226 470386
rect 67725 470328 67730 470384
rect 67786 470328 70226 470384
rect 67725 470326 70226 470328
rect 67725 470323 67791 470326
rect 70166 470084 70226 470326
rect 103421 470250 103487 470253
rect 99790 470248 103487 470250
rect 99790 470192 103426 470248
rect 103482 470192 103487 470248
rect 99790 470190 103487 470192
rect 99790 470084 99850 470190
rect 103421 470187 103487 470190
rect 67633 469706 67699 469709
rect 102777 469706 102843 469709
rect 67633 469704 70226 469706
rect 67633 469648 67638 469704
rect 67694 469648 70226 469704
rect 67633 469646 70226 469648
rect 67633 469643 67699 469646
rect 70166 469404 70226 469646
rect 99790 469704 102843 469706
rect 99790 469648 102782 469704
rect 102838 469648 102843 469704
rect 99790 469646 102843 469648
rect 99790 469404 99850 469646
rect 102777 469643 102843 469646
rect 67633 469026 67699 469029
rect 68921 469026 68987 469029
rect 67633 469024 70226 469026
rect 67633 468968 67638 469024
rect 67694 468968 68926 469024
rect 68982 468968 70226 469024
rect 67633 468966 70226 468968
rect 67633 468963 67699 468966
rect 68921 468963 68987 468966
rect 70166 468724 70226 468966
rect 102317 468890 102383 468893
rect 99790 468888 102383 468890
rect 99790 468832 102322 468888
rect 102378 468832 102383 468888
rect 99790 468830 102383 468832
rect 99790 468724 99850 468830
rect 102317 468827 102383 468830
rect 67633 468210 67699 468213
rect 67633 468208 70226 468210
rect 67633 468152 67638 468208
rect 67694 468152 70226 468208
rect 67633 468150 70226 468152
rect 67633 468147 67699 468150
rect 70166 468044 70226 468150
rect 105486 467876 105492 467940
rect 105556 467938 105562 467940
rect 109125 467938 109191 467941
rect 105556 467936 109191 467938
rect 105556 467880 109130 467936
rect 109186 467880 109191 467936
rect 105556 467878 109191 467880
rect 105556 467876 105562 467878
rect 109125 467875 109191 467878
rect 63217 467802 63283 467805
rect 64638 467802 64644 467804
rect 63217 467800 64644 467802
rect 63217 467744 63222 467800
rect 63278 467744 64644 467800
rect 63217 467742 64644 467744
rect 63217 467739 63283 467742
rect 64638 467740 64644 467742
rect 64708 467740 64714 467804
rect 64638 467196 64644 467260
rect 64708 467258 64714 467260
rect 64708 467198 70226 467258
rect 64708 467196 64714 467198
rect 70166 466684 70226 467198
rect 99790 466986 99850 467228
rect 102777 466986 102843 466989
rect 99790 466984 102843 466986
rect 99790 466928 102782 466984
rect 102838 466928 102843 466984
rect 99790 466926 102843 466928
rect 102777 466923 102843 466926
rect 103421 466850 103487 466853
rect 99790 466848 103487 466850
rect 99790 466792 103426 466848
rect 103482 466792 103487 466848
rect 99790 466790 103487 466792
rect 99790 466684 99850 466790
rect 103421 466787 103487 466790
rect 99966 466244 99972 466308
rect 100036 466306 100042 466308
rect 111977 466306 112043 466309
rect 100036 466304 112043 466306
rect 100036 466248 111982 466304
rect 112038 466248 112043 466304
rect 100036 466246 112043 466248
rect 100036 466244 100042 466246
rect 111977 466243 112043 466246
rect 102317 466170 102383 466173
rect 99790 466168 102383 466170
rect 99790 466112 102322 466168
rect 102378 466112 102383 466168
rect 99790 466110 102383 466112
rect 99790 466004 99850 466110
rect 102317 466107 102383 466110
rect 67633 465626 67699 465629
rect 70350 465626 70410 465868
rect 103421 465762 103487 465765
rect 107694 465762 107700 465764
rect 103421 465760 107700 465762
rect 103421 465704 103426 465760
rect 103482 465704 107700 465760
rect 103421 465702 107700 465704
rect 103421 465699 103487 465702
rect 107694 465700 107700 465702
rect 107764 465700 107770 465764
rect 67633 465624 70410 465626
rect 67633 465568 67638 465624
rect 67694 465568 70410 465624
rect 67633 465566 70410 465568
rect 67633 465563 67699 465566
rect 67633 465490 67699 465493
rect 103421 465490 103487 465493
rect 67633 465488 70226 465490
rect 67633 465432 67638 465488
rect 67694 465432 70226 465488
rect 67633 465430 70226 465432
rect 67633 465427 67699 465430
rect 70166 465324 70226 465430
rect 99790 465488 103487 465490
rect 99790 465432 103426 465488
rect 103482 465432 103487 465488
rect 99790 465430 103487 465432
rect 99790 465324 99850 465430
rect 103421 465427 103487 465430
rect 67633 464810 67699 464813
rect 102409 464810 102475 464813
rect 67633 464808 70226 464810
rect 67633 464752 67638 464808
rect 67694 464752 70226 464808
rect 67633 464750 70226 464752
rect 67633 464747 67699 464750
rect 70166 464644 70226 464750
rect 99790 464808 102475 464810
rect 99790 464752 102414 464808
rect 102470 464752 102475 464808
rect 99790 464750 102475 464752
rect 99790 464644 99850 464750
rect 102409 464747 102475 464750
rect 67725 464266 67791 464269
rect 102317 464266 102383 464269
rect 67725 464264 70226 464266
rect 67725 464208 67730 464264
rect 67786 464208 70226 464264
rect 67725 464206 70226 464208
rect 67725 464203 67791 464206
rect 70166 463964 70226 464206
rect 99606 464264 102383 464266
rect 99606 464208 102322 464264
rect 102378 464208 102383 464264
rect 99606 464206 102383 464208
rect 99606 463964 99666 464206
rect 102317 464203 102383 464206
rect 61377 463586 61443 463589
rect 61878 463586 61884 463588
rect 61377 463584 61884 463586
rect 61377 463528 61382 463584
rect 61438 463528 61884 463584
rect 61377 463526 61884 463528
rect 61377 463523 61443 463526
rect 61878 463524 61884 463526
rect 61948 463524 61954 463588
rect 116526 463524 116532 463588
rect 116596 463586 116602 463588
rect 121637 463586 121703 463589
rect 116596 463584 121703 463586
rect 116596 463528 121642 463584
rect 121698 463528 121703 463584
rect 116596 463526 121703 463528
rect 116596 463524 116602 463526
rect 121637 463523 121703 463526
rect 102317 463450 102383 463453
rect 99790 463448 102383 463450
rect 99790 463392 102322 463448
rect 102378 463392 102383 463448
rect 99790 463390 102383 463392
rect 99790 463284 99850 463390
rect 102317 463387 102383 463390
rect 67633 462906 67699 462909
rect 70350 462906 70410 463148
rect 67633 462904 70410 462906
rect 67633 462848 67638 462904
rect 67694 462848 70410 462904
rect 67633 462846 70410 462848
rect 67633 462843 67699 462846
rect -960 462634 480 462724
rect 64830 462710 70226 462770
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 61377 462362 61443 462365
rect 64830 462362 64890 462710
rect 70166 462604 70226 462710
rect 61377 462360 64890 462362
rect 61377 462304 61382 462360
rect 61438 462304 64890 462360
rect 61377 462302 64890 462304
rect 61377 462299 61443 462302
rect 102317 462090 102383 462093
rect 99790 462088 102383 462090
rect 99790 462032 102322 462088
rect 102378 462032 102383 462088
rect 99790 462030 102383 462032
rect 99790 461924 99850 462030
rect 102317 462027 102383 462030
rect 102726 461484 102732 461548
rect 102796 461546 102802 461548
rect 117497 461546 117563 461549
rect 102796 461544 117563 461546
rect 102796 461488 117502 461544
rect 117558 461488 117563 461544
rect 102796 461486 117563 461488
rect 102796 461484 102802 461486
rect 117497 461483 117563 461486
rect 66069 461410 66135 461413
rect 102317 461410 102383 461413
rect 66069 461408 70226 461410
rect 66069 461352 66074 461408
rect 66130 461352 70226 461408
rect 66069 461350 70226 461352
rect 66069 461347 66135 461350
rect 70166 461244 70226 461350
rect 99790 461408 102383 461410
rect 99790 461352 102322 461408
rect 102378 461352 102383 461408
rect 99790 461350 102383 461352
rect 99790 461244 99850 461350
rect 102317 461347 102383 461350
rect 60590 460940 60596 461004
rect 60660 461002 60666 461004
rect 66069 461002 66135 461005
rect 60660 461000 66135 461002
rect 60660 460944 66074 461000
rect 66130 460944 66135 461000
rect 60660 460942 66135 460944
rect 60660 460940 60666 460942
rect 66069 460939 66135 460942
rect 67633 460730 67699 460733
rect 67633 460728 70226 460730
rect 67633 460672 67638 460728
rect 67694 460672 70226 460728
rect 67633 460670 70226 460672
rect 67633 460667 67699 460670
rect 70166 460564 70226 460670
rect 67725 460186 67791 460189
rect 99790 460186 99850 460428
rect 102869 460186 102935 460189
rect 67725 460184 70226 460186
rect 67725 460128 67730 460184
rect 67786 460128 70226 460184
rect 67725 460126 70226 460128
rect 99790 460184 102935 460186
rect 99790 460128 102874 460184
rect 102930 460128 102935 460184
rect 99790 460126 102935 460128
rect 67725 460123 67791 460126
rect 70166 459884 70226 460126
rect 102869 460123 102935 460126
rect 115933 460186 115999 460189
rect 127249 460186 127315 460189
rect 115933 460184 127315 460186
rect 115933 460128 115938 460184
rect 115994 460128 127254 460184
rect 127310 460128 127315 460184
rect 115933 460126 127315 460128
rect 115933 460123 115999 460126
rect 127249 460123 127315 460126
rect 102317 460050 102383 460053
rect 99790 460048 102383 460050
rect 99790 459992 102322 460048
rect 102378 459992 102383 460048
rect 99790 459990 102383 459992
rect 99790 459884 99850 459990
rect 102317 459987 102383 459990
rect 114645 459778 114711 459781
rect 115933 459778 115999 459781
rect 114645 459776 115999 459778
rect 114645 459720 114650 459776
rect 114706 459720 115938 459776
rect 115994 459720 115999 459776
rect 114645 459718 115999 459720
rect 114645 459715 114711 459718
rect 115933 459715 115999 459718
rect 115790 459580 115796 459644
rect 115860 459642 115866 459644
rect 117497 459642 117563 459645
rect 115860 459640 117563 459642
rect 115860 459584 117502 459640
rect 117558 459584 117563 459640
rect 115860 459582 117563 459584
rect 115860 459580 115866 459582
rect 117497 459579 117563 459582
rect 67265 459506 67331 459509
rect 67265 459504 70226 459506
rect 67265 459448 67270 459504
rect 67326 459448 70226 459504
rect 67265 459446 70226 459448
rect 67265 459443 67331 459446
rect 70166 459204 70226 459446
rect 102317 459370 102383 459373
rect 99790 459368 102383 459370
rect 99790 459312 102322 459368
rect 102378 459312 102383 459368
rect 99790 459310 102383 459312
rect 99790 459204 99850 459310
rect 102317 459307 102383 459310
rect 67633 458826 67699 458829
rect 67633 458824 70226 458826
rect 67633 458768 67638 458824
rect 67694 458768 70226 458824
rect 67633 458766 70226 458768
rect 67633 458763 67699 458766
rect 70166 458524 70226 458766
rect 102409 458690 102475 458693
rect 99790 458688 102475 458690
rect 99790 458632 102414 458688
rect 102470 458632 102475 458688
rect 99790 458630 102475 458632
rect 99790 458524 99850 458630
rect 102409 458627 102475 458630
rect 115197 458282 115263 458285
rect 115606 458282 115612 458284
rect 115197 458280 115612 458282
rect 115197 458224 115202 458280
rect 115258 458224 115612 458280
rect 115197 458222 115612 458224
rect 115197 458219 115263 458222
rect 115606 458220 115612 458222
rect 115676 458220 115682 458284
rect 103513 458146 103579 458149
rect 99790 458144 103579 458146
rect 99790 458088 103518 458144
rect 103574 458088 103579 458144
rect 99790 458086 103579 458088
rect 68093 458010 68159 458013
rect 69197 458010 69263 458013
rect 68093 458008 70226 458010
rect 68093 457952 68098 458008
rect 68154 457952 69202 458008
rect 69258 457952 70226 458008
rect 68093 457950 70226 457952
rect 68093 457947 68159 457950
rect 69197 457947 69263 457950
rect 70166 457844 70226 457950
rect 99790 457844 99850 458086
rect 103513 458083 103579 458086
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect 67633 457466 67699 457469
rect 135437 457466 135503 457469
rect 150433 457466 150499 457469
rect 67633 457464 70226 457466
rect 67633 457408 67638 457464
rect 67694 457408 70226 457464
rect 67633 457406 70226 457408
rect 67633 457403 67699 457406
rect 70166 457164 70226 457406
rect 113130 457464 150499 457466
rect 113130 457408 135442 457464
rect 135498 457408 150438 457464
rect 150494 457408 150499 457464
rect 113130 457406 150499 457408
rect 113130 456922 113190 457406
rect 135437 457403 135503 457406
rect 150433 457403 150499 457406
rect 107702 456862 113190 456922
rect 106089 456786 106155 456789
rect 107702 456786 107762 456862
rect 106089 456784 107762 456786
rect 106089 456728 106094 456784
rect 106150 456728 107762 456784
rect 106089 456726 107762 456728
rect 106089 456723 106155 456726
rect 102409 456650 102475 456653
rect 99790 456648 102475 456650
rect 99790 456592 102414 456648
rect 102470 456592 102475 456648
rect 99790 456590 102475 456592
rect 99790 456484 99850 456590
rect 102409 456587 102475 456590
rect 102225 456106 102291 456109
rect 99606 456104 102291 456106
rect 99606 456048 102230 456104
rect 102286 456048 102291 456104
rect 99606 456046 102291 456048
rect 67633 455970 67699 455973
rect 67633 455968 70226 455970
rect 67633 455912 67638 455968
rect 67694 455912 70226 455968
rect 67633 455910 70226 455912
rect 67633 455907 67699 455910
rect 70166 455804 70226 455910
rect 99606 455804 99666 456046
rect 102225 456043 102291 456046
rect 107561 456106 107627 456109
rect 107878 456106 107884 456108
rect 107561 456104 107884 456106
rect 107561 456048 107566 456104
rect 107622 456048 107884 456104
rect 107561 456046 107884 456048
rect 107561 456043 107627 456046
rect 107878 456044 107884 456046
rect 107948 456106 107954 456108
rect 149053 456106 149119 456109
rect 107948 456104 149119 456106
rect 107948 456048 149058 456104
rect 149114 456048 149119 456104
rect 107948 456046 149119 456048
rect 107948 456044 107954 456046
rect 149053 456043 149119 456046
rect 103513 455426 103579 455429
rect 99790 455424 103579 455426
rect 99790 455368 103518 455424
rect 103574 455368 103579 455424
rect 99790 455366 103579 455368
rect 99790 455124 99850 455366
rect 103513 455363 103579 455366
rect 67633 454610 67699 454613
rect 70166 454610 70226 454988
rect 102225 454746 102291 454749
rect 67633 454608 70226 454610
rect 67633 454552 67638 454608
rect 67694 454552 70226 454608
rect 67633 454550 70226 454552
rect 99790 454744 102291 454746
rect 99790 454688 102230 454744
rect 102286 454688 102291 454744
rect 99790 454686 102291 454688
rect 67633 454547 67699 454550
rect 99790 454444 99850 454686
rect 102225 454683 102291 454686
rect 69105 454066 69171 454069
rect 70350 454066 70410 454308
rect 69105 454064 70410 454066
rect 69105 454008 69110 454064
rect 69166 454008 70410 454064
rect 69105 454006 70410 454008
rect 69105 454003 69171 454006
rect 67725 453930 67791 453933
rect 102225 453930 102291 453933
rect 67725 453928 70226 453930
rect 67725 453872 67730 453928
rect 67786 453872 70226 453928
rect 67725 453870 70226 453872
rect 67725 453867 67791 453870
rect 70166 453764 70226 453870
rect 99790 453928 102291 453930
rect 99790 453872 102230 453928
rect 102286 453872 102291 453928
rect 99790 453870 102291 453872
rect 99790 453764 99850 453870
rect 102225 453867 102291 453870
rect 67633 453250 67699 453253
rect 102225 453250 102291 453253
rect 67633 453248 70226 453250
rect 67633 453192 67638 453248
rect 67694 453192 70226 453248
rect 67633 453190 70226 453192
rect 67633 453187 67699 453190
rect 70166 453084 70226 453190
rect 99790 453248 102291 453250
rect 99790 453192 102230 453248
rect 102286 453192 102291 453248
rect 99790 453190 102291 453192
rect 99790 453084 99850 453190
rect 102225 453187 102291 453190
rect 102225 452570 102291 452573
rect 99790 452568 102291 452570
rect 99790 452512 102230 452568
rect 102286 452512 102291 452568
rect 99790 452510 102291 452512
rect 99790 452404 99850 452510
rect 102225 452507 102291 452510
rect 66989 451890 67055 451893
rect 70166 451890 70226 452268
rect 66989 451888 70226 451890
rect 66989 451832 66994 451888
rect 67050 451832 70226 451888
rect 66989 451830 70226 451832
rect 66989 451827 67055 451830
rect 67725 451346 67791 451349
rect 70350 451346 70410 451588
rect 67725 451344 70410 451346
rect 67725 451288 67730 451344
rect 67786 451288 70410 451344
rect 67725 451286 70410 451288
rect 67725 451283 67791 451286
rect 100845 451210 100911 451213
rect 99790 451208 100911 451210
rect 99790 451152 100850 451208
rect 100906 451152 100911 451208
rect 99790 451150 100911 451152
rect 99790 451044 99850 451150
rect 100845 451147 100911 451150
rect 103513 450666 103579 450669
rect 99790 450664 103579 450666
rect 99790 450608 103518 450664
rect 103574 450608 103579 450664
rect 99790 450606 103579 450608
rect 99790 450364 99850 450606
rect 103513 450603 103579 450606
rect 67633 449986 67699 449989
rect 70166 449986 70226 450228
rect 67633 449984 70226 449986
rect 67633 449928 67638 449984
rect 67694 449928 70226 449984
rect 67633 449926 70226 449928
rect 67633 449923 67699 449926
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 67725 449306 67791 449309
rect 68277 449306 68343 449309
rect 70166 449306 70226 449548
rect 67725 449304 70226 449306
rect 67725 449248 67730 449304
rect 67786 449248 68282 449304
rect 68338 449248 70226 449304
rect 67725 449246 70226 449248
rect 99790 449306 99850 449548
rect 102133 449306 102199 449309
rect 99790 449304 102199 449306
rect 99790 449248 102138 449304
rect 102194 449248 102199 449304
rect 99790 449246 102199 449248
rect 67725 449243 67791 449246
rect 68277 449243 68343 449246
rect 102133 449243 102199 449246
rect 67633 449170 67699 449173
rect 102409 449170 102475 449173
rect 67633 449168 70226 449170
rect 67633 449112 67638 449168
rect 67694 449112 70226 449168
rect 67633 449110 70226 449112
rect 67633 449107 67699 449110
rect 70166 449004 70226 449110
rect 99790 449168 102475 449170
rect 99790 449112 102414 449168
rect 102470 449112 102475 449168
rect 99790 449110 102475 449112
rect 99790 449004 99850 449110
rect 102409 449107 102475 449110
rect 102133 448490 102199 448493
rect 99790 448488 102199 448490
rect 99790 448432 102138 448488
rect 102194 448432 102199 448488
rect 99790 448430 102199 448432
rect 99790 448324 99850 448430
rect 102133 448427 102199 448430
rect 62982 447748 62988 447812
rect 63052 447810 63058 447812
rect 63309 447810 63375 447813
rect 70166 447810 70226 448188
rect 102409 447946 102475 447949
rect 63052 447808 70226 447810
rect 63052 447752 63314 447808
rect 63370 447752 70226 447808
rect 63052 447750 70226 447752
rect 99790 447944 102475 447946
rect 99790 447888 102414 447944
rect 102470 447888 102475 447944
rect 99790 447886 102475 447888
rect 63052 447748 63058 447750
rect 63309 447747 63375 447750
rect 99790 447644 99850 447886
rect 102409 447883 102475 447886
rect 67633 447266 67699 447269
rect 70350 447266 70410 447508
rect 67633 447264 70410 447266
rect 67633 447208 67638 447264
rect 67694 447208 70410 447264
rect 67633 447206 70410 447208
rect 67633 447203 67699 447206
rect 67633 446450 67699 446453
rect 70166 446450 70226 446828
rect 99373 446586 99439 446589
rect 99790 446586 99850 446828
rect 99373 446584 99850 446586
rect 99373 446528 99378 446584
rect 99434 446528 99850 446584
rect 99373 446526 99850 446528
rect 99373 446523 99439 446526
rect 67633 446448 70226 446450
rect 67633 446392 67638 446448
rect 67694 446392 70226 446448
rect 67633 446390 70226 446392
rect 67633 446387 67699 446390
rect 99790 446314 99850 446526
rect 102133 446314 102199 446317
rect 99790 446312 102199 446314
rect 99790 446256 102138 446312
rect 102194 446256 102199 446312
rect 99790 446254 102199 446256
rect 102133 446251 102199 446254
rect 67725 445906 67791 445909
rect 70166 445906 70226 446148
rect 67725 445904 70226 445906
rect 67725 445848 67730 445904
rect 67786 445848 70226 445904
rect 67725 445846 70226 445848
rect 67725 445843 67791 445846
rect 103830 445770 103836 445772
rect 99790 445710 103836 445770
rect 99790 445604 99850 445710
rect 103830 445708 103836 445710
rect 103900 445708 103906 445772
rect 104065 445770 104131 445773
rect 133086 445770 133092 445772
rect 104065 445768 133092 445770
rect 104065 445712 104070 445768
rect 104126 445712 133092 445768
rect 104065 445710 133092 445712
rect 104065 445707 104131 445710
rect 133086 445708 133092 445710
rect 133156 445708 133162 445772
rect 104065 445226 104131 445229
rect 99790 445224 104131 445226
rect 99790 445168 104070 445224
rect 104126 445168 104131 445224
rect 99790 445166 104131 445168
rect 67633 445090 67699 445093
rect 67633 445088 70226 445090
rect 67633 445032 67638 445088
rect 67694 445032 70226 445088
rect 67633 445030 70226 445032
rect 67633 445027 67699 445030
rect 70166 444924 70226 445030
rect 99790 444924 99850 445166
rect 104065 445163 104131 445166
rect 583520 444668 584960 444908
rect 69982 444350 70226 444410
rect 67725 444274 67791 444277
rect 69982 444274 70042 444350
rect 67725 444272 70042 444274
rect 67725 444216 67730 444272
rect 67786 444216 70042 444272
rect 70166 444244 70226 444350
rect 99790 444390 100034 444410
rect 99790 444350 100218 444390
rect 99790 444244 99850 444350
rect 99974 444330 100218 444350
rect 103830 444348 103836 444412
rect 103900 444410 103906 444412
rect 104157 444410 104223 444413
rect 103900 444408 104223 444410
rect 103900 444352 104162 444408
rect 104218 444352 104223 444408
rect 103900 444350 104223 444352
rect 103900 444348 103906 444350
rect 104157 444347 104223 444350
rect 100158 444274 100218 444330
rect 103513 444274 103579 444277
rect 100158 444272 103579 444274
rect 67725 444214 70042 444216
rect 100158 444216 103518 444272
rect 103574 444216 103579 444272
rect 100158 444214 103579 444216
rect 67725 444211 67791 444214
rect 103513 444211 103579 444214
rect 67633 443866 67699 443869
rect 67633 443864 70226 443866
rect 67633 443808 67638 443864
rect 67694 443808 70226 443864
rect 67633 443806 70226 443808
rect 67633 443803 67699 443806
rect 70166 443564 70226 443806
rect 99741 443730 99807 443733
rect 102593 443730 102659 443733
rect 99660 443728 102659 443730
rect 99660 443672 99746 443728
rect 99802 443672 102598 443728
rect 102654 443672 102659 443728
rect 99660 443670 102659 443672
rect 99741 443667 99850 443670
rect 102593 443667 102659 443670
rect 99790 443564 99850 443667
rect 102869 443050 102935 443053
rect 69982 442990 70226 443050
rect 60733 442914 60799 442917
rect 61878 442914 61884 442916
rect 60733 442912 61884 442914
rect 60733 442856 60738 442912
rect 60794 442856 61884 442912
rect 60733 442854 61884 442856
rect 60733 442851 60799 442854
rect 61878 442852 61884 442854
rect 61948 442852 61954 442916
rect 67725 442914 67791 442917
rect 69982 442914 70042 442990
rect 67725 442912 70042 442914
rect 67725 442856 67730 442912
rect 67786 442856 70042 442912
rect 70166 442884 70226 442990
rect 99790 443048 102935 443050
rect 99790 442992 102874 443048
rect 102930 442992 102935 443048
rect 99790 442990 102935 442992
rect 99790 442884 99850 442990
rect 102869 442987 102935 442990
rect 67725 442854 70042 442856
rect 67725 442851 67791 442854
rect 67633 442506 67699 442509
rect 99281 442506 99347 442509
rect 120349 442506 120415 442509
rect 67633 442504 70226 442506
rect 67633 442448 67638 442504
rect 67694 442448 70226 442504
rect 67633 442446 70226 442448
rect 67633 442443 67699 442446
rect 70166 442204 70226 442446
rect 99281 442504 120415 442506
rect 99281 442448 99286 442504
rect 99342 442448 120354 442504
rect 120410 442448 120415 442504
rect 99281 442446 120415 442448
rect 99281 442443 99347 442446
rect 120349 442443 120415 442446
rect 99606 441826 99666 442068
rect 102041 441826 102107 441829
rect 103329 441826 103395 441829
rect 99606 441824 103395 441826
rect 99606 441768 102046 441824
rect 102102 441768 103334 441824
rect 103390 441768 103395 441824
rect 99606 441766 103395 441768
rect 102041 441763 102107 441766
rect 103329 441763 103395 441766
rect 61878 441628 61884 441692
rect 61948 441690 61954 441692
rect 67725 441690 67791 441693
rect 61948 441688 67791 441690
rect 61948 441632 67730 441688
rect 67786 441632 67791 441688
rect 61948 441630 67791 441632
rect 61948 441628 61954 441630
rect 67725 441627 67791 441630
rect 69841 441282 69907 441285
rect 64830 441280 69907 441282
rect 64830 441224 69846 441280
rect 69902 441224 69907 441280
rect 64830 441222 69907 441224
rect 53598 441084 53604 441148
rect 53668 441146 53674 441148
rect 64830 441146 64890 441222
rect 69841 441219 69907 441222
rect 53668 441086 64890 441146
rect 67725 441146 67791 441149
rect 70166 441146 70226 441388
rect 67725 441144 70226 441146
rect 67725 441088 67730 441144
rect 67786 441088 70226 441144
rect 67725 441086 70226 441088
rect 53668 441084 53674 441086
rect 67725 441083 67791 441086
rect 99046 441084 99052 441148
rect 99116 441146 99122 441148
rect 99281 441146 99347 441149
rect 99116 441144 99347 441146
rect 99116 441088 99286 441144
rect 99342 441088 99347 441144
rect 99116 441086 99347 441088
rect 99606 441146 99666 441388
rect 100293 441146 100359 441149
rect 102869 441146 102935 441149
rect 99606 441144 102935 441146
rect 99606 441088 100298 441144
rect 100354 441088 102874 441144
rect 102930 441088 102935 441144
rect 99606 441086 102935 441088
rect 99116 441084 99122 441086
rect 99281 441083 99347 441086
rect 100293 441083 100359 441086
rect 102869 441083 102935 441086
rect 59118 440948 59124 441012
rect 59188 441010 59194 441012
rect 59188 440950 74550 441010
rect 59188 440948 59194 440950
rect 74490 440738 74550 440950
rect 79317 440738 79383 440741
rect 81433 440738 81499 440741
rect 74490 440736 81499 440738
rect 65977 440332 66043 440333
rect 65926 440330 65932 440332
rect 65886 440270 65932 440330
rect 65996 440328 66043 440332
rect 66038 440272 66043 440328
rect 65926 440268 65932 440270
rect 65996 440268 66043 440272
rect 65977 440267 66043 440268
rect 67633 440330 67699 440333
rect 70166 440330 70226 440708
rect 74490 440680 79322 440736
rect 79378 440680 81438 440736
rect 81494 440680 81499 440736
rect 74490 440678 81499 440680
rect 79317 440675 79383 440678
rect 81433 440675 81499 440678
rect 67633 440328 70226 440330
rect 67633 440272 67638 440328
rect 67694 440272 70226 440328
rect 67633 440270 70226 440272
rect 67633 440267 67699 440270
rect 102041 440194 102107 440197
rect 102726 440194 102732 440196
rect 102041 440192 102732 440194
rect 102041 440136 102046 440192
rect 102102 440136 102732 440192
rect 102041 440134 102732 440136
rect 102041 440131 102107 440134
rect 102726 440132 102732 440134
rect 102796 440132 102802 440196
rect 99606 439786 99666 440028
rect 100753 439786 100819 439789
rect 103053 439786 103119 439789
rect 99606 439784 103119 439786
rect 99606 439728 100758 439784
rect 100814 439728 103058 439784
rect 103114 439728 103119 439784
rect 99606 439726 103119 439728
rect 100753 439723 100819 439726
rect 103053 439723 103119 439726
rect 37089 439514 37155 439517
rect 64638 439514 64644 439516
rect 37089 439512 64644 439514
rect 37089 439456 37094 439512
rect 37150 439456 64644 439512
rect 37089 439454 64644 439456
rect 37089 439451 37155 439454
rect 64638 439452 64644 439454
rect 64708 439514 64714 439516
rect 67633 439514 67699 439517
rect 64708 439512 67699 439514
rect 64708 439456 67638 439512
rect 67694 439456 67699 439512
rect 64708 439454 67699 439456
rect 64708 439452 64714 439454
rect 67633 439451 67699 439454
rect 69054 439452 69060 439516
rect 69124 439514 69130 439516
rect 77937 439514 78003 439517
rect 69124 439512 78003 439514
rect 69124 439456 77942 439512
rect 77998 439456 78003 439512
rect 69124 439454 78003 439456
rect 69124 439452 69130 439454
rect 77937 439451 78003 439454
rect 121545 439378 121611 439381
rect 122097 439378 122163 439381
rect 124254 439378 124260 439380
rect 121545 439376 124260 439378
rect 121545 439320 121550 439376
rect 121606 439320 122102 439376
rect 122158 439320 124260 439376
rect 121545 439318 124260 439320
rect 121545 439315 121611 439318
rect 122097 439315 122163 439318
rect 124254 439316 124260 439318
rect 124324 439316 124330 439380
rect 92565 439106 92631 439109
rect 99414 439106 99420 439108
rect 92565 439104 99420 439106
rect 92565 439048 92570 439104
rect 92626 439048 99420 439104
rect 92565 439046 99420 439048
rect 92565 439043 92631 439046
rect 99414 439044 99420 439046
rect 99484 439044 99490 439108
rect 68686 438908 68692 438972
rect 68756 438970 68762 438972
rect 71037 438970 71103 438973
rect 68756 438968 71103 438970
rect 68756 438912 71042 438968
rect 71098 438912 71103 438968
rect 68756 438910 71103 438912
rect 68756 438908 68762 438910
rect 71037 438907 71103 438910
rect 84193 438970 84259 438973
rect 102041 438970 102107 438973
rect 84193 438968 102107 438970
rect 84193 438912 84198 438968
rect 84254 438912 102046 438968
rect 102102 438912 102107 438968
rect 84193 438910 102107 438912
rect 84193 438907 84259 438910
rect 102041 438907 102107 438910
rect 55070 438772 55076 438836
rect 55140 438834 55146 438836
rect 79685 438834 79751 438837
rect 55140 438832 79751 438834
rect 55140 438776 79690 438832
rect 79746 438776 79751 438832
rect 55140 438774 79751 438776
rect 55140 438772 55146 438774
rect 79685 438771 79751 438774
rect 91277 438834 91343 438837
rect 124438 438834 124444 438836
rect 91277 438832 124444 438834
rect 91277 438776 91282 438832
rect 91338 438776 124444 438832
rect 91277 438774 124444 438776
rect 91277 438771 91343 438774
rect 124438 438772 124444 438774
rect 124508 438834 124514 438836
rect 125726 438834 125732 438836
rect 124508 438774 125732 438834
rect 124508 438772 124514 438774
rect 125726 438772 125732 438774
rect 125796 438772 125802 438836
rect 90357 438698 90423 438701
rect 99966 438698 99972 438700
rect 90357 438696 99972 438698
rect 90357 438640 90362 438696
rect 90418 438640 99972 438696
rect 90357 438638 99972 438640
rect 90357 438635 90423 438638
rect 99966 438636 99972 438638
rect 100036 438636 100042 438700
rect 70342 437684 70348 437748
rect 70412 437746 70418 437748
rect 70669 437746 70735 437749
rect 70412 437744 70735 437746
rect 70412 437688 70674 437744
rect 70730 437688 70735 437744
rect 70412 437686 70735 437688
rect 70412 437684 70418 437686
rect 70669 437683 70735 437686
rect 78673 437610 78739 437613
rect 79685 437610 79751 437613
rect 78673 437608 79751 437610
rect 78673 437552 78678 437608
rect 78734 437552 79690 437608
rect 79746 437552 79751 437608
rect 78673 437550 79751 437552
rect 78673 437547 78739 437550
rect 79685 437547 79751 437550
rect 57830 437412 57836 437476
rect 57900 437474 57906 437476
rect 81893 437474 81959 437477
rect 57900 437472 81959 437474
rect 57900 437416 81898 437472
rect 81954 437416 81959 437472
rect 57900 437414 81959 437416
rect 57900 437412 57906 437414
rect 81893 437411 81959 437414
rect -960 436508 480 436748
rect 89621 435978 89687 435981
rect 105486 435978 105492 435980
rect 89621 435976 105492 435978
rect 89621 435920 89626 435976
rect 89682 435920 105492 435976
rect 89621 435918 105492 435920
rect 89621 435915 89687 435918
rect 105486 435916 105492 435918
rect 105556 435916 105562 435980
rect 44030 434556 44036 434620
rect 44100 434618 44106 434620
rect 74533 434618 74599 434621
rect 44100 434616 74599 434618
rect 44100 434560 74538 434616
rect 74594 434560 74599 434616
rect 44100 434558 74599 434560
rect 44100 434556 44106 434558
rect 74533 434555 74599 434558
rect 48078 433196 48084 433260
rect 48148 433258 48154 433260
rect 48957 433258 49023 433261
rect 48148 433256 49023 433258
rect 48148 433200 48962 433256
rect 49018 433200 49023 433256
rect 48148 433198 49023 433200
rect 48148 433196 48154 433198
rect 48957 433195 49023 433198
rect 49325 431898 49391 431901
rect 71773 431898 71839 431901
rect 49325 431896 71839 431898
rect 49325 431840 49330 431896
rect 49386 431840 71778 431896
rect 71834 431840 71839 431896
rect 49325 431838 71839 431840
rect 49325 431835 49391 431838
rect 71773 431835 71839 431838
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 48078 430612 48084 430676
rect 48148 430674 48154 430676
rect 49325 430674 49391 430677
rect 48148 430672 49391 430674
rect 48148 430616 49330 430672
rect 49386 430616 49391 430672
rect 48148 430614 49391 430616
rect 48148 430612 48154 430614
rect 49325 430611 49391 430614
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 93669 404970 93735 404973
rect 128670 404970 128676 404972
rect 93669 404968 128676 404970
rect 93669 404912 93674 404968
rect 93730 404912 128676 404968
rect 93669 404910 128676 404912
rect 93669 404907 93735 404910
rect 128670 404908 128676 404910
rect 128740 404908 128746 404972
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 61694 401644 61700 401708
rect 61764 401706 61770 401708
rect 62021 401706 62087 401709
rect 160737 401706 160803 401709
rect 61764 401704 160803 401706
rect 61764 401648 62026 401704
rect 62082 401648 160742 401704
rect 160798 401648 160803 401704
rect 61764 401646 160803 401648
rect 61764 401644 61770 401646
rect 62021 401643 62087 401646
rect 160737 401643 160803 401646
rect 109534 401236 109540 401300
rect 109604 401298 109610 401300
rect 113817 401298 113883 401301
rect 109604 401296 113883 401298
rect 109604 401240 113822 401296
rect 113878 401240 113883 401296
rect 109604 401238 113883 401240
rect 109604 401236 109610 401238
rect 113817 401235 113883 401238
rect 66110 400284 66116 400348
rect 66180 400346 66186 400348
rect 264237 400346 264303 400349
rect 66180 400344 264303 400346
rect 66180 400288 264242 400344
rect 264298 400288 264303 400344
rect 66180 400286 264303 400288
rect 66180 400284 66186 400286
rect 264237 400283 264303 400286
rect 53598 399604 53604 399668
rect 53668 399666 53674 399668
rect 84193 399666 84259 399669
rect 53668 399664 84259 399666
rect 53668 399608 84198 399664
rect 84254 399608 84259 399664
rect 53668 399606 84259 399608
rect 53668 399604 53674 399606
rect 84193 399603 84259 399606
rect 50838 399468 50844 399532
rect 50908 399530 50914 399532
rect 85113 399530 85179 399533
rect 50908 399528 85179 399530
rect 50908 399472 85118 399528
rect 85174 399472 85179 399528
rect 50908 399470 85179 399472
rect 50908 399468 50914 399470
rect 85113 399467 85179 399470
rect 93761 399530 93827 399533
rect 129774 399530 129780 399532
rect 93761 399528 129780 399530
rect 93761 399472 93766 399528
rect 93822 399472 129780 399528
rect 93761 399470 129780 399472
rect 93761 399467 93827 399470
rect 129774 399468 129780 399470
rect 129844 399468 129850 399532
rect 64781 398850 64847 398853
rect 168414 398850 168420 398852
rect 64781 398848 168420 398850
rect 64781 398792 64786 398848
rect 64842 398792 168420 398848
rect 64781 398790 168420 398792
rect 64781 398787 64847 398790
rect 168414 398788 168420 398790
rect 168484 398788 168490 398852
rect 52310 397972 52316 398036
rect 52380 398034 52386 398036
rect 92473 398034 92539 398037
rect 52380 398032 92539 398034
rect 52380 397976 92478 398032
rect 92534 397976 92539 398032
rect 52380 397974 92539 397976
rect 52380 397972 52386 397974
rect 92473 397971 92539 397974
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 103421 394090 103487 394093
rect 115974 394090 115980 394092
rect 103421 394088 115980 394090
rect 103421 394032 103426 394088
rect 103482 394032 115980 394088
rect 103421 394030 115980 394032
rect 103421 394027 103487 394030
rect 115974 394028 115980 394030
rect 116044 394028 116050 394092
rect 110413 393954 110479 393957
rect 173014 393954 173020 393956
rect 110413 393952 173020 393954
rect 110413 393896 110418 393952
rect 110474 393896 173020 393952
rect 110413 393894 173020 393896
rect 110413 393891 110479 393894
rect 173014 393892 173020 393894
rect 173084 393892 173090 393956
rect 100753 393410 100819 393413
rect 101990 393410 101996 393412
rect 100753 393408 101996 393410
rect 100753 393352 100758 393408
rect 100814 393352 101996 393408
rect 100753 393350 101996 393352
rect 100753 393347 100819 393350
rect 101990 393348 101996 393350
rect 102060 393410 102066 393412
rect 133822 393410 133828 393412
rect 102060 393350 133828 393410
rect 102060 393348 102066 393350
rect 133822 393348 133828 393350
rect 133892 393348 133898 393412
rect 99189 392594 99255 392597
rect 124213 392594 124279 392597
rect 238017 392594 238083 392597
rect 99189 392592 238083 392594
rect 99189 392536 99194 392592
rect 99250 392536 124218 392592
rect 124274 392536 238022 392592
rect 238078 392536 238083 392592
rect 99189 392534 238083 392536
rect 99189 392531 99255 392534
rect 124213 392531 124279 392534
rect 238017 392531 238083 392534
rect 583520 391628 584960 391868
rect 57830 391172 57836 391236
rect 57900 391234 57906 391236
rect 81525 391234 81591 391237
rect 57900 391232 81591 391234
rect 57900 391176 81530 391232
rect 81586 391176 81591 391232
rect 57900 391174 81591 391176
rect 57900 391172 57906 391174
rect 81525 391171 81591 391174
rect 91553 390690 91619 390693
rect 91921 390690 91987 390693
rect 121678 390690 121684 390692
rect 91553 390688 121684 390690
rect 91553 390632 91558 390688
rect 91614 390632 91926 390688
rect 91982 390632 121684 390688
rect 91553 390630 121684 390632
rect 91553 390627 91619 390630
rect 91921 390627 91987 390630
rect 121678 390628 121684 390630
rect 121748 390628 121754 390692
rect 96521 389874 96587 389877
rect 122598 389874 122604 389876
rect 96521 389872 122604 389874
rect 96521 389816 96526 389872
rect 96582 389816 122604 389872
rect 96521 389814 122604 389816
rect 96521 389811 96587 389814
rect 122598 389812 122604 389814
rect 122668 389812 122674 389876
rect 59118 389132 59124 389196
rect 59188 389194 59194 389196
rect 95877 389194 95943 389197
rect 96521 389194 96587 389197
rect 59188 389192 96587 389194
rect 59188 389136 95882 389192
rect 95938 389136 96526 389192
rect 96582 389136 96587 389192
rect 59188 389134 96587 389136
rect 59188 389132 59194 389134
rect 95877 389131 95943 389134
rect 96521 389131 96587 389134
rect 111006 389132 111012 389196
rect 111076 389194 111082 389196
rect 114921 389194 114987 389197
rect 313273 389194 313339 389197
rect 111076 389192 313339 389194
rect 111076 389136 114926 389192
rect 114982 389136 313278 389192
rect 313334 389136 313339 389192
rect 111076 389134 313339 389136
rect 111076 389132 111082 389134
rect 114921 389131 114987 389134
rect 313273 389131 313339 389134
rect 121913 388922 121979 388925
rect 122414 388922 122420 388924
rect 121913 388920 122420 388922
rect 121913 388864 121918 388920
rect 121974 388864 122420 388920
rect 121913 388862 122420 388864
rect 121913 388859 121979 388862
rect 122414 388860 122420 388862
rect 122484 388922 122490 388924
rect 123017 388922 123083 388925
rect 122484 388920 123083 388922
rect 122484 388864 123022 388920
rect 123078 388864 123083 388920
rect 122484 388862 123083 388864
rect 122484 388860 122490 388862
rect 123017 388859 123083 388862
rect 98821 388378 98887 388381
rect 99046 388378 99052 388380
rect 98821 388376 99052 388378
rect 98821 388320 98826 388376
rect 98882 388320 99052 388376
rect 98821 388318 99052 388320
rect 98821 388315 98887 388318
rect 99046 388316 99052 388318
rect 99116 388378 99122 388380
rect 123334 388378 123340 388380
rect 99116 388318 123340 388378
rect 99116 388316 99122 388318
rect 123334 388316 123340 388318
rect 123404 388316 123410 388380
rect 71037 387834 71103 387837
rect 73521 387834 73587 387837
rect 115422 387834 115428 387836
rect 71037 387832 115428 387834
rect 71037 387776 71042 387832
rect 71098 387776 73526 387832
rect 73582 387776 115428 387832
rect 71037 387774 115428 387776
rect 71037 387771 71103 387774
rect 73521 387771 73587 387774
rect 115422 387772 115428 387774
rect 115492 387772 115498 387836
rect 120625 387834 120691 387837
rect 120758 387834 120764 387836
rect 120625 387832 120764 387834
rect 120625 387776 120630 387832
rect 120686 387776 120764 387832
rect 120625 387774 120764 387776
rect 120625 387771 120691 387774
rect 120758 387772 120764 387774
rect 120828 387772 120834 387836
rect 122097 387834 122163 387837
rect 122598 387834 122604 387836
rect 122097 387832 122604 387834
rect 122097 387776 122102 387832
rect 122158 387776 122604 387832
rect 122097 387774 122604 387776
rect 122097 387771 122163 387774
rect 122598 387772 122604 387774
rect 122668 387772 122674 387836
rect 70526 387636 70532 387700
rect 70596 387698 70602 387700
rect 76005 387698 76071 387701
rect 70596 387696 76071 387698
rect 70596 387640 76010 387696
rect 76066 387640 76071 387696
rect 70596 387638 76071 387640
rect 70596 387636 70602 387638
rect 76005 387635 76071 387638
rect 53046 387500 53052 387564
rect 53116 387562 53122 387564
rect 53465 387562 53531 387565
rect 53116 387560 53531 387562
rect 53116 387504 53470 387560
rect 53526 387504 53531 387560
rect 53116 387502 53531 387504
rect 53116 387500 53122 387502
rect 53465 387499 53531 387502
rect 85941 386474 86007 386477
rect 306373 386474 306439 386477
rect 85941 386472 306439 386474
rect 85941 386416 85946 386472
rect 86002 386416 306378 386472
rect 306434 386416 306439 386472
rect 85941 386414 306439 386416
rect 85941 386411 86007 386414
rect 306373 386411 306439 386414
rect 68829 385794 68895 385797
rect 68829 385792 70226 385794
rect 68829 385736 68834 385792
rect 68890 385736 70226 385792
rect 68829 385734 70226 385736
rect 68829 385731 68895 385734
rect 70166 385250 70226 385734
rect 134609 385658 134675 385661
rect 251214 385658 251220 385660
rect 134609 385656 251220 385658
rect 134609 385600 134614 385656
rect 134670 385600 251220 385656
rect 134609 385598 251220 385600
rect 134609 385595 134675 385598
rect 251214 385596 251220 385598
rect 251284 385596 251290 385660
rect 112294 385324 112300 385388
rect 112364 385386 112370 385388
rect 117313 385386 117379 385389
rect 112364 385384 117379 385386
rect 112364 385328 117318 385384
rect 117374 385328 117379 385384
rect 112364 385326 117379 385328
rect 112364 385324 112370 385326
rect 117313 385323 117379 385326
rect 122097 385250 122163 385253
rect 70166 385248 122163 385250
rect 70166 385192 122102 385248
rect 122158 385192 122163 385248
rect 70166 385190 122163 385192
rect 122097 385187 122163 385190
rect 117497 384978 117563 384981
rect 118233 384978 118299 384981
rect 115828 384976 118299 384978
rect 66110 384780 66116 384844
rect 66180 384842 66186 384844
rect 70166 384842 70226 384948
rect 115828 384920 117502 384976
rect 117558 384920 118238 384976
rect 118294 384920 118299 384976
rect 115828 384918 118299 384920
rect 117497 384915 117563 384918
rect 118233 384915 118299 384918
rect 66180 384782 70226 384842
rect 66180 384780 66186 384782
rect -960 384284 480 384524
rect 115422 384508 115428 384572
rect 115492 384570 115498 384572
rect 300853 384570 300919 384573
rect 115492 384568 300919 384570
rect 115492 384512 300858 384568
rect 300914 384512 300919 384568
rect 115492 384510 300919 384512
rect 115492 384508 115498 384510
rect 300853 384507 300919 384510
rect 116117 384298 116183 384301
rect 116669 384298 116735 384301
rect 115828 384296 116735 384298
rect 115828 384240 116122 384296
rect 116178 384240 116674 384296
rect 116730 384240 116735 384296
rect 115828 384238 116735 384240
rect 116117 384235 116183 384238
rect 116669 384235 116735 384238
rect 116117 383618 116183 383621
rect 116761 383618 116827 383621
rect 115828 383616 116827 383618
rect 68737 383482 68803 383485
rect 70166 383482 70226 383588
rect 115828 383560 116122 383616
rect 116178 383560 116766 383616
rect 116822 383560 116827 383616
rect 115828 383558 116827 383560
rect 116117 383555 116183 383558
rect 116761 383555 116827 383558
rect 68737 383480 70226 383482
rect 68737 383424 68742 383480
rect 68798 383424 70226 383480
rect 68737 383422 70226 383424
rect 68737 383419 68803 383422
rect 42609 383210 42675 383213
rect 69974 383210 69980 383212
rect 42609 383208 69980 383210
rect 42609 383152 42614 383208
rect 42670 383152 69980 383208
rect 42609 383150 69980 383152
rect 42609 383147 42675 383150
rect 69974 383148 69980 383150
rect 70044 383148 70050 383212
rect 67725 382530 67791 382533
rect 70166 382530 70226 382908
rect 67725 382528 70226 382530
rect 67725 382472 67730 382528
rect 67786 382472 70226 382528
rect 67725 382470 70226 382472
rect 67725 382467 67791 382470
rect 117313 382258 117379 382261
rect 115828 382256 117379 382258
rect 67633 382122 67699 382125
rect 70166 382122 70226 382228
rect 115828 382200 117318 382256
rect 117374 382200 117379 382256
rect 115828 382198 117379 382200
rect 117313 382195 117379 382198
rect 67633 382120 70226 382122
rect 67633 382064 67638 382120
rect 67694 382064 70226 382120
rect 67633 382062 70226 382064
rect 67633 382059 67699 382062
rect 118918 381578 118924 381580
rect 115828 381518 118924 381578
rect 118918 381516 118924 381518
rect 118988 381516 118994 381580
rect 118918 380972 118924 381036
rect 118988 381034 118994 381036
rect 120257 381034 120323 381037
rect 118988 381032 120323 381034
rect 118988 380976 120262 381032
rect 120318 380976 120323 381032
rect 118988 380974 120323 380976
rect 118988 380972 118994 380974
rect 120257 380971 120323 380974
rect 117313 380898 117379 380901
rect 115828 380896 117379 380898
rect 67633 380762 67699 380765
rect 70166 380762 70226 380868
rect 115828 380840 117318 380896
rect 117374 380840 117379 380896
rect 115828 380838 117379 380840
rect 117313 380835 117379 380838
rect 67633 380760 70226 380762
rect 67633 380704 67638 380760
rect 67694 380704 70226 380760
rect 67633 380702 70226 380704
rect 67633 380699 67699 380702
rect 68001 380354 68067 380357
rect 69054 380354 69060 380356
rect 68001 380352 69060 380354
rect 68001 380296 68006 380352
rect 68062 380296 69060 380352
rect 68001 380294 69060 380296
rect 68001 380291 68067 380294
rect 69054 380292 69060 380294
rect 69124 380354 69130 380356
rect 69124 380294 70226 380354
rect 69124 380292 69130 380294
rect 70166 380188 70226 380294
rect 67449 379946 67515 379949
rect 67449 379944 70226 379946
rect 67449 379888 67454 379944
rect 67510 379888 70226 379944
rect 67449 379886 70226 379888
rect 67449 379883 67515 379886
rect 70166 379508 70226 379886
rect 117681 379538 117747 379541
rect 115828 379536 117747 379538
rect 115828 379480 117686 379536
rect 117742 379480 117747 379536
rect 115828 379478 117747 379480
rect 117681 379475 117747 379478
rect 118601 378858 118667 378861
rect 115828 378856 118667 378858
rect 115828 378800 118606 378856
rect 118662 378800 118667 378856
rect 115828 378798 118667 378800
rect 118601 378795 118667 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 67633 378314 67699 378317
rect 67633 378312 70226 378314
rect 67633 378256 67638 378312
rect 67694 378256 70226 378312
rect 583520 378300 584960 378390
rect 67633 378254 70226 378256
rect 67633 378251 67699 378254
rect 70166 378148 70226 378254
rect 118785 378178 118851 378181
rect 115828 378176 118851 378178
rect 115828 378120 118790 378176
rect 118846 378120 118851 378176
rect 115828 378118 118851 378120
rect 118785 378115 118851 378118
rect 52310 377708 52316 377772
rect 52380 377770 52386 377772
rect 70526 377770 70532 377772
rect 52380 377710 70532 377770
rect 52380 377708 52386 377710
rect 70526 377708 70532 377710
rect 70596 377708 70602 377772
rect 62982 377300 62988 377364
rect 63052 377362 63058 377364
rect 67633 377362 67699 377365
rect 70166 377362 70226 377468
rect 63052 377302 64890 377362
rect 63052 377300 63058 377302
rect 64830 377226 64890 377302
rect 67633 377360 70226 377362
rect 67633 377304 67638 377360
rect 67694 377304 70226 377360
rect 67633 377302 70226 377304
rect 119337 377362 119403 377365
rect 252502 377362 252508 377364
rect 119337 377360 252508 377362
rect 119337 377304 119342 377360
rect 119398 377304 252508 377360
rect 119337 377302 252508 377304
rect 67633 377299 67699 377302
rect 119337 377299 119403 377302
rect 252502 377300 252508 377302
rect 252572 377300 252578 377364
rect 68870 377226 68876 377228
rect 64830 377166 68876 377226
rect 68870 377164 68876 377166
rect 68940 377226 68946 377228
rect 68940 377166 70226 377226
rect 68940 377164 68946 377166
rect 70166 376788 70226 377166
rect 118601 376818 118667 376821
rect 115828 376816 118667 376818
rect 115828 376760 118606 376816
rect 118662 376760 118667 376816
rect 115828 376758 118667 376760
rect 118601 376755 118667 376758
rect 118601 376138 118667 376141
rect 115828 376136 118667 376138
rect 115828 376080 118606 376136
rect 118662 376080 118667 376136
rect 115828 376078 118667 376080
rect 118601 376075 118667 376078
rect 30281 376002 30347 376005
rect 65374 376002 65380 376004
rect 30281 376000 65380 376002
rect 30281 375944 30286 376000
rect 30342 375944 65380 376000
rect 30281 375942 65380 375944
rect 30281 375939 30347 375942
rect 65374 375940 65380 375942
rect 65444 376002 65450 376004
rect 122281 376002 122347 376005
rect 255262 376002 255268 376004
rect 65444 375942 70226 376002
rect 65444 375940 65450 375942
rect 70166 375428 70226 375942
rect 122281 376000 255268 376002
rect 122281 375944 122286 376000
rect 122342 375944 255268 376000
rect 122281 375942 255268 375944
rect 122281 375939 122347 375942
rect 255262 375940 255268 375942
rect 255332 375940 255338 376004
rect 118509 375458 118575 375461
rect 115828 375456 118575 375458
rect 115828 375400 118514 375456
rect 118570 375400 118575 375456
rect 115828 375398 118575 375400
rect 118509 375395 118575 375398
rect 67633 375186 67699 375189
rect 67633 375184 70226 375186
rect 67633 375128 67638 375184
rect 67694 375128 70226 375184
rect 67633 375126 70226 375128
rect 67633 375123 67699 375126
rect 70166 374748 70226 375126
rect 67725 374234 67791 374237
rect 67725 374232 70226 374234
rect 67725 374176 67730 374232
rect 67786 374176 70226 374232
rect 67725 374174 70226 374176
rect 67725 374171 67791 374174
rect 70166 374068 70226 374174
rect 118601 374098 118667 374101
rect 115828 374096 118667 374098
rect 115828 374040 118606 374096
rect 118662 374040 118667 374096
rect 115828 374038 118667 374040
rect 118601 374035 118667 374038
rect 117497 373418 117563 373421
rect 115828 373416 117563 373418
rect 115828 373360 117502 373416
rect 117558 373360 117563 373416
rect 115828 373358 117563 373360
rect 117497 373355 117563 373358
rect 68921 372876 68987 372877
rect 68870 372874 68876 372876
rect 68794 372814 68876 372874
rect 68940 372874 68987 372876
rect 68940 372872 70226 372874
rect 68982 372816 70226 372872
rect 68870 372812 68876 372814
rect 68940 372814 70226 372816
rect 68940 372812 68987 372814
rect 68921 372811 68987 372812
rect 70166 372708 70226 372814
rect 117078 372738 117084 372740
rect 115828 372678 117084 372738
rect 117078 372676 117084 372678
rect 117148 372738 117154 372740
rect 118417 372738 118483 372741
rect 117148 372736 118483 372738
rect 117148 372680 118422 372736
rect 118478 372680 118483 372736
rect 117148 372678 118483 372680
rect 117148 372676 117154 372678
rect 118417 372675 118483 372678
rect 67633 372466 67699 372469
rect 67633 372464 70226 372466
rect 67633 372408 67638 372464
rect 67694 372408 70226 372464
rect 67633 372406 70226 372408
rect 67633 372403 67699 372406
rect 70166 372028 70226 372406
rect 67633 371514 67699 371517
rect 67633 371512 70226 371514
rect -960 371378 480 371468
rect 67633 371456 67638 371512
rect 67694 371456 70226 371512
rect 67633 371454 70226 371456
rect 67633 371451 67699 371454
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect 70166 371348 70226 371454
rect 117998 371378 118004 371380
rect -960 371318 3299 371320
rect 115828 371318 118004 371378
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 117998 371316 118004 371318
rect 118068 371378 118074 371380
rect 118601 371378 118667 371381
rect 118068 371376 118667 371378
rect 118068 371320 118606 371376
rect 118662 371320 118667 371376
rect 118068 371318 118667 371320
rect 118068 371316 118074 371318
rect 118601 371315 118667 371318
rect 48037 370562 48103 370565
rect 55070 370562 55076 370564
rect 48037 370560 55076 370562
rect 48037 370504 48042 370560
rect 48098 370504 55076 370560
rect 48037 370502 55076 370504
rect 48037 370499 48103 370502
rect 55070 370500 55076 370502
rect 55140 370562 55146 370564
rect 55140 370502 70226 370562
rect 55140 370500 55146 370502
rect 70166 369988 70226 370502
rect 115798 370290 115858 370668
rect 122230 370500 122236 370564
rect 122300 370562 122306 370564
rect 304942 370562 304948 370564
rect 122300 370502 304948 370562
rect 122300 370500 122306 370502
rect 304942 370500 304948 370502
rect 305012 370500 305018 370564
rect 116025 370290 116091 370293
rect 115798 370288 116091 370290
rect 115798 370232 116030 370288
rect 116086 370232 116091 370288
rect 115798 370230 116091 370232
rect 116025 370227 116091 370230
rect 118877 370018 118943 370021
rect 115828 370016 118943 370018
rect 115828 369960 118882 370016
rect 118938 369960 118943 370016
rect 115828 369958 118943 369960
rect 118877 369955 118943 369958
rect 67725 369202 67791 369205
rect 70166 369202 70226 369308
rect 67725 369200 70226 369202
rect 67725 369144 67730 369200
rect 67786 369144 70226 369200
rect 67725 369142 70226 369144
rect 67725 369139 67791 369142
rect 67633 369066 67699 369069
rect 123845 369066 123911 369069
rect 299606 369066 299612 369068
rect 67633 369064 70226 369066
rect 67633 369008 67638 369064
rect 67694 369008 70226 369064
rect 67633 369006 70226 369008
rect 67633 369003 67699 369006
rect 70166 368628 70226 369006
rect 123845 369064 299612 369066
rect 123845 369008 123850 369064
rect 123906 369008 299612 369064
rect 123845 369006 299612 369008
rect 123845 369003 123911 369006
rect 299606 369004 299612 369006
rect 299676 369004 299682 369068
rect 118734 368658 118740 368660
rect 115828 368598 118740 368658
rect 118734 368596 118740 368598
rect 118804 368658 118810 368660
rect 118969 368658 119035 368661
rect 118804 368656 119035 368658
rect 118804 368600 118974 368656
rect 119030 368600 119035 368656
rect 118804 368598 119035 368600
rect 118804 368596 118810 368598
rect 118969 368595 119035 368598
rect 118509 367978 118575 367981
rect 115828 367976 118575 367978
rect 115828 367920 118514 367976
rect 118570 367920 118575 367976
rect 115828 367918 118575 367920
rect 118509 367915 118575 367918
rect 122097 367706 122163 367709
rect 259494 367706 259500 367708
rect 122097 367704 259500 367706
rect 122097 367648 122102 367704
rect 122158 367648 259500 367704
rect 122097 367646 259500 367648
rect 122097 367643 122163 367646
rect 259494 367644 259500 367646
rect 259564 367644 259570 367708
rect 118601 367298 118667 367301
rect 115828 367296 118667 367298
rect 67633 367162 67699 367165
rect 70166 367162 70226 367268
rect 115828 367240 118606 367296
rect 118662 367240 118667 367296
rect 115828 367238 118667 367240
rect 118601 367235 118667 367238
rect 67633 367160 70226 367162
rect 67633 367104 67638 367160
rect 67694 367104 70226 367160
rect 67633 367102 70226 367104
rect 67633 367099 67699 367102
rect 67633 366482 67699 366485
rect 70166 366482 70226 366588
rect 67633 366480 70226 366482
rect 67633 366424 67638 366480
rect 67694 366424 70226 366480
rect 67633 366422 70226 366424
rect 67633 366419 67699 366422
rect 67725 366346 67791 366349
rect 67725 366344 70226 366346
rect 67725 366288 67730 366344
rect 67786 366288 70226 366344
rect 67725 366286 70226 366288
rect 67725 366283 67791 366286
rect 70166 365908 70226 366286
rect 120758 366284 120764 366348
rect 120828 366346 120834 366348
rect 316033 366346 316099 366349
rect 120828 366344 316099 366346
rect 120828 366288 316038 366344
rect 316094 366288 316099 366344
rect 120828 366286 316099 366288
rect 120828 366284 120834 366286
rect 316033 366283 316099 366286
rect 118601 365938 118667 365941
rect 115828 365936 118667 365938
rect 115828 365880 118606 365936
rect 118662 365880 118667 365936
rect 115828 365878 118667 365880
rect 118601 365875 118667 365878
rect 118601 365258 118667 365261
rect 115828 365256 118667 365258
rect 115828 365200 118606 365256
rect 118662 365200 118667 365256
rect 115828 365198 118667 365200
rect 118601 365195 118667 365198
rect 68369 365122 68435 365125
rect 580349 365122 580415 365125
rect 583520 365122 584960 365212
rect 68369 365120 70226 365122
rect 68369 365064 68374 365120
rect 68430 365064 70226 365120
rect 68369 365062 70226 365064
rect 68369 365059 68435 365062
rect 70166 364548 70226 365062
rect 580349 365120 584960 365122
rect 580349 365064 580354 365120
rect 580410 365064 584960 365120
rect 580349 365062 584960 365064
rect 580349 365059 580415 365062
rect 583520 364972 584960 365062
rect 118601 364578 118667 364581
rect 115828 364576 118667 364578
rect 115828 364520 118606 364576
rect 118662 364520 118667 364576
rect 115828 364518 118667 364520
rect 118601 364515 118667 364518
rect 67633 363762 67699 363765
rect 70166 363762 70226 363868
rect 67633 363760 70226 363762
rect 67633 363704 67638 363760
rect 67694 363704 70226 363760
rect 67633 363702 70226 363704
rect 67633 363699 67699 363702
rect 67725 363626 67791 363629
rect 117589 363626 117655 363629
rect 302734 363626 302740 363628
rect 67725 363624 70226 363626
rect 67725 363568 67730 363624
rect 67786 363568 70226 363624
rect 67725 363566 70226 363568
rect 67725 363563 67791 363566
rect 70166 363188 70226 363566
rect 115798 363624 302740 363626
rect 115798 363568 117594 363624
rect 117650 363568 302740 363624
rect 115798 363566 302740 363568
rect 115798 363188 115858 363566
rect 117589 363563 117655 363566
rect 302734 363564 302740 363566
rect 302804 363564 302810 363628
rect 117957 362538 118023 362541
rect 115828 362536 118023 362538
rect 67633 362130 67699 362133
rect 70166 362130 70226 362508
rect 115828 362480 117962 362536
rect 118018 362480 118023 362536
rect 115828 362478 118023 362480
rect 117957 362475 118023 362478
rect 153101 362266 153167 362269
rect 242014 362266 242020 362268
rect 153101 362264 242020 362266
rect 153101 362208 153106 362264
rect 153162 362208 242020 362264
rect 153101 362206 242020 362208
rect 153101 362203 153167 362206
rect 242014 362204 242020 362206
rect 242084 362204 242090 362268
rect 67633 362128 70226 362130
rect 67633 362072 67638 362128
rect 67694 362072 70226 362128
rect 67633 362070 70226 362072
rect 67633 362067 67699 362070
rect 118601 361858 118667 361861
rect 115828 361856 118667 361858
rect 115828 361800 118606 361856
rect 118662 361800 118667 361856
rect 115828 361798 118667 361800
rect 118601 361795 118667 361798
rect 118601 361178 118667 361181
rect 115828 361176 118667 361178
rect 67633 361042 67699 361045
rect 70166 361042 70226 361148
rect 115828 361120 118606 361176
rect 118662 361120 118667 361176
rect 115828 361118 118667 361120
rect 118601 361115 118667 361118
rect 67633 361040 70226 361042
rect 67633 360984 67638 361040
rect 67694 360984 70226 361040
rect 67633 360982 70226 360984
rect 67633 360979 67699 360982
rect 69197 360906 69263 360909
rect 69197 360904 70226 360906
rect 69197 360848 69202 360904
rect 69258 360848 70226 360904
rect 69197 360846 70226 360848
rect 69197 360843 69263 360846
rect 70166 360468 70226 360846
rect 123334 360844 123340 360908
rect 123404 360906 123410 360908
rect 318793 360906 318859 360909
rect 123404 360904 318859 360906
rect 123404 360848 318798 360904
rect 318854 360848 318859 360904
rect 123404 360846 318859 360848
rect 123404 360844 123410 360846
rect 318793 360843 318859 360846
rect 116669 359818 116735 359821
rect 115828 359816 116735 359818
rect 67633 359546 67699 359549
rect 70166 359546 70226 359788
rect 115828 359760 116674 359816
rect 116730 359760 116735 359816
rect 115828 359758 116735 359760
rect 116669 359755 116735 359758
rect 67633 359544 70226 359546
rect 67633 359488 67638 359544
rect 67694 359488 70226 359544
rect 67633 359486 70226 359488
rect 67633 359483 67699 359486
rect 118141 359138 118207 359141
rect 115828 359136 118207 359138
rect 115828 359080 118146 359136
rect 118202 359080 118207 359136
rect 115828 359078 118207 359080
rect 118141 359075 118207 359078
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 118601 358458 118667 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect 115828 358456 118667 358458
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 67725 358186 67791 358189
rect 70166 358186 70226 358428
rect 115828 358400 118606 358456
rect 118662 358400 118667 358456
rect 115828 358398 118667 358400
rect 118601 358395 118667 358398
rect 67725 358184 70226 358186
rect 67725 358128 67730 358184
rect 67786 358128 70226 358184
rect 67725 358126 70226 358128
rect 67725 358123 67791 358126
rect 67633 358050 67699 358053
rect 67633 358048 70226 358050
rect 67633 357992 67638 358048
rect 67694 357992 70226 358048
rect 67633 357990 70226 357992
rect 67633 357987 67699 357990
rect 70166 357748 70226 357990
rect 115974 357370 115980 357372
rect 115798 357310 115980 357370
rect 115798 357098 115858 357310
rect 115974 357308 115980 357310
rect 116044 357308 116050 357372
rect 117681 357098 117747 357101
rect 115798 357096 117747 357098
rect 115798 357068 117686 357096
rect 69105 356962 69171 356965
rect 69473 356962 69539 356965
rect 70166 356962 70226 357068
rect 115828 357040 117686 357068
rect 117742 357040 117747 357096
rect 115828 357038 117747 357040
rect 117681 357035 117747 357038
rect 69105 356960 70226 356962
rect 69105 356904 69110 356960
rect 69166 356904 69478 356960
rect 69534 356904 70226 356960
rect 69105 356902 70226 356904
rect 69105 356899 69171 356902
rect 69473 356899 69539 356902
rect 115798 356146 115858 356388
rect 119981 356146 120047 356149
rect 124806 356146 124812 356148
rect 115798 356144 124812 356146
rect 115798 356088 119986 356144
rect 120042 356088 124812 356144
rect 115798 356086 124812 356088
rect 119981 356083 120047 356086
rect 124806 356084 124812 356086
rect 124876 356084 124882 356148
rect 118601 355738 118667 355741
rect 115828 355736 118667 355738
rect 67633 355602 67699 355605
rect 70166 355602 70226 355708
rect 115828 355680 118606 355736
rect 118662 355680 118667 355736
rect 115828 355678 118667 355680
rect 118601 355675 118667 355678
rect 67633 355600 70226 355602
rect 67633 355544 67638 355600
rect 67694 355544 70226 355600
rect 67633 355542 70226 355544
rect 67633 355539 67699 355542
rect 67725 355466 67791 355469
rect 67725 355464 70226 355466
rect 67725 355408 67730 355464
rect 67786 355408 70226 355464
rect 67725 355406 70226 355408
rect 67725 355403 67791 355406
rect 49601 355330 49667 355333
rect 61694 355330 61700 355332
rect 49601 355328 61700 355330
rect 49601 355272 49606 355328
rect 49662 355272 61700 355328
rect 49601 355270 61700 355272
rect 49601 355267 49667 355270
rect 61694 355268 61700 355270
rect 61764 355330 61770 355332
rect 63493 355330 63559 355333
rect 61764 355328 63559 355330
rect 61764 355272 63498 355328
rect 63554 355272 63559 355328
rect 61764 355270 63559 355272
rect 61764 355268 61770 355270
rect 63493 355267 63559 355270
rect 70166 355028 70226 355406
rect 118049 354378 118115 354381
rect 115828 354376 118115 354378
rect 67633 353834 67699 353837
rect 70166 353834 70226 354348
rect 115828 354320 118054 354376
rect 118110 354320 118115 354376
rect 115828 354318 118115 354320
rect 118049 354315 118115 354318
rect 67633 353832 70226 353834
rect 67633 353776 67638 353832
rect 67694 353776 70226 353832
rect 67633 353774 70226 353776
rect 67633 353771 67699 353774
rect 118601 353698 118667 353701
rect 115828 353696 118667 353698
rect 115828 353640 118606 353696
rect 118662 353640 118667 353696
rect 115828 353638 118667 353640
rect 118601 353635 118667 353638
rect 115933 353290 115999 353293
rect 115798 353288 115999 353290
rect 115798 353232 115938 353288
rect 115994 353232 115999 353288
rect 115798 353230 115999 353232
rect 115798 353018 115858 353230
rect 115933 353227 115999 353230
rect 117957 353018 118023 353021
rect 115798 353016 118023 353018
rect 115798 352988 117962 353016
rect 67633 352610 67699 352613
rect 70166 352610 70226 352988
rect 115828 352960 117962 352988
rect 118018 352960 118023 353016
rect 115828 352958 118023 352960
rect 117957 352955 118023 352958
rect 67633 352608 70226 352610
rect 67633 352552 67638 352608
rect 67694 352552 70226 352608
rect 67633 352550 70226 352552
rect 67633 352547 67699 352550
rect 67909 352474 67975 352477
rect 68737 352474 68803 352477
rect 67909 352472 70226 352474
rect 67909 352416 67914 352472
rect 67970 352416 68742 352472
rect 68798 352416 70226 352472
rect 67909 352414 70226 352416
rect 67909 352411 67975 352414
rect 68737 352411 68803 352414
rect 70166 352308 70226 352414
rect 580257 351930 580323 351933
rect 583520 351930 584960 352020
rect 580257 351928 584960 351930
rect 580257 351872 580262 351928
rect 580318 351872 584960 351928
rect 580257 351870 584960 351872
rect 580257 351867 580323 351870
rect 583520 351780 584960 351870
rect 117405 351658 117471 351661
rect 118509 351658 118575 351661
rect 115828 351656 118575 351658
rect 67725 351522 67791 351525
rect 68277 351522 68343 351525
rect 70166 351522 70226 351628
rect 115828 351600 117410 351656
rect 117466 351600 118514 351656
rect 118570 351600 118575 351656
rect 115828 351598 118575 351600
rect 117405 351595 117471 351598
rect 118509 351595 118575 351598
rect 67725 351520 70226 351522
rect 67725 351464 67730 351520
rect 67786 351464 68282 351520
rect 68338 351464 70226 351520
rect 67725 351462 70226 351464
rect 67725 351459 67791 351462
rect 68277 351459 68343 351462
rect 117313 350978 117379 350981
rect 118417 350978 118483 350981
rect 115828 350976 118483 350978
rect 115828 350920 117318 350976
rect 117374 350920 118422 350976
rect 118478 350920 118483 350976
rect 115828 350918 118483 350920
rect 117313 350915 117379 350918
rect 118417 350915 118483 350918
rect 118601 350298 118667 350301
rect 115828 350296 118667 350298
rect 67633 349890 67699 349893
rect 70166 349890 70226 350268
rect 115828 350240 118606 350296
rect 118662 350240 118667 350296
rect 115828 350238 118667 350240
rect 118601 350235 118667 350238
rect 67633 349888 70226 349890
rect 67633 349832 67638 349888
rect 67694 349832 70226 349888
rect 67633 349830 70226 349832
rect 67633 349827 67699 349830
rect 68001 349754 68067 349757
rect 68921 349754 68987 349757
rect 68001 349752 70226 349754
rect 68001 349696 68006 349752
rect 68062 349696 68926 349752
rect 68982 349696 70226 349752
rect 68001 349694 70226 349696
rect 68001 349691 68067 349694
rect 68921 349691 68987 349694
rect 70166 349588 70226 349694
rect 115289 349210 115355 349213
rect 115289 349208 115490 349210
rect 115289 349152 115294 349208
rect 115350 349152 115490 349208
rect 115289 349150 115490 349152
rect 115289 349147 115355 349150
rect 115430 349074 115490 349150
rect 115430 349014 115858 349074
rect 115798 348938 115858 349014
rect 117773 348938 117839 348941
rect 115798 348936 117839 348938
rect 115798 348908 117778 348936
rect 68829 348394 68895 348397
rect 70166 348394 70226 348908
rect 115828 348880 117778 348908
rect 117834 348880 117839 348936
rect 115828 348878 117839 348880
rect 117773 348875 117839 348878
rect 68829 348392 70226 348394
rect 68829 348336 68834 348392
rect 68890 348336 70226 348392
rect 68829 348334 70226 348336
rect 68829 348331 68895 348334
rect 118601 348258 118667 348261
rect 115828 348256 118667 348258
rect 115828 348200 118606 348256
rect 118662 348200 118667 348256
rect 115828 348198 118667 348200
rect 118601 348195 118667 348198
rect 117405 347578 117471 347581
rect 115828 347576 117471 347578
rect 68553 347170 68619 347173
rect 70166 347170 70226 347548
rect 115828 347520 117410 347576
rect 117466 347520 117471 347576
rect 115828 347518 117471 347520
rect 117405 347515 117471 347518
rect 68553 347168 70226 347170
rect 68553 347112 68558 347168
rect 68614 347112 70226 347168
rect 68553 347110 70226 347112
rect 68553 347107 68619 347110
rect 67633 346762 67699 346765
rect 70166 346762 70226 346868
rect 67633 346760 70226 346762
rect 67633 346704 67638 346760
rect 67694 346704 70226 346760
rect 67633 346702 70226 346704
rect 67633 346699 67699 346702
rect 118325 346218 118391 346221
rect 115828 346216 118391 346218
rect 67725 345674 67791 345677
rect 70166 345674 70226 346188
rect 115828 346160 118330 346216
rect 118386 346160 118391 346216
rect 115828 346158 118391 346160
rect 118325 346155 118391 346158
rect 67725 345672 70226 345674
rect 67725 345616 67730 345672
rect 67786 345616 70226 345672
rect 67725 345614 70226 345616
rect 67725 345611 67791 345614
rect 118601 345538 118667 345541
rect 115828 345536 118667 345538
rect -960 345402 480 345492
rect 115828 345480 118606 345536
rect 118662 345480 118667 345536
rect 115828 345478 118667 345480
rect 118601 345475 118667 345478
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 118601 344858 118667 344861
rect 115828 344856 118667 344858
rect 67725 344450 67791 344453
rect 70166 344450 70226 344828
rect 115828 344800 118606 344856
rect 118662 344800 118667 344856
rect 115828 344798 118667 344800
rect 118601 344795 118667 344798
rect 67725 344448 70226 344450
rect 67725 344392 67730 344448
rect 67786 344392 70226 344448
rect 67725 344390 70226 344392
rect 67725 344387 67791 344390
rect 67633 343770 67699 343773
rect 70166 343770 70226 344148
rect 67633 343768 70226 343770
rect 67633 343712 67638 343768
rect 67694 343712 70226 343768
rect 67633 343710 70226 343712
rect 67633 343707 67699 343710
rect 118141 343498 118207 343501
rect 115828 343496 118207 343498
rect 70350 342956 70410 343468
rect 115828 343440 118146 343496
rect 118202 343440 118207 343496
rect 115828 343438 118207 343440
rect 118141 343435 118207 343438
rect 70342 342892 70348 342956
rect 70412 342892 70418 342956
rect 70350 342818 70410 342892
rect 118601 342818 118667 342821
rect 64830 342758 70410 342818
rect 115828 342816 118667 342818
rect 115828 342760 118606 342816
rect 118662 342760 118667 342816
rect 115828 342758 118667 342760
rect 61878 342212 61884 342276
rect 61948 342274 61954 342276
rect 64830 342274 64890 342758
rect 118601 342755 118667 342758
rect 61948 342214 64890 342274
rect 61948 342212 61954 342214
rect 118601 342138 118667 342141
rect 115828 342136 118667 342138
rect 67633 341730 67699 341733
rect 70166 341730 70226 342108
rect 115828 342080 118606 342136
rect 118662 342080 118667 342136
rect 115828 342078 118667 342080
rect 118601 342075 118667 342078
rect 67633 341728 70226 341730
rect 67633 341672 67638 341728
rect 67694 341672 70226 341728
rect 67633 341670 70226 341672
rect 67633 341667 67699 341670
rect 67541 341594 67607 341597
rect 67541 341592 70594 341594
rect 67541 341536 67546 341592
rect 67602 341536 70594 341592
rect 67541 341534 70594 341536
rect 67541 341531 67607 341534
rect 70534 341052 70594 341534
rect 124806 341396 124812 341460
rect 124876 341458 124882 341460
rect 140865 341458 140931 341461
rect 124876 341456 140931 341458
rect 124876 341400 140870 341456
rect 140926 341400 140931 341456
rect 124876 341398 140931 341400
rect 124876 341396 124882 341398
rect 140865 341395 140931 341398
rect 70526 340988 70532 341052
rect 70596 340988 70602 341052
rect 48037 340780 48103 340781
rect 48037 340776 48084 340780
rect 48148 340778 48154 340780
rect 48037 340720 48042 340776
rect 48037 340716 48084 340720
rect 48148 340718 48194 340778
rect 48148 340716 48154 340718
rect 64638 340716 64644 340780
rect 64708 340778 64714 340780
rect 118049 340778 118115 340781
rect 64708 340718 64890 340778
rect 115828 340776 118115 340778
rect 64708 340716 64714 340718
rect 48037 340715 48103 340716
rect 64830 340642 64890 340718
rect 70534 340642 70594 340748
rect 115828 340720 118054 340776
rect 118110 340720 118115 340776
rect 115828 340718 118115 340720
rect 118049 340715 118115 340718
rect 64830 340582 70594 340642
rect 70534 339962 70594 340582
rect 117773 340098 117839 340101
rect 115828 340096 117839 340098
rect 115828 340068 117778 340096
rect 115798 340040 117778 340068
rect 117834 340040 117839 340096
rect 115798 340038 117839 340040
rect 71129 339962 71195 339965
rect 70534 339960 71195 339962
rect 70534 339904 71134 339960
rect 71190 339904 71195 339960
rect 70534 339902 71195 339904
rect 71129 339899 71195 339902
rect 52310 339628 52316 339692
rect 52380 339690 52386 339692
rect 79041 339690 79107 339693
rect 52380 339688 79107 339690
rect 52380 339632 79046 339688
rect 79102 339632 79107 339688
rect 52380 339630 79107 339632
rect 52380 339628 52386 339630
rect 79041 339627 79107 339630
rect 115381 339554 115447 339557
rect 115798 339554 115858 340038
rect 117773 340035 117839 340038
rect 115381 339552 115858 339554
rect 115381 339496 115386 339552
rect 115442 339496 115858 339552
rect 115381 339494 115858 339496
rect 115381 339491 115447 339494
rect 44030 339356 44036 339420
rect 44100 339418 44106 339420
rect 75821 339418 75887 339421
rect 44100 339416 75887 339418
rect 44100 339360 75826 339416
rect 75882 339360 75887 339416
rect 44100 339358 75887 339360
rect 44100 339356 44106 339358
rect 75821 339355 75887 339358
rect 583520 338452 584960 338692
rect 38469 338058 38535 338061
rect 71313 338058 71379 338061
rect 38469 338056 71379 338058
rect 38469 338000 38474 338056
rect 38530 338000 71318 338056
rect 71374 338000 71379 338056
rect 38469 337998 71379 338000
rect 38469 337995 38535 337998
rect 71313 337995 71379 337998
rect 128445 338058 128511 338061
rect 128670 338058 128676 338060
rect 128445 338056 128676 338058
rect 128445 338000 128450 338056
rect 128506 338000 128676 338056
rect 128445 337998 128676 338000
rect 128445 337995 128511 337998
rect 128670 337996 128676 337998
rect 128740 337996 128746 338060
rect 61377 337924 61443 337925
rect 57830 337860 57836 337924
rect 57900 337922 57906 337924
rect 61326 337922 61332 337924
rect 57900 337862 61332 337922
rect 61396 337922 61443 337924
rect 61396 337920 61524 337922
rect 61438 337864 61524 337920
rect 57900 337860 57906 337862
rect 61326 337860 61332 337862
rect 61396 337862 61524 337864
rect 61396 337860 61443 337862
rect 61377 337859 61443 337860
rect 71313 337514 71379 337517
rect 84837 337514 84903 337517
rect 71313 337512 84903 337514
rect 71313 337456 71318 337512
rect 71374 337456 84842 337512
rect 84898 337456 84903 337512
rect 71313 337454 84903 337456
rect 71313 337451 71379 337454
rect 84837 337451 84903 337454
rect 120441 337514 120507 337517
rect 126094 337514 126100 337516
rect 120441 337512 126100 337514
rect 120441 337456 120446 337512
rect 120502 337456 126100 337512
rect 120441 337454 126100 337456
rect 120441 337451 120507 337454
rect 126094 337452 126100 337454
rect 126164 337452 126170 337516
rect 79041 337378 79107 337381
rect 124806 337378 124812 337380
rect 79041 337376 124812 337378
rect 79041 337320 79046 337376
rect 79102 337320 124812 337376
rect 79041 337318 124812 337320
rect 79041 337315 79107 337318
rect 124806 337316 124812 337318
rect 124876 337316 124882 337380
rect 70526 336092 70532 336156
rect 70596 336154 70602 336156
rect 292614 336154 292620 336156
rect 70596 336094 292620 336154
rect 70596 336092 70602 336094
rect 292614 336092 292620 336094
rect 292684 336092 292690 336156
rect 70342 335956 70348 336020
rect 70412 336018 70418 336020
rect 328453 336018 328519 336021
rect 70412 336016 328519 336018
rect 70412 335960 328458 336016
rect 328514 335960 328519 336016
rect 70412 335958 328519 335960
rect 70412 335956 70418 335958
rect 328453 335955 328519 335958
rect 68645 334794 68711 334797
rect 248454 334794 248460 334796
rect 68645 334792 248460 334794
rect 68645 334736 68650 334792
rect 68706 334736 248460 334792
rect 68645 334734 248460 334736
rect 68645 334731 68711 334734
rect 248454 334732 248460 334734
rect 248524 334732 248530 334796
rect 72969 334658 73035 334661
rect 291142 334658 291148 334660
rect 72969 334656 291148 334658
rect 72969 334600 72974 334656
rect 73030 334600 291148 334656
rect 72969 334598 291148 334600
rect 72969 334595 73035 334598
rect 291142 334596 291148 334598
rect 291212 334596 291218 334660
rect 53598 333916 53604 333980
rect 53668 333978 53674 333980
rect 89069 333978 89135 333981
rect 53668 333976 89135 333978
rect 53668 333920 89074 333976
rect 89130 333920 89135 333976
rect 53668 333918 89135 333920
rect 53668 333916 53674 333918
rect 89069 333915 89135 333918
rect 68737 333298 68803 333301
rect 288382 333298 288388 333300
rect 68737 333296 288388 333298
rect 68737 333240 68742 333296
rect 68798 333240 288388 333296
rect 68737 333238 288388 333240
rect 68737 333235 68803 333238
rect 288382 333236 288388 333238
rect 288452 333236 288458 333300
rect 125777 332484 125843 332485
rect 125726 332482 125732 332484
rect -960 332196 480 332436
rect 125686 332422 125732 332482
rect 125796 332480 125843 332484
rect 125838 332424 125843 332480
rect 125726 332420 125732 332422
rect 125796 332420 125843 332424
rect 125777 332419 125843 332420
rect 78673 331802 78739 331805
rect 244222 331802 244228 331804
rect 78673 331800 244228 331802
rect 78673 331744 78678 331800
rect 78734 331744 244228 331800
rect 78673 331742 244228 331744
rect 78673 331739 78739 331742
rect 244222 331740 244228 331742
rect 244292 331740 244298 331804
rect 96521 331122 96587 331125
rect 122598 331122 122604 331124
rect 96521 331120 122604 331122
rect 96521 331064 96526 331120
rect 96582 331064 122604 331120
rect 96521 331062 122604 331064
rect 96521 331059 96587 331062
rect 122598 331060 122604 331062
rect 122668 331060 122674 331124
rect 95233 330714 95299 330717
rect 96521 330714 96587 330717
rect 95233 330712 96587 330714
rect 95233 330656 95238 330712
rect 95294 330656 96526 330712
rect 96582 330656 96587 330712
rect 95233 330654 96587 330656
rect 95233 330651 95299 330654
rect 96521 330651 96587 330654
rect 55070 330380 55076 330444
rect 55140 330442 55146 330444
rect 111057 330442 111123 330445
rect 55140 330440 111123 330442
rect 55140 330384 111062 330440
rect 111118 330384 111123 330440
rect 55140 330382 111123 330384
rect 55140 330380 55146 330382
rect 111057 330379 111123 330382
rect 133137 329764 133203 329765
rect 133086 329762 133092 329764
rect 133046 329702 133092 329762
rect 133156 329760 133203 329764
rect 133198 329704 133203 329760
rect 133086 329700 133092 329702
rect 133156 329700 133203 329704
rect 133137 329699 133203 329700
rect 133781 329082 133847 329085
rect 298686 329082 298692 329084
rect 133781 329080 298692 329082
rect 133781 329024 133786 329080
rect 133842 329024 298692 329080
rect 133781 329022 298692 329024
rect 133781 329019 133847 329022
rect 298686 329020 298692 329022
rect 298756 329020 298762 329084
rect 129825 328404 129891 328405
rect 129774 328402 129780 328404
rect 129734 328342 129780 328402
rect 129844 328400 129891 328404
rect 129886 328344 129891 328400
rect 129774 328340 129780 328342
rect 129844 328340 129891 328344
rect 129825 328339 129891 328340
rect 580349 325274 580415 325277
rect 583520 325274 584960 325364
rect 580349 325272 584960 325274
rect 580349 325216 580354 325272
rect 580410 325216 584960 325272
rect 580349 325214 584960 325216
rect 580349 325211 580415 325214
rect 583520 325124 584960 325214
rect 124305 324324 124371 324325
rect 124254 324322 124260 324324
rect 124214 324262 124260 324322
rect 124324 324320 124371 324324
rect 124366 324264 124371 324320
rect 124254 324260 124260 324262
rect 124324 324260 124371 324264
rect 124305 324259 124371 324260
rect 61694 323716 61700 323780
rect 61764 323778 61770 323780
rect 133965 323778 134031 323781
rect 61764 323776 134031 323778
rect 61764 323720 133970 323776
rect 134026 323720 134031 323776
rect 61764 323718 134031 323720
rect 61764 323716 61770 323718
rect 133965 323715 134031 323718
rect 65374 323580 65380 323644
rect 65444 323642 65450 323644
rect 327073 323642 327139 323645
rect 65444 323640 327139 323642
rect 65444 323584 327078 323640
rect 327134 323584 327139 323640
rect 65444 323582 327139 323584
rect 65444 323580 65450 323582
rect 327073 323579 327139 323582
rect 82077 322146 82143 322149
rect 245694 322146 245700 322148
rect 82077 322144 245700 322146
rect 82077 322088 82082 322144
rect 82138 322088 245700 322144
rect 82077 322086 245700 322088
rect 82077 322083 82143 322086
rect 245694 322084 245700 322086
rect 245764 322084 245770 322148
rect 66161 320786 66227 320789
rect 249742 320786 249748 320788
rect 66161 320784 249748 320786
rect 66161 320728 66166 320784
rect 66222 320728 249748 320784
rect 66161 320726 249748 320728
rect 66161 320723 66227 320726
rect 249742 320724 249748 320726
rect 249812 320724 249818 320788
rect -960 319290 480 319380
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 68870 316644 68876 316708
rect 68940 316706 68946 316708
rect 295926 316706 295932 316708
rect 68940 316646 295932 316706
rect 68940 316644 68946 316646
rect 295926 316644 295932 316646
rect 295996 316644 296002 316708
rect 76649 315346 76715 315349
rect 240358 315346 240364 315348
rect 76649 315344 240364 315346
rect 76649 315288 76654 315344
rect 76710 315288 240364 315344
rect 76649 315286 240364 315288
rect 76649 315283 76715 315286
rect 240358 315284 240364 315286
rect 240428 315284 240434 315348
rect 121637 314260 121703 314261
rect 121637 314256 121684 314260
rect 121748 314258 121754 314260
rect 121637 314200 121642 314256
rect 121637 314196 121684 314200
rect 121748 314198 121794 314258
rect 121748 314196 121754 314198
rect 121637 314195 121703 314196
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect 92381 307050 92447 307053
rect 268326 307050 268332 307052
rect 92381 307048 268332 307050
rect 92381 306992 92386 307048
rect 92442 306992 268332 307048
rect 92381 306990 268332 306992
rect 92381 306987 92447 306990
rect 268326 306988 268332 306990
rect 268396 306988 268402 307052
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 69054 305628 69060 305692
rect 69124 305690 69130 305692
rect 115289 305690 115355 305693
rect 69124 305688 115355 305690
rect 69124 305632 115294 305688
rect 115350 305632 115355 305688
rect 69124 305630 115355 305632
rect 69124 305628 69130 305630
rect 115289 305627 115355 305630
rect 70894 304132 70900 304196
rect 70964 304194 70970 304196
rect 94589 304194 94655 304197
rect 70964 304192 94655 304194
rect 70964 304136 94594 304192
rect 94650 304136 94655 304192
rect 70964 304134 94655 304136
rect 70964 304132 70970 304134
rect 94589 304131 94655 304134
rect 73153 302834 73219 302837
rect 249006 302834 249012 302836
rect 73153 302832 249012 302834
rect 73153 302776 73158 302832
rect 73214 302776 249012 302832
rect 73153 302774 249012 302776
rect 73153 302771 73219 302774
rect 249006 302772 249012 302774
rect 249076 302772 249082 302836
rect 113173 300794 113239 300797
rect 114461 300794 114527 300797
rect 113173 300792 114527 300794
rect 113173 300736 113178 300792
rect 113234 300736 114466 300792
rect 114522 300736 114527 300792
rect 113173 300734 114527 300736
rect 113173 300731 113239 300734
rect 114461 300731 114527 300734
rect 96521 300114 96587 300117
rect 322933 300114 322999 300117
rect 96521 300112 322999 300114
rect 96521 300056 96526 300112
rect 96582 300056 322938 300112
rect 322994 300056 322999 300112
rect 96521 300054 322999 300056
rect 96521 300051 96587 300054
rect 322933 300051 322999 300054
rect 114461 299570 114527 299573
rect 582465 299570 582531 299573
rect 114461 299568 582531 299570
rect 114461 299512 114466 299568
rect 114522 299512 582470 299568
rect 582526 299512 582531 299568
rect 114461 299510 582531 299512
rect 114461 299507 114527 299510
rect 582465 299507 582531 299510
rect 580349 298754 580415 298757
rect 583520 298754 584960 298844
rect 580349 298752 584960 298754
rect 580349 298696 580354 298752
rect 580410 298696 584960 298752
rect 580349 298694 584960 298696
rect 580349 298691 580415 298694
rect 583520 298604 584960 298694
rect 90633 298346 90699 298349
rect 247718 298346 247724 298348
rect 90633 298344 247724 298346
rect 90633 298288 90638 298344
rect 90694 298288 247724 298344
rect 90633 298286 247724 298288
rect 90633 298283 90699 298286
rect 247718 298284 247724 298286
rect 247788 298284 247794 298348
rect 70025 298210 70091 298213
rect 227662 298210 227668 298212
rect 70025 298208 227668 298210
rect 70025 298152 70030 298208
rect 70086 298152 227668 298208
rect 70025 298150 227668 298152
rect 70025 298147 70091 298150
rect 227662 298148 227668 298150
rect 227732 298148 227738 298212
rect 111057 297394 111123 297397
rect 129917 297394 129983 297397
rect 111057 297392 129983 297394
rect 111057 297336 111062 297392
rect 111118 297336 129922 297392
rect 129978 297336 129983 297392
rect 111057 297334 129983 297336
rect 111057 297331 111123 297334
rect 129917 297331 129983 297334
rect 69013 296850 69079 296853
rect 185577 296850 185643 296853
rect 69013 296848 185643 296850
rect 69013 296792 69018 296848
rect 69074 296792 185582 296848
rect 185638 296792 185643 296848
rect 69013 296790 185643 296792
rect 69013 296787 69079 296790
rect 185577 296787 185643 296790
rect 107561 296170 107627 296173
rect 127065 296170 127131 296173
rect 107561 296168 127131 296170
rect 107561 296112 107566 296168
rect 107622 296112 127070 296168
rect 127126 296112 127131 296168
rect 107561 296110 127131 296112
rect 107561 296107 107627 296110
rect 127065 296107 127131 296110
rect 76557 296034 76623 296037
rect 118734 296034 118740 296036
rect 76557 296032 118740 296034
rect 76557 295976 76562 296032
rect 76618 295976 118740 296032
rect 76557 295974 118740 295976
rect 76557 295971 76623 295974
rect 118734 295972 118740 295974
rect 118804 295972 118810 296036
rect 115841 295354 115907 295357
rect 310513 295354 310579 295357
rect 115841 295352 310579 295354
rect 115841 295296 115846 295352
rect 115902 295296 310518 295352
rect 310574 295296 310579 295352
rect 115841 295294 310579 295296
rect 115841 295291 115907 295294
rect 310513 295291 310579 295294
rect 115289 294266 115355 294269
rect 115749 294266 115815 294269
rect 123334 294266 123340 294268
rect 115289 294264 123340 294266
rect 115289 294208 115294 294264
rect 115350 294208 115754 294264
rect 115810 294208 123340 294264
rect 115289 294206 123340 294208
rect 115289 294203 115355 294206
rect 115749 294203 115815 294206
rect 123334 294204 123340 294206
rect 123404 294204 123410 294268
rect 95785 294130 95851 294133
rect 178677 294130 178743 294133
rect 95785 294128 178743 294130
rect 95785 294072 95790 294128
rect 95846 294072 178682 294128
rect 178738 294072 178743 294128
rect 95785 294070 178743 294072
rect 95785 294067 95851 294070
rect 178677 294067 178743 294070
rect 68737 293994 68803 293997
rect 287094 293994 287100 293996
rect 68737 293992 287100 293994
rect 68737 293936 68742 293992
rect 68798 293936 287100 293992
rect 68737 293934 287100 293936
rect 68737 293931 68803 293934
rect 287094 293932 287100 293934
rect 287164 293932 287170 293996
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 118601 292906 118667 292909
rect 120165 292906 120231 292909
rect 118601 292904 120231 292906
rect 118601 292848 118606 292904
rect 118662 292848 120170 292904
rect 120226 292848 120231 292904
rect 118601 292846 120231 292848
rect 118601 292843 118667 292846
rect 120165 292843 120231 292846
rect 68921 292770 68987 292773
rect 250294 292770 250300 292772
rect 68921 292768 250300 292770
rect 68921 292712 68926 292768
rect 68982 292712 250300 292768
rect 68921 292710 250300 292712
rect 68921 292707 68987 292710
rect 250294 292708 250300 292710
rect 250364 292708 250370 292772
rect 99005 292634 99071 292637
rect 304993 292634 305059 292637
rect 99005 292632 305059 292634
rect 99005 292576 99010 292632
rect 99066 292576 304998 292632
rect 305054 292576 305059 292632
rect 99005 292574 305059 292576
rect 99005 292571 99071 292574
rect 304993 292571 305059 292574
rect 71037 292362 71103 292365
rect 70718 292360 71103 292362
rect 70718 292304 71042 292360
rect 71098 292304 71103 292360
rect 70718 292302 71103 292304
rect 70718 291788 70778 292302
rect 71037 292299 71103 292302
rect 114277 291954 114343 291957
rect 164877 291954 164943 291957
rect 114277 291952 164943 291954
rect 114277 291896 114282 291952
rect 114338 291896 164882 291952
rect 164938 291896 164943 291952
rect 114277 291894 164943 291896
rect 114277 291891 114343 291894
rect 164877 291891 164943 291894
rect 121637 291818 121703 291821
rect 119876 291816 121703 291818
rect 119876 291760 121642 291816
rect 121698 291760 121703 291816
rect 119876 291758 121703 291760
rect 121637 291755 121703 291758
rect 69982 291214 70226 291274
rect 67633 291138 67699 291141
rect 69982 291138 70042 291214
rect 67633 291136 70042 291138
rect 67633 291080 67638 291136
rect 67694 291080 70042 291136
rect 70166 291108 70226 291214
rect 67633 291078 70042 291080
rect 67633 291075 67699 291078
rect 68829 290866 68895 290869
rect 68829 290864 70226 290866
rect 68829 290808 68834 290864
rect 68890 290808 70226 290864
rect 68829 290806 70226 290808
rect 68829 290803 68895 290806
rect 70166 290428 70226 290806
rect 119846 290594 119906 291108
rect 119846 290534 122850 290594
rect 121637 290458 121703 290461
rect 119876 290456 121703 290458
rect 119876 290400 121642 290456
rect 121698 290400 121703 290456
rect 119876 290398 121703 290400
rect 121637 290395 121703 290398
rect 119797 289914 119863 289917
rect 122790 289914 122850 290534
rect 242934 289914 242940 289916
rect 69982 289854 70226 289914
rect 69013 289778 69079 289781
rect 69982 289778 70042 289854
rect 69013 289776 70042 289778
rect 69013 289720 69018 289776
rect 69074 289720 70042 289776
rect 70166 289748 70226 289854
rect 119797 289912 119906 289914
rect 119797 289856 119802 289912
rect 119858 289856 119906 289912
rect 119797 289851 119906 289856
rect 122790 289854 242940 289914
rect 242934 289852 242940 289854
rect 243004 289852 243010 289916
rect 119846 289748 119906 289851
rect 69013 289718 70042 289720
rect 69013 289715 69079 289718
rect 68185 289506 68251 289509
rect 68185 289504 70226 289506
rect 68185 289448 68190 289504
rect 68246 289448 70226 289504
rect 68185 289446 70226 289448
rect 68185 289443 68251 289446
rect 70166 289068 70226 289446
rect 121729 289098 121795 289101
rect 119876 289096 121795 289098
rect 119876 289040 121734 289096
rect 121790 289040 121795 289096
rect 119876 289038 121795 289040
rect 121729 289035 121795 289038
rect 121821 288418 121887 288421
rect 119876 288416 121887 288418
rect 67633 288146 67699 288149
rect 70350 288146 70410 288388
rect 119876 288360 121826 288416
rect 121882 288360 121887 288416
rect 119876 288358 121887 288360
rect 121821 288355 121887 288358
rect 67633 288144 70410 288146
rect 67633 288088 67638 288144
rect 67694 288088 70410 288144
rect 67633 288086 70410 288088
rect 67633 288083 67699 288086
rect 121637 287738 121703 287741
rect 119876 287736 121703 287738
rect 66897 287466 66963 287469
rect 70166 287466 70226 287708
rect 119876 287680 121642 287736
rect 121698 287680 121703 287736
rect 119876 287678 121703 287680
rect 121637 287675 121703 287678
rect 66897 287464 70226 287466
rect 66897 287408 66902 287464
rect 66958 287408 70226 287464
rect 66897 287406 70226 287408
rect 66897 287403 66963 287406
rect 121637 287058 121703 287061
rect 119876 287056 121703 287058
rect 68277 286514 68343 286517
rect 70166 286514 70226 287028
rect 119876 287000 121642 287056
rect 121698 287000 121703 287056
rect 119876 286998 121703 287000
rect 121637 286995 121703 286998
rect 70526 286724 70532 286788
rect 70596 286724 70602 286788
rect 68277 286512 70226 286514
rect 68277 286456 68282 286512
rect 68338 286456 70226 286512
rect 68277 286454 70226 286456
rect 68277 286451 68343 286454
rect 70534 286348 70594 286724
rect 121545 286378 121611 286381
rect 119876 286376 121611 286378
rect 119876 286320 121550 286376
rect 121606 286320 121611 286376
rect 119876 286318 121611 286320
rect 121545 286315 121611 286318
rect 68737 286106 68803 286109
rect 68737 286104 70226 286106
rect 68737 286048 68742 286104
rect 68798 286048 70226 286104
rect 68737 286046 70226 286048
rect 68737 286043 68803 286046
rect 70166 285668 70226 286046
rect 121729 285698 121795 285701
rect 119876 285696 121795 285698
rect 119876 285640 121734 285696
rect 121790 285640 121795 285696
rect 119876 285638 121795 285640
rect 121729 285635 121795 285638
rect 68645 285426 68711 285429
rect 68645 285424 70226 285426
rect 68645 285368 68650 285424
rect 68706 285368 70226 285424
rect 68645 285366 70226 285368
rect 68645 285363 68711 285366
rect 70166 284988 70226 285366
rect 583520 285276 584960 285516
rect 121637 285018 121703 285021
rect 119876 285016 121703 285018
rect 119876 284960 121642 285016
rect 121698 284960 121703 285016
rect 119876 284958 121703 284960
rect 121637 284955 121703 284958
rect 121545 284746 121611 284749
rect 119846 284744 121611 284746
rect 119846 284688 121550 284744
rect 121606 284688 121611 284744
rect 119846 284686 121611 284688
rect 67633 284474 67699 284477
rect 67633 284472 70226 284474
rect 67633 284416 67638 284472
rect 67694 284416 70226 284472
rect 67633 284414 70226 284416
rect 67633 284411 67699 284414
rect 70166 284308 70226 284414
rect 119846 284308 119906 284686
rect 121545 284683 121611 284686
rect 68921 284066 68987 284069
rect 68921 284064 70226 284066
rect 68921 284008 68926 284064
rect 68982 284008 70226 284064
rect 68921 284006 70226 284008
rect 68921 284003 68987 284006
rect 70166 283628 70226 284006
rect 121545 283658 121611 283661
rect 119876 283656 121611 283658
rect 119876 283600 121550 283656
rect 121606 283600 121611 283656
rect 119876 283598 121611 283600
rect 121545 283595 121611 283598
rect 124806 283460 124812 283524
rect 124876 283522 124882 283524
rect 340873 283522 340939 283525
rect 124876 283520 340939 283522
rect 124876 283464 340878 283520
rect 340934 283464 340939 283520
rect 124876 283462 340939 283464
rect 124876 283460 124882 283462
rect 340873 283459 340939 283462
rect 67725 283386 67791 283389
rect 67725 283384 70226 283386
rect 67725 283328 67730 283384
rect 67786 283328 70226 283384
rect 67725 283326 70226 283328
rect 67725 283323 67791 283326
rect 70166 282948 70226 283326
rect 121545 282978 121611 282981
rect 119876 282976 121611 282978
rect 119876 282920 121550 282976
rect 121606 282920 121611 282976
rect 119876 282918 121611 282920
rect 121545 282915 121611 282918
rect 121637 282298 121703 282301
rect 119876 282296 121703 282298
rect 119876 282240 121642 282296
rect 121698 282240 121703 282296
rect 119876 282238 121703 282240
rect 121637 282235 121703 282238
rect 67633 282162 67699 282165
rect 67633 282160 70226 282162
rect 67633 282104 67638 282160
rect 67694 282104 70226 282160
rect 67633 282102 70226 282104
rect 67633 282099 67699 282102
rect 70166 281588 70226 282102
rect 121545 281618 121611 281621
rect 119876 281616 121611 281618
rect 119876 281560 121550 281616
rect 121606 281560 121611 281616
rect 119876 281558 121611 281560
rect 121545 281555 121611 281558
rect 121545 280938 121611 280941
rect 119876 280936 121611 280938
rect 68369 280530 68435 280533
rect 70166 280530 70226 280908
rect 119876 280880 121550 280936
rect 121606 280880 121611 280936
rect 119876 280878 121611 280880
rect 121545 280875 121611 280878
rect 68369 280528 70226 280530
rect 68369 280472 68374 280528
rect 68430 280472 70226 280528
rect 68369 280470 70226 280472
rect 68369 280467 68435 280470
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 241646 280258 241652 280260
rect -960 279972 480 280212
rect 119876 280198 241652 280258
rect 241646 280196 241652 280198
rect 241716 280196 241722 280260
rect 67725 279986 67791 279989
rect 67725 279984 70226 279986
rect 67725 279928 67730 279984
rect 67786 279928 70226 279984
rect 67725 279926 70226 279928
rect 67725 279923 67791 279926
rect 70166 279548 70226 279926
rect 121637 279578 121703 279581
rect 119876 279576 121703 279578
rect 119876 279520 121642 279576
rect 121698 279520 121703 279576
rect 119876 279518 121703 279520
rect 121637 279515 121703 279518
rect 67633 279306 67699 279309
rect 67633 279304 70226 279306
rect 67633 279248 67638 279304
rect 67694 279248 70226 279304
rect 67633 279246 70226 279248
rect 67633 279243 67699 279246
rect 70166 278868 70226 279246
rect 121545 278898 121611 278901
rect 119876 278896 121611 278898
rect 119876 278840 121550 278896
rect 121606 278840 121611 278896
rect 119876 278838 121611 278840
rect 121545 278835 121611 278838
rect 121637 278218 121703 278221
rect 119876 278216 121703 278218
rect 67725 277810 67791 277813
rect 70166 277810 70226 278188
rect 119876 278160 121642 278216
rect 121698 278160 121703 278216
rect 119876 278158 121703 278160
rect 121637 278155 121703 278158
rect 67725 277808 70226 277810
rect 67725 277752 67730 277808
rect 67786 277752 70226 277808
rect 67725 277750 70226 277752
rect 67725 277747 67791 277750
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 121545 277538 121611 277541
rect 119876 277536 121611 277538
rect 119876 277480 121550 277536
rect 121606 277480 121611 277536
rect 119876 277478 121611 277480
rect 121545 277475 121611 277478
rect 121545 276858 121611 276861
rect 119876 276856 121611 276858
rect 67633 276450 67699 276453
rect 70166 276450 70226 276828
rect 119876 276800 121550 276856
rect 121606 276800 121611 276856
rect 119876 276798 121611 276800
rect 121545 276795 121611 276798
rect 67633 276448 70226 276450
rect 67633 276392 67638 276448
rect 67694 276392 70226 276448
rect 67633 276390 70226 276392
rect 67633 276387 67699 276390
rect 66110 276252 66116 276316
rect 66180 276314 66186 276316
rect 66180 276254 70226 276314
rect 66180 276252 66186 276254
rect 70166 276148 70226 276254
rect 121729 276178 121795 276181
rect 119876 276176 121795 276178
rect 119876 276120 121734 276176
rect 121790 276120 121795 276176
rect 119876 276118 121795 276120
rect 121729 276115 121795 276118
rect 119286 275572 119292 275636
rect 119356 275634 119362 275636
rect 119356 275574 119906 275634
rect 119356 275572 119362 275574
rect 119846 275498 119906 275574
rect 121821 275498 121887 275501
rect 119846 275496 121887 275498
rect 119846 275468 121826 275496
rect 67817 275090 67883 275093
rect 70166 275090 70226 275468
rect 119876 275440 121826 275468
rect 121882 275440 121887 275496
rect 119876 275438 121887 275440
rect 121821 275435 121887 275438
rect 67817 275088 70226 275090
rect 67817 275032 67822 275088
rect 67878 275032 70226 275088
rect 67817 275030 70226 275032
rect 67817 275027 67883 275030
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 121545 274818 121611 274821
rect 119876 274816 121611 274818
rect 119876 274760 121550 274816
rect 121606 274760 121611 274816
rect 119876 274758 121611 274760
rect 121545 274755 121611 274758
rect 67725 274546 67791 274549
rect 67725 274544 70226 274546
rect 67725 274488 67730 274544
rect 67786 274488 70226 274544
rect 67725 274486 70226 274488
rect 67725 274483 67791 274486
rect 70166 274108 70226 274486
rect 121637 274138 121703 274141
rect 119876 274136 121703 274138
rect 119876 274080 121642 274136
rect 121698 274080 121703 274136
rect 119876 274078 121703 274080
rect 121637 274075 121703 274078
rect 67633 273594 67699 273597
rect 67633 273592 70226 273594
rect 67633 273536 67638 273592
rect 67694 273536 70226 273592
rect 67633 273534 70226 273536
rect 67633 273531 67699 273534
rect 70166 273428 70226 273534
rect 121545 273458 121611 273461
rect 119876 273456 121611 273458
rect 119876 273400 121550 273456
rect 121606 273400 121611 273456
rect 119876 273398 121611 273400
rect 121545 273395 121611 273398
rect 121637 272778 121703 272781
rect 119876 272776 121703 272778
rect 67633 272234 67699 272237
rect 70166 272234 70226 272748
rect 119876 272720 121642 272776
rect 121698 272720 121703 272776
rect 119876 272718 121703 272720
rect 121637 272715 121703 272718
rect 67633 272232 70226 272234
rect 67633 272176 67638 272232
rect 67694 272176 70226 272232
rect 67633 272174 70226 272176
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 67633 272171 67699 272174
rect 580257 272171 580323 272174
rect 121545 272098 121611 272101
rect 119876 272096 121611 272098
rect 67541 271962 67607 271965
rect 67541 271960 69858 271962
rect 67541 271904 67546 271960
rect 67602 271904 69858 271960
rect 67541 271902 69858 271904
rect 67541 271899 67607 271902
rect 69798 271826 69858 271902
rect 70350 271826 70410 272068
rect 119876 272040 121550 272096
rect 121606 272040 121611 272096
rect 583520 272084 584960 272174
rect 119876 272038 121611 272040
rect 121545 272035 121611 272038
rect 69798 271766 70410 271826
rect 121545 271418 121611 271421
rect 119876 271416 121611 271418
rect 67633 271010 67699 271013
rect 70166 271010 70226 271388
rect 119876 271360 121550 271416
rect 121606 271360 121611 271416
rect 119876 271358 121611 271360
rect 121545 271355 121611 271358
rect 67633 271008 70226 271010
rect 67633 270952 67638 271008
rect 67694 270952 70226 271008
rect 67633 270950 70226 270952
rect 67633 270947 67699 270950
rect 67725 270874 67791 270877
rect 67725 270872 70226 270874
rect 67725 270816 67730 270872
rect 67786 270816 70226 270872
rect 67725 270814 70226 270816
rect 67725 270811 67791 270814
rect 70166 270708 70226 270814
rect 121545 270058 121611 270061
rect 119876 270056 121611 270058
rect 67725 269650 67791 269653
rect 70166 269650 70226 270028
rect 119876 270000 121550 270056
rect 121606 270000 121611 270056
rect 119876 269998 121611 270000
rect 121545 269995 121611 269998
rect 67725 269648 70226 269650
rect 67725 269592 67730 269648
rect 67786 269592 70226 269648
rect 67725 269590 70226 269592
rect 67725 269587 67791 269590
rect 67633 269514 67699 269517
rect 67633 269512 70226 269514
rect 67633 269456 67638 269512
rect 67694 269456 70226 269512
rect 67633 269454 70226 269456
rect 67633 269451 67699 269454
rect 70166 269348 70226 269454
rect 121637 269378 121703 269381
rect 119876 269376 121703 269378
rect 119876 269320 121642 269376
rect 121698 269320 121703 269376
rect 119876 269318 121703 269320
rect 121637 269315 121703 269318
rect 121545 268698 121611 268701
rect 119876 268696 121611 268698
rect 69105 268290 69171 268293
rect 70166 268290 70226 268668
rect 119876 268640 121550 268696
rect 121606 268640 121611 268696
rect 119876 268638 121611 268640
rect 121545 268635 121611 268638
rect 69105 268288 70226 268290
rect 69105 268232 69110 268288
rect 69166 268232 70226 268288
rect 69105 268230 70226 268232
rect 69105 268227 69171 268230
rect 67633 268154 67699 268157
rect 67633 268152 70226 268154
rect 67633 268096 67638 268152
rect 67694 268096 70226 268152
rect 67633 268094 70226 268096
rect 67633 268091 67699 268094
rect 70166 267988 70226 268094
rect 121545 268018 121611 268021
rect 119876 268016 121611 268018
rect 119876 267960 121550 268016
rect 121606 267960 121611 268016
rect 119876 267958 121611 267960
rect 121545 267955 121611 267958
rect 67633 267474 67699 267477
rect 67633 267472 70226 267474
rect 67633 267416 67638 267472
rect 67694 267416 70226 267472
rect 67633 267414 70226 267416
rect 67633 267411 67699 267414
rect 70166 267308 70226 267414
rect 121729 267338 121795 267341
rect 119876 267336 121795 267338
rect -960 267202 480 267292
rect 119876 267280 121734 267336
rect 121790 267280 121795 267336
rect 119876 267278 121795 267280
rect 121729 267275 121795 267278
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 67725 267066 67791 267069
rect 67725 267064 70226 267066
rect 67725 267008 67730 267064
rect 67786 267008 70226 267064
rect 67725 267006 70226 267008
rect 67725 267003 67791 267006
rect 70166 266628 70226 267006
rect 121453 266658 121519 266661
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 121453 266595 121519 266598
rect 121545 265978 121611 265981
rect 119876 265976 121611 265978
rect 70166 265434 70226 265948
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 121545 265915 121611 265918
rect 64830 265374 70226 265434
rect 50838 265100 50844 265164
rect 50908 265162 50914 265164
rect 64830 265162 64890 265374
rect 121453 265298 121519 265301
rect 119876 265296 121519 265298
rect 50908 265102 64890 265162
rect 50908 265100 50914 265102
rect 67633 265026 67699 265029
rect 70350 265026 70410 265268
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 121453 265235 121519 265238
rect 67633 265024 70410 265026
rect 67633 264968 67638 265024
rect 67694 264968 70410 265024
rect 67633 264966 70410 264968
rect 67633 264963 67699 264966
rect 67633 264890 67699 264893
rect 67633 264888 70226 264890
rect 67633 264832 67638 264888
rect 67694 264832 70226 264888
rect 67633 264830 70226 264832
rect 67633 264827 67699 264830
rect 70166 264588 70226 264830
rect 121453 264618 121519 264621
rect 119876 264616 121519 264618
rect 119876 264560 121458 264616
rect 121514 264560 121519 264616
rect 119876 264558 121519 264560
rect 121453 264555 121519 264558
rect 121545 263938 121611 263941
rect 119876 263936 121611 263938
rect 67725 263666 67791 263669
rect 70166 263666 70226 263908
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 121545 263875 121611 263878
rect 67725 263664 70226 263666
rect 67725 263608 67730 263664
rect 67786 263608 70226 263664
rect 67725 263606 70226 263608
rect 67725 263603 67791 263606
rect 67633 263530 67699 263533
rect 67633 263528 70226 263530
rect 67633 263472 67638 263528
rect 67694 263472 70226 263528
rect 67633 263470 70226 263472
rect 67633 263467 67699 263470
rect 70166 263228 70226 263470
rect 121453 263258 121519 263261
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 121453 263195 121519 263198
rect 121453 262578 121519 262581
rect 119876 262576 121519 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 121453 262515 121519 262518
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121729 261898 121795 261901
rect 119876 261896 121795 261898
rect 67633 261490 67699 261493
rect 70166 261490 70226 261868
rect 119876 261840 121734 261896
rect 121790 261840 121795 261896
rect 119876 261838 121795 261840
rect 121729 261835 121795 261838
rect 67633 261488 70226 261490
rect 67633 261432 67638 261488
rect 67694 261432 70226 261488
rect 67633 261430 70226 261432
rect 67633 261427 67699 261430
rect 121545 261218 121611 261221
rect 119876 261216 121611 261218
rect 67725 260946 67791 260949
rect 70166 260946 70226 261188
rect 119876 261160 121550 261216
rect 121606 261160 121611 261216
rect 119876 261158 121611 261160
rect 121545 261155 121611 261158
rect 67725 260944 70226 260946
rect 67725 260888 67730 260944
rect 67786 260888 70226 260944
rect 67725 260886 70226 260888
rect 67725 260883 67791 260886
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121453 260538 121519 260541
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 121453 260475 121519 260478
rect 121453 259858 121519 259861
rect 119876 259856 121519 259858
rect 67633 259586 67699 259589
rect 70350 259586 70410 259828
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 121453 259795 121519 259798
rect 67633 259584 70410 259586
rect 67633 259528 67638 259584
rect 67694 259528 70410 259584
rect 67633 259526 70410 259528
rect 67633 259523 67699 259526
rect 121545 259178 121611 259181
rect 119876 259176 121611 259178
rect 67725 258634 67791 258637
rect 70166 258634 70226 259148
rect 119876 259120 121550 259176
rect 121606 259120 121611 259176
rect 119876 259118 121611 259120
rect 121545 259115 121611 259118
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 67725 258632 70226 258634
rect 67725 258576 67730 258632
rect 67786 258576 70226 258632
rect 67725 258574 70226 258576
rect 67725 258571 67791 258574
rect 121453 258498 121519 258501
rect 119876 258496 121519 258498
rect 67633 258226 67699 258229
rect 70350 258226 70410 258468
rect 119876 258440 121458 258496
rect 121514 258440 121519 258496
rect 119876 258438 121519 258440
rect 121453 258435 121519 258438
rect 67633 258224 70410 258226
rect 67633 258168 67638 258224
rect 67694 258168 70410 258224
rect 67633 258166 70410 258168
rect 67633 258163 67699 258166
rect 67633 257954 67699 257957
rect 67633 257952 70226 257954
rect 67633 257896 67638 257952
rect 67694 257896 70226 257952
rect 67633 257894 70226 257896
rect 67633 257891 67699 257894
rect 70166 257788 70226 257894
rect 121545 257818 121611 257821
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 121545 257755 121611 257758
rect 120717 257138 120783 257141
rect 119876 257136 120783 257138
rect 67633 256866 67699 256869
rect 70350 256866 70410 257108
rect 119876 257080 120722 257136
rect 120778 257080 120783 257136
rect 119876 257078 120783 257080
rect 120717 257075 120783 257078
rect 67633 256864 70410 256866
rect 67633 256808 67638 256864
rect 67694 256808 70410 256864
rect 67633 256806 70410 256808
rect 67633 256803 67699 256806
rect 120073 256458 120139 256461
rect 119876 256456 120139 256458
rect 69289 255914 69355 255917
rect 70166 255914 70226 256428
rect 119876 256400 120078 256456
rect 120134 256400 120139 256456
rect 119876 256398 120139 256400
rect 120073 256395 120139 256398
rect 69289 255912 70226 255914
rect 69289 255856 69294 255912
rect 69350 255856 70226 255912
rect 69289 255854 70226 255856
rect 69289 255851 69355 255854
rect 123334 255852 123340 255916
rect 123404 255914 123410 255916
rect 580257 255914 580323 255917
rect 123404 255912 580323 255914
rect 123404 255856 580262 255912
rect 580318 255856 580323 255912
rect 123404 255854 580323 255856
rect 123404 255852 123410 255854
rect 580257 255851 580323 255854
rect 121453 255778 121519 255781
rect 119876 255776 121519 255778
rect 67725 255370 67791 255373
rect 70166 255370 70226 255748
rect 119876 255720 121458 255776
rect 121514 255720 121519 255776
rect 119876 255718 121519 255720
rect 121453 255715 121519 255718
rect 67725 255368 70226 255370
rect 67725 255312 67730 255368
rect 67786 255312 70226 255368
rect 67725 255310 70226 255312
rect 67725 255307 67791 255310
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 121545 255098 121611 255101
rect 119876 255096 121611 255098
rect 119876 255040 121550 255096
rect 121606 255040 121611 255096
rect 119876 255038 121611 255040
rect 121545 255035 121611 255038
rect 121453 254418 121519 254421
rect 119876 254416 121519 254418
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 67725 254010 67791 254013
rect 70166 254010 70226 254388
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 121453 254355 121519 254358
rect 67725 254008 70226 254010
rect 67725 253952 67730 254008
rect 67786 253952 70226 254008
rect 67725 253950 70226 253952
rect 67725 253947 67791 253950
rect 56409 253874 56475 253877
rect 60917 253874 60983 253877
rect 61510 253874 61516 253876
rect 56409 253872 61516 253874
rect 56409 253816 56414 253872
rect 56470 253816 60922 253872
rect 60978 253816 61516 253872
rect 56409 253814 61516 253816
rect 56409 253811 56475 253814
rect 60917 253811 60983 253814
rect 61510 253812 61516 253814
rect 61580 253812 61586 253876
rect 67633 253874 67699 253877
rect 67633 253872 70226 253874
rect 67633 253816 67638 253872
rect 67694 253816 70226 253872
rect 67633 253814 70226 253816
rect 67633 253811 67699 253814
rect 70166 253708 70226 253814
rect 121545 253738 121611 253741
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 121545 253675 121611 253678
rect 126094 253132 126100 253196
rect 126164 253194 126170 253196
rect 343633 253194 343699 253197
rect 126164 253192 343699 253194
rect 126164 253136 343638 253192
rect 343694 253136 343699 253192
rect 126164 253134 343699 253136
rect 126164 253132 126170 253134
rect 343633 253131 343699 253134
rect 121453 253058 121519 253061
rect 119876 253056 121519 253058
rect 67633 252650 67699 252653
rect 70166 252650 70226 253028
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 121453 252995 121519 252998
rect 67633 252648 70226 252650
rect 67633 252592 67638 252648
rect 67694 252592 70226 252648
rect 67633 252590 70226 252592
rect 67633 252587 67699 252590
rect 121637 252378 121703 252381
rect 119876 252376 121703 252378
rect 68829 251834 68895 251837
rect 70166 251834 70226 252348
rect 119876 252320 121642 252376
rect 121698 252320 121703 252376
rect 119876 252318 121703 252320
rect 121637 252315 121703 252318
rect 68829 251832 70226 251834
rect 68829 251776 68834 251832
rect 68890 251776 70226 251832
rect 68829 251774 70226 251776
rect 68829 251771 68895 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 57830 251364 57836 251428
rect 57900 251426 57906 251428
rect 70166 251426 70226 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 57900 251366 70226 251426
rect 57900 251364 57906 251366
rect 120073 251018 120139 251021
rect 122925 251018 122991 251021
rect 119876 251016 122991 251018
rect 65926 250412 65932 250476
rect 65996 250474 66002 250476
rect 70166 250474 70226 250988
rect 119876 250960 120078 251016
rect 120134 250960 122930 251016
rect 122986 250960 122991 251016
rect 119876 250958 122991 250960
rect 120073 250955 120139 250958
rect 122925 250955 122991 250958
rect 65996 250414 70226 250474
rect 65996 250412 66002 250414
rect 121545 250338 121611 250341
rect 119876 250336 121611 250338
rect 67725 249930 67791 249933
rect 70166 249930 70226 250308
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 121545 250275 121611 250278
rect 67725 249928 70226 249930
rect 67725 249872 67730 249928
rect 67786 249872 70226 249928
rect 67725 249870 70226 249872
rect 67725 249867 67791 249870
rect 67633 249794 67699 249797
rect 67633 249792 70226 249794
rect 67633 249736 67638 249792
rect 67694 249736 70226 249792
rect 67633 249734 70226 249736
rect 67633 249731 67699 249734
rect 70166 249628 70226 249734
rect 121453 249658 121519 249661
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 121453 249595 121519 249598
rect 121453 248978 121519 248981
rect 119876 248976 121519 248978
rect 70534 248436 70594 248948
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 121453 248915 121519 248918
rect 70526 248372 70532 248436
rect 70596 248372 70602 248436
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67633 247754 67699 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67633 247752 70226 247754
rect 67633 247696 67638 247752
rect 67694 247696 70226 247752
rect 67633 247694 70226 247696
rect 67633 247691 67699 247694
rect 122741 247618 122807 247621
rect 119876 247616 122807 247618
rect 67725 247210 67791 247213
rect 70166 247210 70226 247588
rect 119876 247560 122746 247616
rect 122802 247560 122807 247616
rect 119876 247558 122807 247560
rect 122741 247555 122807 247558
rect 67725 247208 70226 247210
rect 67725 247152 67730 247208
rect 67786 247152 70226 247208
rect 67725 247150 70226 247152
rect 67725 247147 67791 247150
rect 67633 246666 67699 246669
rect 70350 246666 70410 246908
rect 67633 246664 70410 246666
rect 67633 246608 67638 246664
rect 67694 246608 70410 246664
rect 67633 246606 70410 246608
rect 67633 246603 67699 246606
rect 119846 246394 119906 246908
rect 120022 246468 120028 246532
rect 120092 246530 120098 246532
rect 120092 246470 132510 246530
rect 120092 246468 120098 246470
rect 132450 246394 132510 246470
rect 580349 246394 580415 246397
rect 119846 246334 122850 246394
rect 132450 246392 580415 246394
rect 132450 246336 580354 246392
rect 580410 246336 580415 246392
rect 132450 246334 580415 246336
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 69013 245714 69079 245717
rect 70166 245714 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 69013 245712 70226 245714
rect 69013 245656 69018 245712
rect 69074 245656 70226 245712
rect 69013 245654 70226 245656
rect 122790 245714 122850 246334
rect 580349 246331 580415 246334
rect 240542 245714 240548 245716
rect 122790 245654 240548 245714
rect 69013 245651 69079 245654
rect 240542 245652 240548 245654
rect 240612 245652 240618 245716
rect 121545 245578 121611 245581
rect 119876 245576 121611 245578
rect 67633 245306 67699 245309
rect 70350 245306 70410 245548
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 121545 245515 121611 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 67633 245304 70410 245306
rect 67633 245248 67638 245304
rect 67694 245248 70410 245304
rect 67633 245246 70410 245248
rect 67633 245243 67699 245246
rect 120165 244898 120231 244901
rect 119876 244896 120231 244898
rect 67633 244626 67699 244629
rect 70166 244626 70226 244868
rect 119876 244840 120170 244896
rect 120226 244840 120231 244896
rect 119876 244838 120231 244840
rect 120165 244835 120231 244838
rect 67633 244624 70226 244626
rect 67633 244568 67638 244624
rect 67694 244568 70226 244624
rect 67633 244566 70226 244568
rect 67633 244563 67699 244566
rect 69982 244294 70226 244354
rect 67817 244218 67883 244221
rect 69982 244218 70042 244294
rect 67817 244216 70042 244218
rect 67817 244160 67822 244216
rect 67878 244160 70042 244216
rect 70166 244188 70226 244294
rect 121545 244218 121611 244221
rect 119876 244216 121611 244218
rect 67817 244158 70042 244160
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 67817 244155 67883 244158
rect 121545 244155 121611 244158
rect 67725 243946 67791 243949
rect 67725 243944 70226 243946
rect 67725 243888 67730 243944
rect 67786 243888 70226 243944
rect 67725 243886 70226 243888
rect 67725 243883 67791 243886
rect 70166 243508 70226 243886
rect 121453 243538 121519 243541
rect 119876 243536 121519 243538
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 121453 243475 121519 243478
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 67633 242586 67699 242589
rect 70350 242586 70410 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 67633 242584 70410 242586
rect 67633 242528 67638 242584
rect 67694 242528 70410 242584
rect 67633 242526 70410 242528
rect 67633 242523 67699 242526
rect 121545 242178 121611 242181
rect 119876 242176 121611 242178
rect 67633 241906 67699 241909
rect 70166 241906 70226 242148
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 121545 242115 121611 242118
rect 67633 241904 70226 241906
rect 67633 241848 67638 241904
rect 67694 241848 70226 241904
rect 67633 241846 70226 241848
rect 67633 241843 67699 241846
rect 122097 241498 122163 241501
rect 119876 241496 122163 241498
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 70166 240954 70226 241468
rect 119876 241440 122102 241496
rect 122158 241440 122163 241496
rect 119876 241438 122163 241440
rect 122097 241435 122163 241438
rect 64830 240894 70226 240954
rect 119981 240954 120047 240957
rect 129825 240954 129891 240957
rect 119981 240952 129891 240954
rect 119981 240896 119986 240952
rect 120042 240896 129830 240952
rect 129886 240896 129891 240952
rect 119981 240894 129891 240896
rect 59118 240348 59124 240412
rect 59188 240410 59194 240412
rect 64830 240410 64890 240894
rect 119981 240891 120047 240894
rect 129825 240891 129891 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 67633 240546 67699 240549
rect 70166 240546 70226 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 67633 240544 70226 240546
rect 67633 240488 67638 240544
rect 67694 240488 70226 240544
rect 67633 240486 70226 240488
rect 67633 240483 67699 240486
rect 59188 240350 64890 240410
rect 59188 240348 59194 240350
rect 122373 240138 122439 240141
rect 119876 240136 122439 240138
rect 119876 240080 122378 240136
rect 122434 240080 122439 240136
rect 119876 240078 122439 240080
rect 122373 240075 122439 240078
rect 103513 238778 103579 238781
rect 104801 238778 104867 238781
rect 103513 238776 104867 238778
rect 103513 238720 103518 238776
rect 103574 238720 104806 238776
rect 104862 238720 104867 238776
rect 103513 238718 104867 238720
rect 103513 238715 103579 238718
rect 104801 238715 104867 238718
rect 75821 238642 75887 238645
rect 138013 238642 138079 238645
rect 75821 238640 138079 238642
rect 75821 238584 75826 238640
rect 75882 238584 138018 238640
rect 138074 238584 138079 238640
rect 75821 238582 138079 238584
rect 75821 238579 75887 238582
rect 138013 238579 138079 238582
rect 61326 238444 61332 238508
rect 61396 238506 61402 238508
rect 86217 238506 86283 238509
rect 61396 238504 86283 238506
rect 61396 238448 86222 238504
rect 86278 238448 86283 238504
rect 61396 238446 86283 238448
rect 61396 238444 61402 238446
rect 86217 238443 86283 238446
rect 91921 238506 91987 238509
rect 119286 238506 119292 238508
rect 91921 238504 119292 238506
rect 91921 238448 91926 238504
rect 91982 238448 119292 238504
rect 91921 238446 119292 238448
rect 91921 238443 91987 238446
rect 119286 238444 119292 238446
rect 119356 238444 119362 238508
rect 61510 235180 61516 235244
rect 61580 235242 61586 235244
rect 582741 235242 582807 235245
rect 61580 235240 582807 235242
rect 61580 235184 582746 235240
rect 582802 235184 582807 235240
rect 61580 235182 582807 235184
rect 61580 235180 61586 235182
rect 582741 235179 582807 235182
rect 580533 232386 580599 232389
rect 583520 232386 584960 232476
rect 580533 232384 584960 232386
rect 580533 232328 580538 232384
rect 580594 232328 584960 232384
rect 580533 232326 584960 232328
rect 580533 232323 580599 232326
rect 583520 232236 584960 232326
rect 75913 228306 75979 228309
rect 288566 228306 288572 228308
rect 75913 228304 288572 228306
rect 75913 228248 75918 228304
rect 75974 228248 288572 228304
rect 75913 228246 288572 228248
rect 75913 228243 75979 228246
rect 288566 228244 288572 228246
rect 288636 228244 288642 228308
rect -960 227884 480 228124
rect 66069 227082 66135 227085
rect 230422 227082 230428 227084
rect 66069 227080 230428 227082
rect 66069 227024 66074 227080
rect 66130 227024 230428 227080
rect 66069 227022 230428 227024
rect 66069 227019 66135 227022
rect 230422 227020 230428 227022
rect 230492 227020 230498 227084
rect 84377 226946 84443 226949
rect 285622 226946 285628 226948
rect 84377 226944 285628 226946
rect 84377 226888 84382 226944
rect 84438 226888 285628 226944
rect 84377 226886 285628 226888
rect 84377 226883 84443 226886
rect 285622 226884 285628 226886
rect 285692 226884 285698 226948
rect 133873 226268 133939 226269
rect 133822 226266 133828 226268
rect 133782 226206 133828 226266
rect 133892 226264 133939 226268
rect 133934 226208 133939 226264
rect 133822 226204 133828 226206
rect 133892 226204 133939 226208
rect 133873 226203 133939 226204
rect 50838 225524 50844 225588
rect 50908 225586 50914 225588
rect 298093 225586 298159 225589
rect 50908 225584 298159 225586
rect 50908 225528 298098 225584
rect 298154 225528 298159 225584
rect 50908 225526 298159 225528
rect 50908 225524 50914 225526
rect 298093 225523 298159 225526
rect 49509 222866 49575 222869
rect 291326 222866 291332 222868
rect 49509 222864 291332 222866
rect 49509 222808 49514 222864
rect 49570 222808 291332 222864
rect 49509 222806 291332 222808
rect 49509 222803 49575 222806
rect 291326 222804 291332 222806
rect 291396 222804 291402 222868
rect 582557 219058 582623 219061
rect 583520 219058 584960 219148
rect 582557 219056 584960 219058
rect 582557 219000 582562 219056
rect 582618 219000 584960 219056
rect 582557 218998 584960 219000
rect 582557 218995 582623 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 99465 213210 99531 213213
rect 278814 213210 278820 213212
rect 99465 213208 278820 213210
rect 99465 213152 99470 213208
rect 99526 213152 278820 213208
rect 99465 213150 278820 213152
rect 99465 213147 99531 213150
rect 278814 213148 278820 213150
rect 278884 213148 278890 213212
rect 87045 208994 87111 208997
rect 285806 208994 285812 208996
rect 87045 208992 285812 208994
rect 87045 208936 87050 208992
rect 87106 208936 285812 208992
rect 87045 208934 285812 208936
rect 87045 208931 87111 208934
rect 285806 208932 285812 208934
rect 285876 208932 285882 208996
rect 580441 205730 580507 205733
rect 583520 205730 584960 205820
rect 580441 205728 584960 205730
rect 580441 205672 580446 205728
rect 580502 205672 584960 205728
rect 580441 205670 584960 205672
rect 580441 205667 580507 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 74533 197978 74599 197981
rect 233182 197978 233188 197980
rect 74533 197976 233188 197978
rect 74533 197920 74538 197976
rect 74594 197920 233188 197976
rect 74533 197918 233188 197920
rect 74533 197915 74599 197918
rect 233182 197916 233188 197918
rect 233252 197916 233258 197980
rect 63125 196754 63191 196757
rect 236494 196754 236500 196756
rect 63125 196752 236500 196754
rect 63125 196696 63130 196752
rect 63186 196696 236500 196752
rect 63125 196694 236500 196696
rect 63125 196691 63191 196694
rect 236494 196692 236500 196694
rect 236564 196692 236570 196756
rect 65926 196556 65932 196620
rect 65996 196618 66002 196620
rect 298185 196618 298251 196621
rect 65996 196616 298251 196618
rect 65996 196560 298190 196616
rect 298246 196560 298251 196616
rect 65996 196558 298251 196560
rect 65996 196556 66002 196558
rect 298185 196555 298251 196558
rect 78673 192538 78739 192541
rect 280286 192538 280292 192540
rect 78673 192536 280292 192538
rect 78673 192480 78678 192536
rect 78734 192480 280292 192536
rect 78673 192478 280292 192480
rect 78673 192475 78739 192478
rect 280286 192476 280292 192478
rect 280356 192476 280362 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 141417 191042 141483 191045
rect 237598 191042 237604 191044
rect 141417 191040 237604 191042
rect 141417 190984 141422 191040
rect 141478 190984 237604 191040
rect 141417 190982 237604 190984
rect 141417 190979 141483 190982
rect 237598 190980 237604 190982
rect 237668 190980 237674 191044
rect 77293 189682 77359 189685
rect 287278 189682 287284 189684
rect 77293 189680 287284 189682
rect 77293 189624 77298 189680
rect 77354 189624 287284 189680
rect 77293 189622 287284 189624
rect 77293 189619 77359 189622
rect 287278 189620 287284 189622
rect 287348 189620 287354 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 171777 187098 171843 187101
rect 290590 187098 290596 187100
rect 171777 187096 290596 187098
rect 171777 187040 171782 187096
rect 171838 187040 290596 187096
rect 171777 187038 290596 187040
rect 171777 187035 171843 187038
rect 290590 187036 290596 187038
rect 290660 187036 290666 187100
rect 57789 186962 57855 186965
rect 237414 186962 237420 186964
rect 57789 186960 237420 186962
rect 57789 186904 57794 186960
rect 57850 186904 237420 186960
rect 57789 186902 237420 186904
rect 57789 186899 57855 186902
rect 237414 186900 237420 186902
rect 237484 186900 237490 186964
rect 66110 184180 66116 184244
rect 66180 184242 66186 184244
rect 281809 184242 281875 184245
rect 66180 184240 281875 184242
rect 66180 184184 281814 184240
rect 281870 184184 281875 184240
rect 66180 184182 281875 184184
rect 66180 184180 66186 184182
rect 281809 184179 281875 184182
rect 67357 182882 67423 182885
rect 245878 182882 245884 182884
rect 67357 182880 245884 182882
rect 67357 182824 67362 182880
rect 67418 182824 245884 182880
rect 67357 182822 245884 182824
rect 67357 182819 67423 182822
rect 245878 182820 245884 182822
rect 245948 182820 245954 182884
rect 164877 181386 164943 181389
rect 189717 181386 189783 181389
rect 164877 181384 189783 181386
rect 164877 181328 164882 181384
rect 164938 181328 189722 181384
rect 189778 181328 189783 181384
rect 164877 181326 189783 181328
rect 164877 181323 164943 181326
rect 189717 181323 189783 181326
rect 70894 180100 70900 180164
rect 70964 180162 70970 180164
rect 259453 180162 259519 180165
rect 70964 180160 259519 180162
rect 70964 180104 259458 180160
rect 259514 180104 259519 180160
rect 70964 180102 259519 180104
rect 70964 180100 70970 180102
rect 259453 180099 259519 180102
rect 67449 180026 67515 180029
rect 305269 180026 305335 180029
rect 67449 180024 305335 180026
rect 67449 179968 67454 180024
rect 67510 179968 305274 180024
rect 305330 179968 305335 180024
rect 67449 179966 305335 179968
rect 67449 179963 67515 179966
rect 305269 179963 305335 179966
rect 110137 179482 110203 179485
rect 166206 179482 166212 179484
rect 110137 179480 166212 179482
rect 110137 179424 110142 179480
rect 110198 179424 166212 179480
rect 110137 179422 166212 179424
rect 110137 179419 110203 179422
rect 166206 179420 166212 179422
rect 166276 179420 166282 179484
rect 582833 179210 582899 179213
rect 583520 179210 584960 179300
rect 582833 179208 584960 179210
rect 582833 179152 582838 179208
rect 582894 179152 584960 179208
rect 582833 179150 584960 179152
rect 582833 179147 582899 179150
rect 583520 179060 584960 179150
rect 269113 178802 269179 178805
rect 294270 178802 294276 178804
rect 269113 178800 294276 178802
rect 269113 178744 269118 178800
rect 269174 178744 294276 178800
rect 269113 178742 294276 178744
rect 269113 178739 269179 178742
rect 294270 178740 294276 178742
rect 294340 178740 294346 178804
rect 238017 178666 238083 178669
rect 295374 178666 295380 178668
rect 238017 178664 295380 178666
rect 238017 178608 238022 178664
rect 238078 178608 295380 178664
rect 238017 178606 295380 178608
rect 238017 178603 238083 178606
rect 295374 178604 295380 178606
rect 295444 178604 295450 178668
rect 97022 177652 97028 177716
rect 97092 177714 97098 177716
rect 97717 177714 97783 177717
rect 97092 177712 97783 177714
rect 97092 177656 97722 177712
rect 97778 177656 97783 177712
rect 97092 177654 97783 177656
rect 97092 177652 97098 177654
rect 97717 177651 97783 177654
rect 98310 177652 98316 177716
rect 98380 177714 98386 177716
rect 99281 177714 99347 177717
rect 98380 177712 99347 177714
rect 98380 177656 99286 177712
rect 99342 177656 99347 177712
rect 98380 177654 99347 177656
rect 98380 177652 98386 177654
rect 99281 177651 99347 177654
rect 100702 177652 100708 177716
rect 100772 177714 100778 177716
rect 101949 177714 102015 177717
rect 100772 177712 102015 177714
rect 100772 177656 101954 177712
rect 102010 177656 102015 177712
rect 100772 177654 102015 177656
rect 100772 177652 100778 177654
rect 101949 177651 102015 177654
rect 104566 177652 104572 177716
rect 104636 177714 104642 177716
rect 104801 177714 104867 177717
rect 104636 177712 104867 177714
rect 104636 177656 104806 177712
rect 104862 177656 104867 177712
rect 104636 177654 104867 177656
rect 104636 177652 104642 177654
rect 104801 177651 104867 177654
rect 113214 177652 113220 177716
rect 113284 177714 113290 177716
rect 114093 177714 114159 177717
rect 113284 177712 114159 177714
rect 113284 177656 114098 177712
rect 114154 177656 114159 177712
rect 113284 177654 114159 177656
rect 113284 177652 113290 177654
rect 114093 177651 114159 177654
rect 114318 177652 114324 177716
rect 114388 177714 114394 177716
rect 114461 177714 114527 177717
rect 118417 177716 118483 177717
rect 118366 177714 118372 177716
rect 114388 177712 114527 177714
rect 114388 177656 114466 177712
rect 114522 177656 114527 177712
rect 114388 177654 114527 177656
rect 118326 177654 118372 177714
rect 118436 177712 118483 177716
rect 118478 177656 118483 177712
rect 114388 177652 114394 177654
rect 114461 177651 114527 177654
rect 118366 177652 118372 177654
rect 118436 177652 118483 177656
rect 119470 177652 119476 177716
rect 119540 177714 119546 177716
rect 119981 177714 120047 177717
rect 119540 177712 120047 177714
rect 119540 177656 119986 177712
rect 120042 177656 120047 177712
rect 119540 177654 120047 177656
rect 119540 177652 119546 177654
rect 118417 177651 118483 177652
rect 119981 177651 120047 177654
rect 121862 177652 121868 177716
rect 121932 177714 121938 177716
rect 122649 177714 122715 177717
rect 121932 177712 122715 177714
rect 121932 177656 122654 177712
rect 122710 177656 122715 177712
rect 121932 177654 122715 177656
rect 121932 177652 121938 177654
rect 122649 177651 122715 177654
rect 127014 177652 127020 177716
rect 127084 177714 127090 177716
rect 128261 177714 128327 177717
rect 129457 177716 129523 177717
rect 129406 177714 129412 177716
rect 127084 177712 128327 177714
rect 127084 177656 128266 177712
rect 128322 177656 128327 177712
rect 127084 177654 128327 177656
rect 129366 177654 129412 177714
rect 129476 177712 129523 177716
rect 129518 177656 129523 177712
rect 127084 177652 127090 177654
rect 128261 177651 128327 177654
rect 129406 177652 129412 177654
rect 129476 177652 129523 177656
rect 129457 177651 129523 177652
rect 227069 177578 227135 177581
rect 234654 177578 234660 177580
rect 227069 177576 234660 177578
rect 227069 177520 227074 177576
rect 227130 177520 234660 177576
rect 227069 177518 234660 177520
rect 227069 177515 227135 177518
rect 234654 177516 234660 177518
rect 234724 177516 234730 177580
rect 160737 177442 160803 177445
rect 193857 177442 193923 177445
rect 160737 177440 193923 177442
rect 160737 177384 160742 177440
rect 160798 177384 193862 177440
rect 193918 177384 193923 177440
rect 160737 177382 193923 177384
rect 160737 177379 160803 177382
rect 193857 177379 193923 177382
rect 206461 177442 206527 177445
rect 228950 177442 228956 177444
rect 206461 177440 228956 177442
rect 206461 177384 206466 177440
rect 206522 177384 228956 177440
rect 206461 177382 228956 177384
rect 206461 177379 206527 177382
rect 228950 177380 228956 177382
rect 229020 177380 229026 177444
rect 265617 177442 265683 177445
rect 291285 177442 291351 177445
rect 265617 177440 291351 177442
rect 265617 177384 265622 177440
rect 265678 177384 291290 177440
rect 291346 177384 291351 177440
rect 265617 177382 291351 177384
rect 265617 177379 265683 177382
rect 291285 177379 291351 177382
rect 181437 177306 181503 177309
rect 238518 177306 238524 177308
rect 181437 177304 238524 177306
rect 181437 177248 181442 177304
rect 181498 177248 238524 177304
rect 181437 177246 238524 177248
rect 181437 177243 181503 177246
rect 238518 177244 238524 177246
rect 238588 177244 238594 177308
rect 258717 177306 258783 177309
rect 329833 177306 329899 177309
rect 258717 177304 329899 177306
rect 258717 177248 258722 177304
rect 258778 177248 329838 177304
rect 329894 177248 329899 177304
rect 258717 177246 329899 177248
rect 258717 177243 258783 177246
rect 329833 177243 329899 177246
rect 278773 177170 278839 177173
rect 279366 177170 279372 177172
rect 278773 177168 279372 177170
rect 278773 177112 278778 177168
rect 278834 177112 279372 177168
rect 278773 177110 279372 177112
rect 278773 177107 278839 177110
rect 279366 177108 279372 177110
rect 279436 177108 279442 177172
rect 109534 176972 109540 177036
rect 109604 177034 109610 177036
rect 110137 177034 110203 177037
rect 109604 177032 110203 177034
rect 109604 176976 110142 177032
rect 110198 176976 110203 177032
rect 109604 176974 110203 176976
rect 109604 176972 109610 176974
rect 110137 176971 110203 176974
rect 125726 176972 125732 177036
rect 125796 177034 125802 177036
rect 126789 177034 126855 177037
rect 133137 177036 133203 177037
rect 133086 177034 133092 177036
rect 125796 177032 126855 177034
rect 125796 176976 126794 177032
rect 126850 176976 126855 177032
rect 125796 176974 126855 176976
rect 133046 176974 133092 177034
rect 133156 177032 133203 177036
rect 133198 176976 133203 177032
rect 125796 176972 125802 176974
rect 126789 176971 126855 176974
rect 133086 176972 133092 176974
rect 133156 176972 133203 176976
rect 133137 176971 133203 176972
rect 100661 176762 100727 176765
rect 102041 176764 102107 176765
rect 101990 176762 101996 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 103329 176762 103395 176765
rect 105721 176764 105787 176765
rect 107009 176764 107075 176765
rect 108113 176764 108179 176765
rect 115841 176764 115907 176765
rect 105670 176762 105676 176764
rect 102102 176704 102107 176760
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 102041 176699 102107 176700
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 105630 176702 105676 176762
rect 105740 176760 105787 176764
rect 106958 176762 106964 176764
rect 105782 176704 105787 176760
rect 105670 176700 105676 176702
rect 105740 176700 105787 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 108062 176762 108068 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 115790 176762 115796 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 115902 176704 115907 176760
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 123150 176700 123156 176764
rect 123220 176762 123226 176764
rect 123753 176762 123819 176765
rect 128169 176762 128235 176765
rect 130745 176764 130811 176765
rect 132401 176764 132467 176765
rect 130694 176762 130700 176764
rect 123220 176760 123819 176762
rect 123220 176704 123758 176760
rect 123814 176704 123819 176760
rect 123220 176702 123819 176704
rect 123220 176700 123226 176702
rect 105721 176699 105787 176700
rect 107009 176699 107075 176700
rect 108113 176699 108179 176700
rect 115841 176699 115907 176700
rect 123753 176699 123819 176702
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 130654 176702 130700 176762
rect 130764 176760 130811 176764
rect 132350 176762 132356 176764
rect 130806 176704 130811 176760
rect 130694 176700 130700 176702
rect 130764 176700 130811 176704
rect 132310 176702 132356 176762
rect 132420 176760 132467 176764
rect 132462 176704 132467 176760
rect 132350 176700 132356 176702
rect 132420 176700 132467 176704
rect 134374 176700 134380 176764
rect 134444 176762 134450 176764
rect 134793 176762 134859 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 136030 176762 136036 176764
rect 134444 176760 134859 176762
rect 134444 176704 134798 176760
rect 134854 176704 134859 176760
rect 134444 176702 134859 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 134444 176700 134450 176702
rect 130745 176699 130811 176700
rect 132401 176699 132467 176700
rect 134793 176699 134859 176702
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 103286 176492 103346 176699
rect 128126 176492 128186 176699
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 278037 176218 278103 176221
rect 281574 176218 281580 176220
rect 278037 176216 281580 176218
rect 278037 176160 278042 176216
rect 278098 176160 281580 176216
rect 278037 176158 281580 176160
rect 278037 176155 278103 176158
rect 281574 176156 281580 176158
rect 281644 176156 281650 176220
rect -960 175796 480 176036
rect 202229 175946 202295 175949
rect 229502 175946 229508 175948
rect 202229 175944 229508 175946
rect 202229 175888 202234 175944
rect 202290 175888 229508 175944
rect 202229 175886 229508 175888
rect 202229 175883 202295 175886
rect 229502 175884 229508 175886
rect 229572 175884 229578 175948
rect 213821 175810 213887 175813
rect 227713 175810 227779 175813
rect 264421 175810 264487 175813
rect 268510 175810 268516 175812
rect 213821 175808 217242 175810
rect 213821 175752 213826 175808
rect 213882 175752 217242 175808
rect 213821 175750 217242 175752
rect 213821 175747 213887 175750
rect 217182 175644 217242 175750
rect 227713 175808 228282 175810
rect 227713 175752 227718 175808
rect 227774 175752 228282 175808
rect 227713 175750 228282 175752
rect 227713 175747 227779 175750
rect 228222 175644 228282 175750
rect 264421 175808 268516 175810
rect 264421 175752 264426 175808
rect 264482 175752 268516 175808
rect 264421 175750 268516 175752
rect 264421 175747 264487 175750
rect 268510 175748 268516 175750
rect 268580 175748 268586 175812
rect 269941 175810 270007 175813
rect 269941 175808 279434 175810
rect 269941 175752 269946 175808
rect 270002 175752 279434 175808
rect 269941 175750 279434 175752
rect 269941 175747 270007 175750
rect 116945 175540 117011 175541
rect 120809 175540 120875 175541
rect 124489 175540 124555 175541
rect 158897 175540 158963 175541
rect 116894 175538 116900 175540
rect 116854 175478 116900 175538
rect 116964 175536 117011 175540
rect 120758 175538 120764 175540
rect 117006 175480 117011 175536
rect 116894 175476 116900 175478
rect 116964 175476 117011 175480
rect 120718 175478 120764 175538
rect 120828 175536 120875 175540
rect 124438 175538 124444 175540
rect 120870 175480 120875 175536
rect 120758 175476 120764 175478
rect 120828 175476 120875 175480
rect 124398 175478 124444 175538
rect 124508 175536 124555 175540
rect 158846 175538 158852 175540
rect 124550 175480 124555 175536
rect 124438 175476 124444 175478
rect 124508 175476 124555 175480
rect 158806 175478 158852 175538
rect 158916 175536 158963 175540
rect 158958 175480 158963 175536
rect 158846 175476 158852 175478
rect 158916 175476 158963 175480
rect 116945 175475 117011 175476
rect 120809 175475 120875 175476
rect 124489 175475 124555 175476
rect 158897 175475 158963 175476
rect 110689 175404 110755 175405
rect 110638 175402 110644 175404
rect 110598 175342 110644 175402
rect 110708 175400 110755 175404
rect 110750 175344 110755 175400
rect 110638 175340 110644 175342
rect 110708 175340 110755 175344
rect 112110 175340 112116 175404
rect 112180 175402 112186 175404
rect 166390 175402 166396 175404
rect 112180 175342 166396 175402
rect 112180 175340 112186 175342
rect 166390 175340 166396 175342
rect 166460 175340 166466 175404
rect 267089 175402 267155 175405
rect 268150 175402 268210 175644
rect 279374 175508 279434 175750
rect 267089 175400 268210 175402
rect 267089 175344 267094 175400
rect 267150 175344 268210 175400
rect 267089 175342 268210 175344
rect 110689 175339 110755 175340
rect 267089 175339 267155 175342
rect 228896 175162 229202 175222
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 217182 174964 217242 175070
rect 229142 174996 229202 175162
rect 229134 174932 229140 174996
rect 229204 174932 229210 174996
rect 265709 174994 265775 174997
rect 268150 174994 268210 175236
rect 279366 175204 279372 175268
rect 279436 175204 279442 175268
rect 265709 174992 268210 174994
rect 265709 174936 265714 174992
rect 265770 174936 268210 174992
rect 265709 174934 268210 174936
rect 265709 174931 265775 174934
rect 268510 174932 268516 174996
rect 268580 174932 268586 174996
rect 268518 174828 268578 174932
rect 214005 174722 214071 174725
rect 229093 174722 229159 174725
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 228968 174720 229159 174722
rect 228968 174664 229098 174720
rect 229154 174664 229159 174720
rect 279374 174692 279434 175204
rect 228968 174662 229159 174664
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 229093 174659 229159 174662
rect 267966 174526 268210 174586
rect 261477 174450 261543 174453
rect 267966 174450 268026 174526
rect 261477 174448 268026 174450
rect 261477 174392 261482 174448
rect 261538 174392 268026 174448
rect 268150 174420 268210 174526
rect 261477 174390 268026 174392
rect 261477 174387 261543 174390
rect 229134 174314 229140 174316
rect 228968 174254 229140 174314
rect 229134 174252 229140 174254
rect 229204 174252 229210 174316
rect 265801 174178 265867 174181
rect 265801 174176 268210 174178
rect 265801 174120 265806 174176
rect 265862 174120 268210 174176
rect 265801 174118 268210 174120
rect 265801 174115 265867 174118
rect 268150 174012 268210 174118
rect 281809 174042 281875 174045
rect 279956 174040 281875 174042
rect 279956 173984 281814 174040
rect 281870 173984 281875 174040
rect 279956 173982 281875 173984
rect 281809 173979 281875 173982
rect 213913 173770 213979 173773
rect 231761 173770 231827 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 228968 173768 231827 173770
rect 228968 173712 231766 173768
rect 231822 173712 231827 173768
rect 228968 173710 231827 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 231761 173707 231827 173710
rect 279325 173770 279391 173773
rect 279325 173768 279434 173770
rect 279325 173712 279330 173768
rect 279386 173712 279434 173768
rect 279325 173707 279434 173712
rect 214097 173362 214163 173365
rect 231117 173362 231183 173365
rect 214097 173360 217242 173362
rect 214097 173304 214102 173360
rect 214158 173304 217242 173360
rect 214097 173302 217242 173304
rect 228968 173360 231183 173362
rect 228968 173304 231122 173360
rect 231178 173304 231183 173360
rect 228968 173302 231183 173304
rect 214097 173299 214163 173302
rect 217182 172924 217242 173302
rect 231117 173299 231183 173302
rect 265893 173226 265959 173229
rect 268150 173226 268210 173604
rect 265893 173224 268210 173226
rect 265893 173168 265898 173224
rect 265954 173168 268210 173224
rect 279374 173196 279434 173707
rect 265893 173166 268210 173168
rect 265893 173163 265959 173166
rect 231485 172818 231551 172821
rect 228968 172816 231551 172818
rect 228968 172760 231490 172816
rect 231546 172760 231551 172816
rect 228968 172758 231551 172760
rect 231485 172755 231551 172758
rect 265525 172818 265591 172821
rect 268150 172818 268210 173060
rect 265525 172816 268210 172818
rect 265525 172760 265530 172816
rect 265586 172760 268210 172816
rect 265525 172758 268210 172760
rect 265525 172755 265591 172758
rect 265709 172546 265775 172549
rect 265709 172544 267842 172546
rect 265709 172488 265714 172544
rect 265770 172488 267842 172544
rect 265709 172486 267842 172488
rect 265709 172483 265775 172486
rect 213913 172410 213979 172413
rect 229185 172410 229251 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 228968 172408 229251 172410
rect 228968 172352 229190 172408
rect 229246 172352 229251 172408
rect 228968 172350 229251 172352
rect 267782 172410 267842 172486
rect 268334 172410 268394 172652
rect 282085 172410 282151 172413
rect 267782 172350 268394 172410
rect 279956 172408 282151 172410
rect 279956 172352 282090 172408
rect 282146 172352 282151 172408
rect 279956 172350 282151 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 229185 172347 229251 172350
rect 282085 172347 282151 172350
rect 214005 172002 214071 172005
rect 265893 172002 265959 172005
rect 268150 172002 268210 172244
rect 214005 172000 217242 172002
rect 214005 171944 214010 172000
rect 214066 171944 217242 172000
rect 214005 171942 217242 171944
rect 214005 171939 214071 171942
rect 167545 171594 167611 171597
rect 164694 171592 167611 171594
rect 164694 171536 167550 171592
rect 167606 171536 167611 171592
rect 217182 171564 217242 171942
rect 265893 172000 268210 172002
rect 265893 171944 265898 172000
rect 265954 171944 268210 172000
rect 265893 171942 268210 171944
rect 265893 171939 265959 171942
rect 231761 171866 231827 171869
rect 228968 171864 231827 171866
rect 228968 171808 231766 171864
rect 231822 171808 231827 171864
rect 228968 171806 231827 171808
rect 231761 171803 231827 171806
rect 265617 171594 265683 171597
rect 268150 171594 268210 171836
rect 281574 171730 281580 171732
rect 279956 171670 281580 171730
rect 281574 171668 281580 171670
rect 281644 171668 281650 171732
rect 265617 171592 268210 171594
rect 164694 171534 167611 171536
rect 167545 171531 167611 171534
rect 265617 171536 265622 171592
rect 265678 171536 268210 171592
rect 265617 171534 268210 171536
rect 265617 171531 265683 171534
rect 229277 171458 229343 171461
rect 228968 171456 229343 171458
rect 228968 171400 229282 171456
rect 229338 171400 229343 171456
rect 228968 171398 229343 171400
rect 229277 171395 229343 171398
rect 215109 171186 215175 171189
rect 265801 171186 265867 171189
rect 268334 171186 268394 171428
rect 215109 171184 217242 171186
rect 215109 171128 215114 171184
rect 215170 171128 217242 171184
rect 215109 171126 217242 171128
rect 215109 171123 215175 171126
rect 217182 171020 217242 171126
rect 265801 171184 268394 171186
rect 265801 171128 265806 171184
rect 265862 171128 268394 171184
rect 265801 171126 268394 171128
rect 265801 171123 265867 171126
rect 231761 170914 231827 170917
rect 228968 170912 231827 170914
rect 228968 170856 231766 170912
rect 231822 170856 231827 170912
rect 228968 170854 231827 170856
rect 231761 170851 231827 170854
rect 214005 170778 214071 170781
rect 214005 170776 217242 170778
rect 214005 170720 214010 170776
rect 214066 170720 217242 170776
rect 214005 170718 217242 170720
rect 214005 170715 214071 170718
rect 217182 170340 217242 170718
rect 265433 170642 265499 170645
rect 268150 170642 268210 171020
rect 282269 170914 282335 170917
rect 279956 170912 282335 170914
rect 279956 170856 282274 170912
rect 282330 170856 282335 170912
rect 279956 170854 282335 170856
rect 282269 170851 282335 170854
rect 265433 170640 268210 170642
rect 265433 170584 265438 170640
rect 265494 170584 268210 170640
rect 265433 170582 268210 170584
rect 265433 170579 265499 170582
rect 231117 170506 231183 170509
rect 228968 170504 231183 170506
rect 228968 170448 231122 170504
rect 231178 170448 231183 170504
rect 228968 170446 231183 170448
rect 231117 170443 231183 170446
rect 265249 170234 265315 170237
rect 268150 170234 268210 170476
rect 265249 170232 268210 170234
rect 265249 170176 265254 170232
rect 265310 170176 268210 170232
rect 265249 170174 268210 170176
rect 265249 170171 265315 170174
rect 281625 170098 281691 170101
rect 279956 170096 281691 170098
rect 231485 169962 231551 169965
rect 228968 169960 231551 169962
rect 228968 169904 231490 169960
rect 231546 169904 231551 169960
rect 228968 169902 231551 169904
rect 231485 169899 231551 169902
rect 265617 169826 265683 169829
rect 268150 169826 268210 170068
rect 279956 170040 281630 170096
rect 281686 170040 281691 170096
rect 279956 170038 281691 170040
rect 281625 170035 281691 170038
rect 216998 169766 217242 169826
rect 214005 169690 214071 169693
rect 216998 169690 217058 169766
rect 214005 169688 217058 169690
rect 214005 169632 214010 169688
rect 214066 169632 217058 169688
rect 217182 169660 217242 169766
rect 265617 169824 268210 169826
rect 265617 169768 265622 169824
rect 265678 169768 268210 169824
rect 265617 169766 268210 169768
rect 265617 169763 265683 169766
rect 214005 169630 217058 169632
rect 214005 169627 214071 169630
rect 230749 169554 230815 169557
rect 228968 169552 230815 169554
rect 228968 169496 230754 169552
rect 230810 169496 230815 169552
rect 228968 169494 230815 169496
rect 230749 169491 230815 169494
rect 213913 169418 213979 169421
rect 265801 169418 265867 169421
rect 268150 169418 268210 169660
rect 280429 169418 280495 169421
rect 213913 169416 217242 169418
rect 213913 169360 213918 169416
rect 213974 169360 217242 169416
rect 213913 169358 217242 169360
rect 213913 169355 213979 169358
rect 217182 168980 217242 169358
rect 265801 169416 268210 169418
rect 265801 169360 265806 169416
rect 265862 169360 268210 169416
rect 265801 169358 268210 169360
rect 279956 169416 280495 169418
rect 279956 169360 280434 169416
rect 280490 169360 280495 169416
rect 279956 169358 280495 169360
rect 265801 169355 265867 169358
rect 280429 169355 280495 169358
rect 231485 169010 231551 169013
rect 228968 169008 231551 169010
rect 228968 168952 231490 169008
rect 231546 168952 231551 169008
rect 228968 168950 231551 168952
rect 231485 168947 231551 168950
rect 265341 169010 265407 169013
rect 268150 169010 268210 169252
rect 265341 169008 268210 169010
rect 265341 168952 265346 169008
rect 265402 168952 268210 169008
rect 265341 168950 268210 168952
rect 265341 168947 265407 168950
rect 229369 168602 229435 168605
rect 228968 168600 229435 168602
rect 228968 168544 229374 168600
rect 229430 168544 229435 168600
rect 228968 168542 229435 168544
rect 229369 168539 229435 168542
rect 265617 168602 265683 168605
rect 268150 168602 268210 168844
rect 282821 168602 282887 168605
rect 265617 168600 268210 168602
rect 265617 168544 265622 168600
rect 265678 168544 268210 168600
rect 265617 168542 268210 168544
rect 279956 168600 282887 168602
rect 279956 168544 282826 168600
rect 282882 168544 282887 168600
rect 279956 168542 282887 168544
rect 265617 168539 265683 168542
rect 282821 168539 282887 168542
rect 168414 168404 168420 168468
rect 168484 168466 168490 168468
rect 169661 168466 169727 168469
rect 265249 168466 265315 168469
rect 168484 168464 169727 168466
rect 168484 168408 169666 168464
rect 169722 168408 169727 168464
rect 168484 168406 169727 168408
rect 168484 168404 168490 168406
rect 169661 168403 169727 168406
rect 216998 168406 217242 168466
rect 213913 168330 213979 168333
rect 216998 168330 217058 168406
rect 213913 168328 217058 168330
rect 213913 168272 213918 168328
rect 213974 168272 217058 168328
rect 217182 168300 217242 168406
rect 265249 168464 267842 168466
rect 265249 168408 265254 168464
rect 265310 168408 267842 168464
rect 265249 168406 267842 168408
rect 265249 168403 265315 168406
rect 238753 168332 238819 168333
rect 213913 168270 217058 168272
rect 213913 168267 213979 168270
rect 238702 168268 238708 168332
rect 238772 168330 238819 168332
rect 238772 168328 238864 168330
rect 238814 168272 238864 168328
rect 238772 168270 238864 168272
rect 238772 168268 238819 168270
rect 238753 168267 238819 168268
rect 267782 168194 267842 168406
rect 268334 168194 268394 168436
rect 267782 168134 268394 168194
rect 214005 168058 214071 168061
rect 231761 168058 231827 168061
rect 214005 168056 217242 168058
rect 214005 168000 214010 168056
rect 214066 168000 217242 168056
rect 214005 167998 217242 168000
rect 228968 168056 231827 168058
rect 228968 168000 231766 168056
rect 231822 168000 231827 168056
rect 228968 167998 231827 168000
rect 214005 167995 214071 167998
rect 217182 167620 217242 167998
rect 231761 167995 231827 167998
rect 237598 167650 237604 167652
rect 228968 167590 237604 167650
rect 237598 167588 237604 167590
rect 237668 167588 237674 167652
rect 265341 167650 265407 167653
rect 268150 167650 268210 167892
rect 281717 167786 281783 167789
rect 279956 167784 281783 167786
rect 279956 167728 281722 167784
rect 281778 167728 281783 167784
rect 279956 167726 281783 167728
rect 281717 167723 281783 167726
rect 265341 167648 268210 167650
rect 265341 167592 265346 167648
rect 265402 167592 268210 167648
rect 265341 167590 268210 167592
rect 265341 167587 265407 167590
rect 268518 167244 268578 167484
rect 258030 167182 268210 167242
rect 231761 167106 231827 167109
rect 228968 167104 231827 167106
rect 228968 167048 231766 167104
rect 231822 167048 231827 167104
rect 228968 167046 231827 167048
rect 231761 167043 231827 167046
rect 239070 167044 239076 167108
rect 239140 167106 239146 167108
rect 258030 167106 258090 167182
rect 239140 167046 258090 167106
rect 268150 167076 268210 167182
rect 268510 167180 268516 167244
rect 268580 167180 268586 167244
rect 282453 167106 282519 167109
rect 279956 167104 282519 167106
rect 279956 167048 282458 167104
rect 282514 167048 282519 167104
rect 279956 167046 282519 167048
rect 239140 167044 239146 167046
rect 282453 167043 282519 167046
rect 213913 166970 213979 166973
rect 216998 166970 217242 167010
rect 213913 166968 217242 166970
rect 213913 166912 213918 166968
rect 213974 166950 217242 166968
rect 213974 166912 217058 166950
rect 217182 166940 217242 166950
rect 213913 166910 217058 166912
rect 213913 166907 213979 166910
rect 264421 166834 264487 166837
rect 268510 166834 268516 166836
rect 264421 166832 268516 166834
rect 264421 166776 264426 166832
rect 264482 166776 268516 166832
rect 264421 166774 268516 166776
rect 264421 166771 264487 166774
rect 268510 166772 268516 166774
rect 268580 166772 268586 166836
rect 214005 166698 214071 166701
rect 232037 166698 232103 166701
rect 214005 166696 217242 166698
rect 214005 166640 214010 166696
rect 214066 166640 217242 166696
rect 214005 166638 217242 166640
rect 228968 166696 232103 166698
rect 228968 166640 232042 166696
rect 232098 166640 232103 166696
rect 228968 166638 232103 166640
rect 214005 166635 214071 166638
rect 217182 166396 217242 166638
rect 232037 166635 232103 166638
rect 265709 166426 265775 166429
rect 268150 166426 268210 166668
rect 265709 166424 268210 166426
rect 265709 166368 265714 166424
rect 265770 166368 268210 166424
rect 265709 166366 268210 166368
rect 265709 166363 265775 166366
rect 282085 166290 282151 166293
rect 279956 166288 282151 166290
rect 213269 166154 213335 166157
rect 231669 166154 231735 166157
rect 213269 166152 217242 166154
rect 213269 166096 213274 166152
rect 213330 166096 217242 166152
rect 213269 166094 217242 166096
rect 228968 166152 231735 166154
rect 228968 166096 231674 166152
rect 231730 166096 231735 166152
rect 228968 166094 231735 166096
rect 213269 166091 213335 166094
rect 217182 165716 217242 166094
rect 231669 166091 231735 166094
rect 265341 166018 265407 166021
rect 268150 166018 268210 166260
rect 279956 166232 282090 166288
rect 282146 166232 282151 166288
rect 279956 166230 282151 166232
rect 282085 166227 282151 166230
rect 265341 166016 268210 166018
rect 265341 165960 265346 166016
rect 265402 165960 268210 166016
rect 265341 165958 268210 165960
rect 265341 165955 265407 165958
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 231761 165746 231827 165749
rect 228968 165744 231827 165746
rect 228968 165688 231766 165744
rect 231822 165688 231827 165744
rect 228968 165686 231827 165688
rect 231761 165683 231827 165686
rect 265801 165746 265867 165749
rect 265801 165744 267842 165746
rect 265801 165688 265806 165744
rect 265862 165688 267842 165744
rect 265801 165686 267842 165688
rect 265801 165683 265867 165686
rect 267782 165610 267842 165686
rect 268334 165610 268394 165852
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 267782 165550 268394 165610
rect 280337 165474 280403 165477
rect 279956 165472 280403 165474
rect 279956 165416 280342 165472
rect 280398 165416 280403 165472
rect 279956 165414 280403 165416
rect 280337 165411 280403 165414
rect 213913 165338 213979 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 231761 165202 231827 165205
rect 228968 165200 231827 165202
rect 228968 165144 231766 165200
rect 231822 165144 231827 165200
rect 228968 165142 231827 165144
rect 231761 165139 231827 165142
rect 265341 165066 265407 165069
rect 268150 165066 268210 165308
rect 265341 165064 268210 165066
rect 265341 165008 265346 165064
rect 265402 165008 268210 165064
rect 265341 165006 268210 165008
rect 265341 165003 265407 165006
rect 213453 164794 213519 164797
rect 231669 164794 231735 164797
rect 213453 164792 217242 164794
rect 213453 164736 213458 164792
rect 213514 164736 217242 164792
rect 213453 164734 217242 164736
rect 228968 164792 231735 164794
rect 228968 164736 231674 164792
rect 231730 164736 231735 164792
rect 228968 164734 231735 164736
rect 213453 164731 213519 164734
rect 217182 164356 217242 164734
rect 231669 164731 231735 164734
rect 265157 164658 265223 164661
rect 268150 164658 268210 164900
rect 282085 164794 282151 164797
rect 279956 164792 282151 164794
rect 279956 164736 282090 164792
rect 282146 164736 282151 164792
rect 279956 164734 282151 164736
rect 282085 164731 282151 164734
rect 265157 164656 268210 164658
rect 265157 164600 265162 164656
rect 265218 164600 268210 164656
rect 265157 164598 268210 164600
rect 265157 164595 265223 164598
rect 231117 164386 231183 164389
rect 228968 164384 231183 164386
rect 228968 164328 231122 164384
rect 231178 164328 231183 164384
rect 228968 164326 231183 164328
rect 231117 164323 231183 164326
rect 265157 164250 265223 164253
rect 268150 164250 268210 164492
rect 265157 164248 268210 164250
rect 265157 164192 265162 164248
rect 265218 164192 268210 164248
rect 265157 164190 268210 164192
rect 265157 164187 265223 164190
rect 213913 163978 213979 163981
rect 213913 163976 217242 163978
rect 213913 163920 213918 163976
rect 213974 163920 217242 163976
rect 213913 163918 217242 163920
rect 213913 163915 213979 163918
rect 217182 163676 217242 163918
rect 231761 163842 231827 163845
rect 228968 163840 231827 163842
rect 228968 163784 231766 163840
rect 231822 163784 231827 163840
rect 228968 163782 231827 163784
rect 231761 163779 231827 163782
rect 264237 163842 264303 163845
rect 268150 163842 268210 164084
rect 282637 163978 282703 163981
rect 279956 163976 282703 163978
rect 279956 163920 282642 163976
rect 282698 163920 282703 163976
rect 279956 163918 282703 163920
rect 282637 163915 282703 163918
rect 264237 163840 268210 163842
rect 264237 163784 264242 163840
rect 264298 163784 268210 163840
rect 264237 163782 268210 163784
rect 264237 163779 264303 163782
rect 231669 163434 231735 163437
rect 228968 163432 231735 163434
rect 228968 163376 231674 163432
rect 231730 163376 231735 163432
rect 228968 163374 231735 163376
rect 231669 163371 231735 163374
rect 265801 163434 265867 163437
rect 268150 163434 268210 163676
rect 265801 163432 268210 163434
rect 265801 163376 265806 163432
rect 265862 163376 268210 163432
rect 265801 163374 268210 163376
rect 265801 163371 265867 163374
rect 200070 163102 217242 163162
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 166390 162828 166396 162892
rect 166460 162890 166466 162892
rect 200070 162890 200130 163102
rect 217182 162996 217242 163102
rect 265525 163026 265591 163029
rect 268518 163028 268578 163268
rect 282821 163162 282887 163165
rect 279956 163160 282887 163162
rect 279956 163104 282826 163160
rect 282882 163104 282887 163160
rect 279956 163102 282887 163104
rect 282821 163099 282887 163102
rect 265525 163024 268210 163026
rect 265525 162968 265530 163024
rect 265586 162968 268210 163024
rect 265525 162966 268210 162968
rect 265525 162963 265591 162966
rect 231117 162890 231183 162893
rect 166460 162830 200130 162890
rect 228968 162888 231183 162890
rect 228968 162832 231122 162888
rect 231178 162832 231183 162888
rect 268150 162860 268210 162966
rect 268510 162964 268516 163028
rect 268580 162964 268586 163028
rect 228968 162830 231183 162832
rect 166460 162828 166466 162830
rect 231117 162827 231183 162830
rect 213913 162618 213979 162621
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 231761 162482 231827 162485
rect 228968 162480 231827 162482
rect 228968 162424 231766 162480
rect 231822 162424 231827 162480
rect 228968 162422 231827 162424
rect 231761 162419 231827 162422
rect 264513 162482 264579 162485
rect 282821 162482 282887 162485
rect 264513 162480 268210 162482
rect 264513 162424 264518 162480
rect 264574 162424 268210 162480
rect 264513 162422 268210 162424
rect 279956 162480 282887 162482
rect 279956 162424 282826 162480
rect 282882 162424 282887 162480
rect 279956 162422 282887 162424
rect 264513 162419 264579 162422
rect 268150 162316 268210 162422
rect 282821 162419 282887 162422
rect 267966 162014 268210 162074
rect 231669 161938 231735 161941
rect 228968 161936 231735 161938
rect 228968 161880 231674 161936
rect 231730 161880 231735 161936
rect 228968 161878 231735 161880
rect 231669 161875 231735 161878
rect 264421 161938 264487 161941
rect 267966 161938 268026 162014
rect 264421 161936 268026 161938
rect 264421 161880 264426 161936
rect 264482 161880 268026 161936
rect 268150 161908 268210 162014
rect 264421 161878 268026 161880
rect 264421 161875 264487 161878
rect 166206 161604 166212 161668
rect 166276 161666 166282 161668
rect 166276 161606 200130 161666
rect 166276 161604 166282 161606
rect 200070 161530 200130 161606
rect 217366 161530 217426 161772
rect 265525 161666 265591 161669
rect 282545 161666 282611 161669
rect 265525 161664 268210 161666
rect 265525 161608 265530 161664
rect 265586 161608 268210 161664
rect 265525 161606 268210 161608
rect 279956 161664 282611 161666
rect 279956 161608 282550 161664
rect 282606 161608 282611 161664
rect 279956 161606 282611 161608
rect 265525 161603 265591 161606
rect 231025 161530 231091 161533
rect 200070 161470 217426 161530
rect 228968 161528 231091 161530
rect 228968 161472 231030 161528
rect 231086 161472 231091 161528
rect 268150 161500 268210 161606
rect 282545 161603 282611 161606
rect 228968 161470 231091 161472
rect 231025 161467 231091 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 231761 160986 231827 160989
rect 228968 160984 231827 160986
rect 228968 160928 231766 160984
rect 231822 160928 231827 160984
rect 228968 160926 231827 160928
rect 231761 160923 231827 160926
rect 214557 160850 214623 160853
rect 265985 160850 266051 160853
rect 268150 160850 268210 161092
rect 282821 160850 282887 160853
rect 214557 160848 217242 160850
rect 214557 160792 214562 160848
rect 214618 160792 217242 160848
rect 214557 160790 217242 160792
rect 214557 160787 214623 160790
rect 217182 160412 217242 160790
rect 265985 160848 268210 160850
rect 265985 160792 265990 160848
rect 266046 160792 268210 160848
rect 265985 160790 268210 160792
rect 279956 160848 282887 160850
rect 279956 160792 282826 160848
rect 282882 160792 282887 160848
rect 279956 160790 282887 160792
rect 265985 160787 266051 160790
rect 282821 160787 282887 160790
rect 231669 160578 231735 160581
rect 228968 160576 231735 160578
rect 228968 160520 231674 160576
rect 231730 160520 231735 160576
rect 228968 160518 231735 160520
rect 231669 160515 231735 160518
rect 265893 160442 265959 160445
rect 268150 160442 268210 160684
rect 265893 160440 268210 160442
rect 265893 160384 265898 160440
rect 265954 160384 268210 160440
rect 265893 160382 268210 160384
rect 265893 160379 265959 160382
rect 265801 160170 265867 160173
rect 265801 160168 267842 160170
rect 265801 160112 265806 160168
rect 265862 160112 267842 160168
rect 265801 160110 267842 160112
rect 265801 160107 265867 160110
rect 213913 160034 213979 160037
rect 231761 160034 231827 160037
rect 213913 160032 217242 160034
rect 213913 159976 213918 160032
rect 213974 159976 217242 160032
rect 213913 159974 217242 159976
rect 228968 160032 231827 160034
rect 228968 159976 231766 160032
rect 231822 159976 231827 160032
rect 228968 159974 231827 159976
rect 267782 160034 267842 160110
rect 268334 160034 268394 160276
rect 282361 160170 282427 160173
rect 279956 160168 282427 160170
rect 279956 160112 282366 160168
rect 282422 160112 282427 160168
rect 279956 160110 282427 160112
rect 282361 160107 282427 160110
rect 267782 159974 268394 160034
rect 213913 159971 213979 159974
rect 217182 159732 217242 159974
rect 231761 159971 231827 159974
rect 265617 159898 265683 159901
rect 268510 159898 268516 159900
rect 265617 159896 268516 159898
rect 265617 159840 265622 159896
rect 265678 159840 268516 159896
rect 265617 159838 268516 159840
rect 265617 159835 265683 159838
rect 268510 159836 268516 159838
rect 268580 159836 268586 159900
rect 231669 159626 231735 159629
rect 228968 159624 231735 159626
rect 228968 159568 231674 159624
rect 231730 159568 231735 159624
rect 228968 159566 231735 159568
rect 231669 159563 231735 159566
rect 214005 159490 214071 159493
rect 265525 159490 265591 159493
rect 268150 159490 268210 159732
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 265525 159488 268210 159490
rect 265525 159432 265530 159488
rect 265586 159432 268210 159488
rect 265525 159430 268210 159432
rect 265525 159427 265591 159430
rect 282729 159354 282795 159357
rect 279956 159352 282795 159354
rect 231669 159082 231735 159085
rect 228968 159080 231735 159082
rect 228968 159024 231674 159080
rect 231730 159024 231735 159080
rect 228968 159022 231735 159024
rect 231669 159019 231735 159022
rect 237966 159020 237972 159084
rect 238036 159082 238042 159084
rect 268150 159082 268210 159324
rect 279956 159296 282734 159352
rect 282790 159296 282795 159352
rect 279956 159294 282795 159296
rect 282729 159291 282795 159294
rect 238036 159022 268210 159082
rect 238036 159020 238042 159022
rect 231485 158810 231551 158813
rect 237414 158810 237420 158812
rect 231485 158808 237420 158810
rect 231485 158752 231490 158808
rect 231546 158752 237420 158808
rect 231485 158750 237420 158752
rect 231485 158747 231551 158750
rect 237414 158748 237420 158750
rect 237484 158748 237490 158812
rect 265801 158810 265867 158813
rect 265801 158808 267842 158810
rect 265801 158752 265806 158808
rect 265862 158752 267842 158808
rect 265801 158750 267842 158752
rect 265801 158747 265867 158750
rect 214097 158674 214163 158677
rect 230565 158674 230631 158677
rect 214097 158672 217242 158674
rect 214097 158616 214102 158672
rect 214158 158616 217242 158672
rect 214097 158614 217242 158616
rect 228968 158672 230631 158674
rect 228968 158616 230570 158672
rect 230626 158616 230631 158672
rect 228968 158614 230631 158616
rect 267782 158674 267842 158750
rect 268334 158674 268394 158916
rect 267782 158614 268394 158674
rect 214097 158611 214163 158614
rect 217182 158372 217242 158614
rect 230565 158611 230631 158614
rect 280153 158538 280219 158541
rect 279956 158536 280219 158538
rect 265985 158266 266051 158269
rect 268150 158266 268210 158508
rect 279956 158480 280158 158536
rect 280214 158480 280219 158536
rect 279956 158478 280219 158480
rect 280153 158475 280219 158478
rect 265985 158264 268210 158266
rect 265985 158208 265990 158264
rect 266046 158208 268210 158264
rect 265985 158206 268210 158208
rect 265985 158203 266051 158206
rect 215017 158130 215083 158133
rect 229502 158130 229508 158132
rect 215017 158128 217242 158130
rect 215017 158072 215022 158128
rect 215078 158072 217242 158128
rect 215017 158070 217242 158072
rect 228968 158070 229508 158130
rect 215017 158067 215083 158070
rect 217182 157692 217242 158070
rect 229502 158068 229508 158070
rect 229572 158068 229578 158132
rect 265801 157858 265867 157861
rect 268150 157858 268210 158100
rect 282269 157858 282335 157861
rect 265801 157856 268210 157858
rect 265801 157800 265806 157856
rect 265862 157800 268210 157856
rect 265801 157798 268210 157800
rect 279956 157856 282335 157858
rect 279956 157800 282274 157856
rect 282330 157800 282335 157856
rect 279956 157798 282335 157800
rect 265801 157795 265867 157798
rect 282269 157795 282335 157798
rect 230473 157722 230539 157725
rect 228968 157720 230539 157722
rect 228968 157664 230478 157720
rect 230534 157664 230539 157720
rect 228968 157662 230539 157664
rect 230473 157659 230539 157662
rect 265065 157450 265131 157453
rect 268334 157450 268394 157692
rect 265065 157448 268394 157450
rect 265065 157392 265070 157448
rect 265126 157392 268394 157448
rect 265065 157390 268394 157392
rect 265065 157387 265131 157390
rect 213913 157314 213979 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 231761 157178 231827 157181
rect 228968 157176 231827 157178
rect 228968 157120 231766 157176
rect 231822 157120 231827 157176
rect 228968 157118 231827 157120
rect 231761 157115 231827 157118
rect 214005 156906 214071 156909
rect 265893 156906 265959 156909
rect 268150 156906 268210 157148
rect 282821 157042 282887 157045
rect 279956 157040 282887 157042
rect 279956 156984 282826 157040
rect 282882 156984 282887 157040
rect 279956 156982 282887 156984
rect 282821 156979 282887 156982
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 265893 156904 268210 156906
rect 265893 156848 265898 156904
rect 265954 156848 268210 156904
rect 265893 156846 268210 156848
rect 265893 156843 265959 156846
rect 231669 156770 231735 156773
rect 228968 156768 231735 156770
rect 228968 156712 231674 156768
rect 231730 156712 231735 156768
rect 228968 156710 231735 156712
rect 231669 156707 231735 156710
rect 266077 156498 266143 156501
rect 268150 156498 268210 156740
rect 279366 156708 279372 156772
rect 279436 156708 279442 156772
rect 266077 156496 268210 156498
rect 266077 156440 266082 156496
rect 266138 156440 268210 156496
rect 266077 156438 268210 156440
rect 266077 156435 266143 156438
rect 279374 156332 279434 156708
rect 230933 156226 230999 156229
rect 228968 156224 230999 156226
rect 228968 156168 230938 156224
rect 230994 156168 230999 156224
rect 228968 156166 230999 156168
rect 230933 156163 230999 156166
rect 265801 156090 265867 156093
rect 268150 156090 268210 156332
rect 265801 156088 268210 156090
rect 265801 156032 265806 156088
rect 265862 156032 268210 156088
rect 265801 156030 268210 156032
rect 265801 156027 265867 156030
rect 214833 155954 214899 155957
rect 214833 155952 217242 155954
rect 214833 155896 214838 155952
rect 214894 155896 217242 155952
rect 214833 155894 217242 155896
rect 214833 155891 214899 155894
rect 217182 155788 217242 155894
rect 230565 155818 230631 155821
rect 228968 155816 230631 155818
rect 228968 155760 230570 155816
rect 230626 155760 230631 155816
rect 228968 155758 230631 155760
rect 230565 155755 230631 155758
rect 265709 155682 265775 155685
rect 268150 155682 268210 155924
rect 265709 155680 268210 155682
rect 265709 155624 265714 155680
rect 265770 155624 268210 155680
rect 265709 155622 268210 155624
rect 265709 155619 265775 155622
rect 213913 155546 213979 155549
rect 282821 155546 282887 155549
rect 213913 155544 217242 155546
rect 213913 155488 213918 155544
rect 213974 155488 217242 155544
rect 279956 155544 282887 155546
rect 213913 155486 217242 155488
rect 213913 155483 213979 155486
rect 217182 155108 217242 155486
rect 230933 155274 230999 155277
rect 228968 155272 230999 155274
rect 228968 155216 230938 155272
rect 230994 155216 230999 155272
rect 228968 155214 230999 155216
rect 230933 155211 230999 155214
rect 265985 155274 266051 155277
rect 268150 155274 268210 155516
rect 279956 155488 282826 155544
rect 282882 155488 282887 155544
rect 279956 155486 282887 155488
rect 282821 155483 282887 155486
rect 265985 155272 268210 155274
rect 265985 155216 265990 155272
rect 266046 155216 268210 155272
rect 265985 155214 268210 155216
rect 265985 155211 266051 155214
rect 247718 154866 247724 154868
rect 228968 154806 247724 154866
rect 247718 154804 247724 154806
rect 247788 154804 247794 154868
rect 265801 154866 265867 154869
rect 268150 154866 268210 155108
rect 265801 154864 268210 154866
rect 265801 154808 265806 154864
rect 265862 154808 268210 154864
rect 265801 154806 268210 154808
rect 265801 154803 265867 154806
rect 265893 154730 265959 154733
rect 281533 154730 281599 154733
rect 265893 154728 268210 154730
rect 265893 154672 265898 154728
rect 265954 154672 268210 154728
rect 265893 154670 268210 154672
rect 279956 154728 281599 154730
rect 279956 154672 281538 154728
rect 281594 154672 281599 154728
rect 279956 154670 281599 154672
rect 265893 154667 265959 154670
rect 268150 154564 268210 154670
rect 281533 154667 281599 154670
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 231761 154322 231827 154325
rect 228968 154320 231827 154322
rect 228968 154264 231766 154320
rect 231822 154264 231827 154320
rect 228968 154262 231827 154264
rect 231761 154259 231827 154262
rect 231393 153914 231459 153917
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 228968 153912 231459 153914
rect 228968 153856 231398 153912
rect 231454 153856 231459 153912
rect 228968 153854 231459 153856
rect 214005 153851 214071 153854
rect 231393 153851 231459 153854
rect 265341 153914 265407 153917
rect 268150 153914 268210 154156
rect 281901 154050 281967 154053
rect 279956 154048 281967 154050
rect 279956 153992 281906 154048
rect 281962 153992 281967 154048
rect 279956 153990 281967 153992
rect 281901 153987 281967 153990
rect 265341 153912 268210 153914
rect 265341 153856 265346 153912
rect 265402 153856 268210 153912
rect 265341 153854 268210 153856
rect 265341 153851 265407 153854
rect 213913 153370 213979 153373
rect 217182 153370 217242 153748
rect 265801 153506 265867 153509
rect 268150 153506 268210 153748
rect 265801 153504 268210 153506
rect 265801 153448 265806 153504
rect 265862 153448 268210 153504
rect 265801 153446 268210 153448
rect 265801 153443 265867 153446
rect 231301 153370 231367 153373
rect 213913 153368 217242 153370
rect 213913 153312 213918 153368
rect 213974 153312 217242 153368
rect 213913 153310 217242 153312
rect 228968 153368 231367 153370
rect 228968 153312 231306 153368
rect 231362 153312 231367 153368
rect 228968 153310 231367 153312
rect 213913 153307 213979 153310
rect 231301 153307 231367 153310
rect 232681 153234 232747 153237
rect 240542 153234 240548 153236
rect 232681 153232 240548 153234
rect 232681 153176 232686 153232
rect 232742 153176 240548 153232
rect 232681 153174 240548 153176
rect 232681 153171 232747 153174
rect 240542 153172 240548 153174
rect 240612 153172 240618 153236
rect 265893 153234 265959 153237
rect 265893 153232 267842 153234
rect 265893 153176 265898 153232
rect 265954 153176 267842 153232
rect 265893 153174 267842 153176
rect 265893 153171 265959 153174
rect 267782 153098 267842 153174
rect 268334 153098 268394 153340
rect 281717 153234 281783 153237
rect 279956 153232 281783 153234
rect 279956 153176 281722 153232
rect 281778 153176 281783 153232
rect 279956 153174 281783 153176
rect 281717 153171 281783 153174
rect 213913 152690 213979 152693
rect 217182 152690 217242 153068
rect 267782 153038 268394 153098
rect 230749 152962 230815 152965
rect 228968 152960 230815 152962
rect 228968 152904 230754 152960
rect 230810 152904 230815 152960
rect 228968 152902 230815 152904
rect 230749 152899 230815 152902
rect 213913 152688 217242 152690
rect 213913 152632 213918 152688
rect 213974 152632 217242 152688
rect 213913 152630 217242 152632
rect 264329 152690 264395 152693
rect 268150 152690 268210 152932
rect 264329 152688 268210 152690
rect 264329 152632 264334 152688
rect 264390 152632 268210 152688
rect 264329 152630 268210 152632
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 213913 152627 213979 152630
rect 264329 152627 264395 152630
rect 579797 152627 579863 152630
rect 231669 152554 231735 152557
rect 228968 152552 231735 152554
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 228968 152496 231674 152552
rect 231730 152496 231735 152552
rect 583520 152540 584960 152630
rect 228968 152494 231735 152496
rect 231669 152491 231735 152494
rect 240726 152356 240732 152420
rect 240796 152418 240802 152420
rect 266077 152418 266143 152421
rect 240796 152416 266143 152418
rect 240796 152360 266082 152416
rect 266138 152360 266143 152416
rect 240796 152358 266143 152360
rect 240796 152356 240802 152358
rect 266077 152355 266143 152358
rect 265249 152146 265315 152149
rect 268150 152146 268210 152524
rect 282177 152418 282243 152421
rect 279956 152416 282243 152418
rect 279956 152360 282182 152416
rect 282238 152360 282243 152416
rect 279956 152358 282243 152360
rect 282177 152355 282243 152358
rect 265249 152144 268210 152146
rect 265249 152088 265254 152144
rect 265310 152088 268210 152144
rect 265249 152086 268210 152088
rect 265249 152083 265315 152086
rect 231761 152010 231827 152013
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 228968 152008 231827 152010
rect 228968 151952 231766 152008
rect 231822 151952 231827 152008
rect 228968 151950 231827 151952
rect 213913 151947 213979 151950
rect 231761 151947 231827 151950
rect 214649 151874 214715 151877
rect 265801 151874 265867 151877
rect 214649 151872 217058 151874
rect 214649 151816 214654 151872
rect 214710 151830 217058 151872
rect 265801 151872 267842 151874
rect 217182 151830 217242 151844
rect 214710 151816 217242 151830
rect 214649 151814 217242 151816
rect 214649 151811 214715 151814
rect 216998 151770 217242 151814
rect 265801 151816 265806 151872
rect 265862 151816 267842 151872
rect 265801 151814 267842 151816
rect 265801 151811 265867 151814
rect 267782 151738 267842 151814
rect 268334 151738 268394 151980
rect 282821 151738 282887 151741
rect 267782 151678 268394 151738
rect 279956 151736 282887 151738
rect 279956 151680 282826 151736
rect 282882 151680 282887 151736
rect 279956 151678 282887 151680
rect 282821 151675 282887 151678
rect 231761 151602 231827 151605
rect 228968 151600 231827 151602
rect 228968 151544 231766 151600
rect 231822 151544 231827 151600
rect 228968 151542 231827 151544
rect 231761 151539 231827 151542
rect 265709 151330 265775 151333
rect 268150 151330 268210 151572
rect 265709 151328 268210 151330
rect 265709 151272 265714 151328
rect 265770 151272 268210 151328
rect 265709 151270 268210 151272
rect 265709 151267 265775 151270
rect 213913 150922 213979 150925
rect 217182 150922 217242 151164
rect 229829 151058 229895 151061
rect 228968 151056 229895 151058
rect 228968 151000 229834 151056
rect 229890 151000 229895 151056
rect 228968 150998 229895 151000
rect 229829 150995 229895 150998
rect 213913 150920 217242 150922
rect 213913 150864 213918 150920
rect 213974 150864 217242 150920
rect 213913 150862 217242 150864
rect 265433 150922 265499 150925
rect 268150 150922 268210 151164
rect 281993 150922 282059 150925
rect 265433 150920 268210 150922
rect 265433 150864 265438 150920
rect 265494 150864 268210 150920
rect 265433 150862 268210 150864
rect 279956 150920 282059 150922
rect 279956 150864 281998 150920
rect 282054 150864 282059 150920
rect 279956 150862 282059 150864
rect 213913 150859 213979 150862
rect 265433 150859 265499 150862
rect 281993 150859 282059 150862
rect 214465 150786 214531 150789
rect 214465 150784 217426 150786
rect 214465 150728 214470 150784
rect 214526 150728 217426 150784
rect 214465 150726 217426 150728
rect 214465 150723 214531 150726
rect 217366 150484 217426 150726
rect 231669 150650 231735 150653
rect 228968 150648 231735 150650
rect 228968 150592 231674 150648
rect 231730 150592 231735 150648
rect 228968 150590 231735 150592
rect 231669 150587 231735 150590
rect 265801 150514 265867 150517
rect 268334 150514 268394 150756
rect 265801 150512 268394 150514
rect 265801 150456 265806 150512
rect 265862 150456 268394 150512
rect 265801 150454 268394 150456
rect 265801 150451 265867 150454
rect 214005 150242 214071 150245
rect 214005 150240 217242 150242
rect 214005 150184 214010 150240
rect 214066 150184 217242 150240
rect 214005 150182 217242 150184
rect 214005 150179 214071 150182
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150182
rect 230933 150106 230999 150109
rect 228968 150104 230999 150106
rect 228968 150048 230938 150104
rect 230994 150048 230999 150104
rect 228968 150046 230999 150048
rect 230933 150043 230999 150046
rect 265801 150106 265867 150109
rect 268150 150106 268210 150348
rect 282821 150106 282887 150109
rect 265801 150104 268210 150106
rect 265801 150048 265806 150104
rect 265862 150048 268210 150104
rect 265801 150046 268210 150048
rect 279956 150104 282887 150106
rect 279956 150048 282826 150104
rect 282882 150048 282887 150104
rect 279956 150046 282887 150048
rect 265801 150043 265867 150046
rect 282821 150043 282887 150046
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 231025 149698 231091 149701
rect 228968 149696 231091 149698
rect 228968 149640 231030 149696
rect 231086 149640 231091 149696
rect 228968 149638 231091 149640
rect 231025 149635 231091 149638
rect 265341 149698 265407 149701
rect 268150 149698 268210 149940
rect 265341 149696 268210 149698
rect 265341 149640 265346 149696
rect 265402 149640 268210 149696
rect 265341 149638 268210 149640
rect 265341 149635 265407 149638
rect 214925 149562 214991 149565
rect 214925 149560 217242 149562
rect 214925 149504 214930 149560
rect 214986 149504 217242 149560
rect 214925 149502 217242 149504
rect 214925 149499 214991 149502
rect 217182 149124 217242 149502
rect 231301 149154 231367 149157
rect 228968 149152 231367 149154
rect 228968 149096 231306 149152
rect 231362 149096 231367 149152
rect 228968 149094 231367 149096
rect 231301 149091 231367 149094
rect 265433 149154 265499 149157
rect 268150 149154 268210 149532
rect 282177 149426 282243 149429
rect 279956 149424 282243 149426
rect 279956 149368 282182 149424
rect 282238 149368 282243 149424
rect 279956 149366 282243 149368
rect 282177 149363 282243 149366
rect 265433 149152 268210 149154
rect 265433 149096 265438 149152
rect 265494 149096 268210 149152
rect 265433 149094 268210 149096
rect 265433 149091 265499 149094
rect 213913 148746 213979 148749
rect 233182 148746 233188 148748
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 228968 148686 233188 148746
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 233182 148684 233188 148686
rect 233252 148684 233258 148748
rect 265525 148746 265591 148749
rect 268150 148746 268210 148988
rect 265525 148744 268210 148746
rect 265525 148688 265530 148744
rect 265586 148688 268210 148744
rect 265525 148686 268210 148688
rect 265525 148683 265591 148686
rect 282085 148610 282151 148613
rect 279956 148608 282151 148610
rect 265709 148338 265775 148341
rect 268150 148338 268210 148580
rect 279956 148552 282090 148608
rect 282146 148552 282151 148608
rect 279956 148550 282151 148552
rect 282085 148547 282151 148550
rect 265709 148336 268210 148338
rect 265709 148280 265714 148336
rect 265770 148280 268210 148336
rect 265709 148278 268210 148280
rect 265709 148275 265775 148278
rect 231761 148202 231827 148205
rect 228968 148200 231827 148202
rect 228968 148144 231766 148200
rect 231822 148144 231827 148200
rect 228968 148142 231827 148144
rect 231761 148139 231827 148142
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 265065 147930 265131 147933
rect 268518 147932 268578 148172
rect 265065 147928 268210 147930
rect 265065 147872 265070 147928
rect 265126 147872 268210 147928
rect 265065 147870 268210 147872
rect 265065 147867 265131 147870
rect 230422 147794 230428 147796
rect 228968 147734 230428 147794
rect 230422 147732 230428 147734
rect 230492 147732 230498 147796
rect 268150 147764 268210 147870
rect 268510 147868 268516 147932
rect 268580 147868 268586 147932
rect 283005 147794 283071 147797
rect 279956 147792 283071 147794
rect 279956 147736 283010 147792
rect 283066 147736 283071 147792
rect 279956 147734 283071 147736
rect 283005 147731 283071 147734
rect 230749 147250 230815 147253
rect 228968 147248 230815 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 228968 147192 230754 147248
rect 230810 147192 230815 147248
rect 228968 147190 230815 147192
rect 230749 147187 230815 147190
rect 265893 147114 265959 147117
rect 268150 147114 268210 147356
rect 281717 147114 281783 147117
rect 265893 147112 268210 147114
rect 265893 147056 265898 147112
rect 265954 147056 268210 147112
rect 265893 147054 268210 147056
rect 279956 147112 281783 147114
rect 279956 147056 281722 147112
rect 281778 147056 281783 147112
rect 279956 147054 281783 147056
rect 265893 147051 265959 147054
rect 281717 147051 281783 147054
rect 230933 146842 230999 146845
rect 228968 146840 230999 146842
rect 228968 146784 230938 146840
rect 230994 146784 230999 146840
rect 228968 146782 230999 146784
rect 230933 146779 230999 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 265525 146706 265591 146709
rect 268150 146706 268210 146948
rect 265525 146704 268210 146706
rect 265525 146648 265530 146704
rect 265586 146648 268210 146704
rect 265525 146646 268210 146648
rect 214005 146643 214071 146646
rect 265525 146643 265591 146646
rect 265985 146570 266051 146573
rect 265985 146568 268210 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 265985 146512 265990 146568
rect 266046 146512 268210 146568
rect 265985 146510 268210 146512
rect 265985 146507 266051 146510
rect 268150 146404 268210 146510
rect 231485 146298 231551 146301
rect 282821 146298 282887 146301
rect 216814 146238 217426 146298
rect 228968 146296 231551 146298
rect 228968 146240 231490 146296
rect 231546 146240 231551 146296
rect 228968 146238 231551 146240
rect 279956 146296 282887 146298
rect 279956 146240 282826 146296
rect 282882 146240 282887 146296
rect 279956 146238 282887 146240
rect 231485 146235 231551 146238
rect 282821 146235 282887 146238
rect 230974 146100 230980 146164
rect 231044 146162 231050 146164
rect 238293 146162 238359 146165
rect 231044 146160 238359 146162
rect 231044 146104 238298 146160
rect 238354 146104 238359 146160
rect 231044 146102 238359 146104
rect 231044 146100 231050 146102
rect 238293 146099 238359 146102
rect 265433 146162 265499 146165
rect 268510 146162 268516 146164
rect 265433 146160 268516 146162
rect 265433 146104 265438 146160
rect 265494 146104 268516 146160
rect 265433 146102 268516 146104
rect 265433 146099 265499 146102
rect 268510 146100 268516 146102
rect 268580 146100 268586 146164
rect 231761 145890 231827 145893
rect 228968 145888 231827 145890
rect 217182 145346 217242 145860
rect 228968 145832 231766 145888
rect 231822 145832 231827 145888
rect 228968 145830 231827 145832
rect 231761 145827 231827 145830
rect 265801 145754 265867 145757
rect 268150 145754 268210 145996
rect 265801 145752 268210 145754
rect 265801 145696 265806 145752
rect 265862 145696 268210 145752
rect 265801 145694 268210 145696
rect 265801 145691 265867 145694
rect 231669 145346 231735 145349
rect 200070 145286 217242 145346
rect 228968 145344 231735 145346
rect 228968 145288 231674 145344
rect 231730 145288 231735 145344
rect 228968 145286 231735 145288
rect 166206 144876 166212 144940
rect 166276 144938 166282 144940
rect 200070 144938 200130 145286
rect 231669 145283 231735 145286
rect 265709 145346 265775 145349
rect 268150 145346 268210 145588
rect 282729 145482 282795 145485
rect 279956 145480 282795 145482
rect 279956 145424 282734 145480
rect 282790 145424 282795 145480
rect 279956 145422 282795 145424
rect 282729 145419 282795 145422
rect 265709 145344 268210 145346
rect 265709 145288 265714 145344
rect 265770 145288 268210 145344
rect 265709 145286 268210 145288
rect 265709 145283 265775 145286
rect 166276 144878 200130 144938
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 231669 144938 231735 144941
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 228968 144936 231735 144938
rect 228968 144880 231674 144936
rect 231730 144880 231735 144936
rect 228968 144878 231735 144880
rect 166276 144876 166282 144878
rect 213913 144875 213979 144878
rect 231669 144875 231735 144878
rect 265893 144938 265959 144941
rect 268334 144938 268394 145180
rect 265893 144936 268394 144938
rect 265893 144880 265898 144936
rect 265954 144880 268394 144936
rect 265893 144878 268394 144880
rect 265893 144875 265959 144878
rect 282821 144802 282887 144805
rect 279956 144800 282887 144802
rect 265525 144530 265591 144533
rect 268150 144530 268210 144772
rect 279956 144744 282826 144800
rect 282882 144744 282887 144800
rect 279956 144742 282887 144744
rect 282821 144739 282887 144742
rect 265525 144528 268210 144530
rect 213913 143986 213979 143989
rect 217182 143986 217242 144500
rect 265525 144472 265530 144528
rect 265586 144472 268210 144528
rect 265525 144470 268210 144472
rect 265525 144467 265591 144470
rect 231761 144394 231827 144397
rect 228968 144392 231827 144394
rect 228968 144336 231766 144392
rect 231822 144336 231827 144392
rect 228968 144334 231827 144336
rect 231761 144331 231827 144334
rect 230749 143986 230815 143989
rect 213913 143984 217242 143986
rect 213913 143928 213918 143984
rect 213974 143928 217242 143984
rect 213913 143926 217242 143928
rect 228968 143984 230815 143986
rect 228968 143928 230754 143984
rect 230810 143928 230815 143984
rect 228968 143926 230815 143928
rect 213913 143923 213979 143926
rect 230749 143923 230815 143926
rect 233734 143924 233740 143988
rect 233804 143986 233810 143988
rect 268150 143986 268210 144364
rect 282821 143986 282887 143989
rect 233804 143926 268210 143986
rect 279956 143984 282887 143986
rect 279956 143928 282826 143984
rect 282882 143928 282887 143984
rect 279956 143926 282887 143928
rect 233804 143924 233810 143926
rect 282821 143923 282887 143926
rect 213269 143578 213335 143581
rect 217182 143578 217242 143820
rect 213269 143576 217242 143578
rect 213269 143520 213274 143576
rect 213330 143520 217242 143576
rect 213269 143518 217242 143520
rect 265801 143578 265867 143581
rect 268150 143578 268210 143820
rect 265801 143576 268210 143578
rect 265801 143520 265806 143576
rect 265862 143520 268210 143576
rect 265801 143518 268210 143520
rect 213269 143515 213335 143518
rect 265801 143515 265867 143518
rect 231761 143442 231827 143445
rect 228968 143440 231827 143442
rect 228968 143384 231766 143440
rect 231822 143384 231827 143440
rect 228968 143382 231827 143384
rect 231761 143379 231827 143382
rect 214005 142762 214071 142765
rect 217182 142762 217242 143276
rect 264973 143170 265039 143173
rect 268150 143170 268210 143412
rect 282085 143170 282151 143173
rect 264973 143168 268210 143170
rect 264973 143112 264978 143168
rect 265034 143112 268210 143168
rect 264973 143110 268210 143112
rect 279956 143168 282151 143170
rect 279956 143112 282090 143168
rect 282146 143112 282151 143168
rect 279956 143110 282151 143112
rect 264973 143107 265039 143110
rect 282085 143107 282151 143110
rect 242934 143034 242940 143036
rect 228968 142974 242940 143034
rect 242934 142972 242940 142974
rect 243004 142972 243010 143036
rect 265433 142898 265499 142901
rect 258030 142896 265499 142898
rect 258030 142840 265438 142896
rect 265494 142840 265499 142896
rect 258030 142838 265499 142840
rect 214005 142760 217242 142762
rect 214005 142704 214010 142760
rect 214066 142704 217242 142760
rect 214005 142702 217242 142704
rect 214005 142699 214071 142702
rect 233918 142700 233924 142764
rect 233988 142762 233994 142764
rect 258030 142762 258090 142838
rect 265433 142835 265499 142838
rect 233988 142702 258090 142762
rect 265341 142762 265407 142765
rect 268150 142762 268210 143004
rect 265341 142760 268210 142762
rect 265341 142704 265346 142760
rect 265402 142704 268210 142760
rect 265341 142702 268210 142704
rect 233988 142700 233994 142702
rect 265341 142699 265407 142702
rect 213913 142354 213979 142357
rect 217182 142354 217242 142596
rect 230473 142490 230539 142493
rect 228968 142488 230539 142490
rect 228968 142432 230478 142488
rect 230534 142432 230539 142488
rect 228968 142430 230539 142432
rect 230473 142427 230539 142430
rect 213913 142352 217242 142354
rect 213913 142296 213918 142352
rect 213974 142296 217242 142352
rect 213913 142294 217242 142296
rect 265801 142354 265867 142357
rect 268150 142354 268210 142596
rect 282269 142490 282335 142493
rect 279956 142488 282335 142490
rect 279956 142432 282274 142488
rect 282330 142432 282335 142488
rect 279956 142430 282335 142432
rect 282269 142427 282335 142430
rect 265801 142352 268210 142354
rect 265801 142296 265806 142352
rect 265862 142296 268210 142352
rect 265801 142294 268210 142296
rect 213913 142291 213979 142294
rect 265801 142291 265867 142294
rect 265249 142218 265315 142221
rect 265249 142216 267842 142218
rect 265249 142160 265254 142216
rect 265310 142160 267842 142216
rect 265249 142158 267842 142160
rect 265249 142155 265315 142158
rect 229737 142082 229803 142085
rect 228968 142080 229803 142082
rect 228968 142024 229742 142080
rect 229798 142024 229803 142080
rect 228968 142022 229803 142024
rect 229737 142019 229803 142022
rect 267782 141946 267842 142158
rect 268334 141946 268394 142188
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 267782 141886 268394 141946
rect 245878 141674 245884 141676
rect 228968 141614 245884 141674
rect 245878 141612 245884 141614
rect 245948 141612 245954 141676
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 214005 141339 214071 141342
rect 231342 141340 231348 141404
rect 231412 141402 231418 141404
rect 262949 141402 263015 141405
rect 231412 141400 263015 141402
rect 231412 141344 262954 141400
rect 263010 141344 263015 141400
rect 231412 141342 263015 141344
rect 231412 141340 231418 141342
rect 262949 141339 263015 141342
rect 265893 141402 265959 141405
rect 268150 141402 268210 141780
rect 282821 141674 282887 141677
rect 279956 141672 282887 141674
rect 279956 141616 282826 141672
rect 282882 141616 282887 141672
rect 279956 141614 282887 141616
rect 282821 141611 282887 141614
rect 265893 141400 268210 141402
rect 265893 141344 265898 141400
rect 265954 141344 268210 141400
rect 265893 141342 268210 141344
rect 265893 141339 265959 141342
rect 213913 140994 213979 140997
rect 217182 140994 217242 141236
rect 241646 141130 241652 141132
rect 228968 141070 241652 141130
rect 241646 141068 241652 141070
rect 241716 141068 241722 141132
rect 213913 140992 217242 140994
rect 213913 140936 213918 140992
rect 213974 140936 217242 140992
rect 213913 140934 217242 140936
rect 265525 140994 265591 140997
rect 268518 140996 268578 141236
rect 265525 140992 268210 140994
rect 265525 140936 265530 140992
rect 265586 140936 268210 140992
rect 265525 140934 268210 140936
rect 213913 140931 213979 140934
rect 265525 140931 265591 140934
rect 268150 140828 268210 140934
rect 268510 140932 268516 140996
rect 268580 140932 268586 140996
rect 282729 140858 282795 140861
rect 279956 140856 282795 140858
rect 279956 140800 282734 140856
rect 282790 140800 282795 140856
rect 279956 140798 282795 140800
rect 282729 140795 282795 140798
rect 231761 140722 231827 140725
rect 228968 140720 231827 140722
rect 228968 140664 231766 140720
rect 231822 140664 231827 140720
rect 228968 140662 231827 140664
rect 231761 140659 231827 140662
rect 264421 140586 264487 140589
rect 268510 140586 268516 140588
rect 264421 140584 268516 140586
rect 213913 140042 213979 140045
rect 217182 140042 217242 140556
rect 264421 140528 264426 140584
rect 264482 140528 268516 140584
rect 264421 140526 268516 140528
rect 264421 140523 264487 140526
rect 268510 140524 268516 140526
rect 268580 140524 268586 140588
rect 230933 140178 230999 140181
rect 228968 140176 230999 140178
rect 228968 140120 230938 140176
rect 230994 140120 230999 140176
rect 228968 140118 230999 140120
rect 230933 140115 230999 140118
rect 262806 140116 262812 140180
rect 262876 140178 262882 140180
rect 268150 140178 268210 140420
rect 282821 140178 282887 140181
rect 262876 140118 268210 140178
rect 279956 140176 282887 140178
rect 279956 140120 282826 140176
rect 282882 140120 282887 140176
rect 279956 140118 282887 140120
rect 262876 140116 262882 140118
rect 282821 140115 282887 140118
rect 213913 140040 217242 140042
rect 213913 139984 213918 140040
rect 213974 139984 217242 140040
rect 213913 139982 217242 139984
rect 213913 139979 213979 139982
rect 214005 139498 214071 139501
rect 217182 139498 217242 139876
rect 231485 139770 231551 139773
rect 228968 139768 231551 139770
rect 228968 139712 231490 139768
rect 231546 139712 231551 139768
rect 228968 139710 231551 139712
rect 231485 139707 231551 139710
rect 265709 139770 265775 139773
rect 268150 139770 268210 140012
rect 265709 139768 268210 139770
rect 265709 139712 265714 139768
rect 265770 139712 268210 139768
rect 265709 139710 268210 139712
rect 265709 139707 265775 139710
rect 214005 139496 217242 139498
rect 214005 139440 214010 139496
rect 214066 139440 217242 139496
rect 214005 139438 217242 139440
rect 265801 139498 265867 139501
rect 265801 139496 267842 139498
rect 265801 139440 265806 139496
rect 265862 139440 267842 139496
rect 265801 139438 267842 139440
rect 214005 139435 214071 139438
rect 265801 139435 265867 139438
rect 267782 139362 267842 139438
rect 268334 139362 268394 139604
rect 282821 139362 282887 139365
rect 267782 139302 268394 139362
rect 279956 139360 282887 139362
rect 279956 139304 282826 139360
rect 282882 139304 282887 139360
rect 279956 139302 282887 139304
rect 282821 139299 282887 139302
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 231669 139226 231735 139229
rect 228968 139224 231735 139226
rect 213913 138818 213979 138821
rect 217182 138818 217242 139196
rect 228968 139168 231674 139224
rect 231730 139168 231735 139224
rect 583520 139212 584960 139302
rect 228968 139166 231735 139168
rect 231669 139163 231735 139166
rect 231761 138818 231827 138821
rect 268150 138818 268210 139196
rect 213913 138816 217242 138818
rect 213913 138760 213918 138816
rect 213974 138760 217242 138816
rect 213913 138758 217242 138760
rect 228968 138816 231827 138818
rect 228968 138760 231766 138816
rect 231822 138760 231827 138816
rect 228968 138758 231827 138760
rect 213913 138755 213979 138758
rect 231761 138755 231827 138758
rect 258030 138758 268210 138818
rect 214649 138138 214715 138141
rect 217182 138138 217242 138652
rect 232446 138348 232452 138412
rect 232516 138410 232522 138412
rect 258030 138410 258090 138758
rect 232516 138350 258090 138410
rect 265801 138410 265867 138413
rect 268150 138410 268210 138652
rect 282729 138546 282795 138549
rect 279956 138544 282795 138546
rect 279956 138488 282734 138544
rect 282790 138488 282795 138544
rect 279956 138486 282795 138488
rect 282729 138483 282795 138486
rect 265801 138408 268210 138410
rect 265801 138352 265806 138408
rect 265862 138352 268210 138408
rect 265801 138350 268210 138352
rect 232516 138348 232522 138350
rect 265801 138347 265867 138350
rect 236494 138274 236500 138276
rect 228968 138214 236500 138274
rect 236494 138212 236500 138214
rect 236564 138212 236570 138276
rect 214649 138136 217242 138138
rect 214649 138080 214654 138136
rect 214710 138080 217242 138136
rect 214649 138078 217242 138080
rect 265157 138138 265223 138141
rect 265157 138136 267842 138138
rect 265157 138080 265162 138136
rect 265218 138080 267842 138136
rect 265157 138078 267842 138080
rect 214649 138075 214715 138078
rect 265157 138075 265223 138078
rect 267782 138002 267842 138078
rect 268334 138002 268394 138244
rect 213913 137458 213979 137461
rect 217182 137458 217242 137972
rect 267782 137942 268394 138002
rect 234654 137866 234660 137868
rect 228968 137806 234660 137866
rect 234654 137804 234660 137806
rect 234724 137804 234730 137868
rect 282821 137866 282887 137869
rect 279956 137864 282887 137866
rect 265801 137594 265867 137597
rect 268150 137594 268210 137836
rect 279956 137808 282826 137864
rect 282882 137808 282887 137864
rect 279956 137806 282887 137808
rect 282821 137803 282887 137806
rect 265801 137592 268210 137594
rect 265801 137536 265806 137592
rect 265862 137536 268210 137592
rect 265801 137534 268210 137536
rect 265801 137531 265867 137534
rect 213913 137456 217242 137458
rect 213913 137400 213918 137456
rect 213974 137400 217242 137456
rect 213913 137398 217242 137400
rect 213913 137395 213979 137398
rect 231761 137322 231827 137325
rect 228968 137320 231827 137322
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 170254 136716 170260 136780
rect 170324 136778 170330 136780
rect 217182 136778 217242 137292
rect 228968 137264 231766 137320
rect 231822 137264 231827 137320
rect 228968 137262 231827 137264
rect 231761 137259 231827 137262
rect 265709 137186 265775 137189
rect 268150 137186 268210 137428
rect 265709 137184 268210 137186
rect 265709 137128 265714 137184
rect 265770 137128 268210 137184
rect 265709 137126 268210 137128
rect 265709 137123 265775 137126
rect 280286 137050 280292 137052
rect 231485 136914 231551 136917
rect 228968 136912 231551 136914
rect 228968 136856 231490 136912
rect 231546 136856 231551 136912
rect 228968 136854 231551 136856
rect 231485 136851 231551 136854
rect 170324 136718 217242 136778
rect 266077 136778 266143 136781
rect 268150 136778 268210 137020
rect 279956 136990 280292 137050
rect 280286 136988 280292 136990
rect 280356 136988 280362 137052
rect 266077 136776 268210 136778
rect 266077 136720 266082 136776
rect 266138 136720 268210 136776
rect 266077 136718 268210 136720
rect 170324 136716 170330 136718
rect 266077 136715 266143 136718
rect 217182 136098 217242 136612
rect 231761 136370 231827 136373
rect 228968 136368 231827 136370
rect 228968 136312 231766 136368
rect 231822 136312 231827 136368
rect 228968 136310 231827 136312
rect 231761 136307 231827 136310
rect 265985 136370 266051 136373
rect 268150 136370 268210 136612
rect 282821 136370 282887 136373
rect 265985 136368 268210 136370
rect 265985 136312 265990 136368
rect 266046 136312 268210 136368
rect 265985 136310 268210 136312
rect 279956 136368 282887 136370
rect 279956 136312 282826 136368
rect 282882 136312 282887 136368
rect 279956 136310 282887 136312
rect 265985 136307 266051 136310
rect 282821 136307 282887 136310
rect 200070 136038 217242 136098
rect 166390 135492 166396 135556
rect 166460 135554 166466 135556
rect 200070 135554 200130 136038
rect 231669 135962 231735 135965
rect 228968 135960 231735 135962
rect 214005 135690 214071 135693
rect 217182 135690 217242 135932
rect 228968 135904 231674 135960
rect 231730 135904 231735 135960
rect 228968 135902 231735 135904
rect 231669 135899 231735 135902
rect 231577 135826 231643 135829
rect 239070 135826 239076 135828
rect 231577 135824 239076 135826
rect 231577 135768 231582 135824
rect 231638 135768 239076 135824
rect 231577 135766 239076 135768
rect 231577 135763 231643 135766
rect 239070 135764 239076 135766
rect 239140 135764 239146 135828
rect 239254 135764 239260 135828
rect 239324 135826 239330 135828
rect 268150 135826 268210 136204
rect 239324 135766 268210 135826
rect 239324 135764 239330 135766
rect 214005 135688 217242 135690
rect 214005 135632 214010 135688
rect 214066 135632 217242 135688
rect 214005 135630 217242 135632
rect 214005 135627 214071 135630
rect 166460 135494 200130 135554
rect 166460 135492 166466 135494
rect 213913 135418 213979 135421
rect 231393 135418 231459 135421
rect 213913 135416 217242 135418
rect 213913 135360 213918 135416
rect 213974 135360 217242 135416
rect 213913 135358 217242 135360
rect 228968 135416 231459 135418
rect 228968 135360 231398 135416
rect 231454 135360 231459 135416
rect 228968 135358 231459 135360
rect 213913 135355 213979 135358
rect 217182 135252 217242 135358
rect 231393 135355 231459 135358
rect 265801 135418 265867 135421
rect 268150 135418 268210 135660
rect 282729 135554 282795 135557
rect 279956 135552 282795 135554
rect 279956 135496 282734 135552
rect 282790 135496 282795 135552
rect 279956 135494 282795 135496
rect 282729 135491 282795 135494
rect 265801 135416 268210 135418
rect 265801 135360 265806 135416
rect 265862 135360 268210 135416
rect 265801 135358 268210 135360
rect 265801 135355 265867 135358
rect 265157 135282 265223 135285
rect 265157 135280 267842 135282
rect 265157 135224 265162 135280
rect 265218 135224 267842 135280
rect 265157 135222 267842 135224
rect 265157 135219 265223 135222
rect 231761 135010 231827 135013
rect 228968 135008 231827 135010
rect 228968 134952 231766 135008
rect 231822 134952 231827 135008
rect 228968 134950 231827 134952
rect 267782 135010 267842 135222
rect 268334 135010 268394 135252
rect 267782 134950 268394 135010
rect 231761 134947 231827 134950
rect 265249 134602 265315 134605
rect 268150 134602 268210 134844
rect 282821 134738 282887 134741
rect 279956 134736 282887 134738
rect 279956 134680 282826 134736
rect 282882 134680 282887 134736
rect 279956 134678 282887 134680
rect 282821 134675 282887 134678
rect 265249 134600 268210 134602
rect 214005 134330 214071 134333
rect 217182 134330 217242 134572
rect 265249 134544 265254 134600
rect 265310 134544 268210 134600
rect 265249 134542 268210 134544
rect 265249 134539 265315 134542
rect 231669 134466 231735 134469
rect 228968 134464 231735 134466
rect 228968 134408 231674 134464
rect 231730 134408 231735 134464
rect 228968 134406 231735 134408
rect 231669 134403 231735 134406
rect 214005 134328 217242 134330
rect 214005 134272 214010 134328
rect 214066 134272 217242 134328
rect 214005 134270 217242 134272
rect 214005 134267 214071 134270
rect 265801 134194 265867 134197
rect 268518 134196 268578 134436
rect 265801 134192 268210 134194
rect 265801 134136 265806 134192
rect 265862 134136 268210 134192
rect 265801 134134 268210 134136
rect 265801 134131 265867 134134
rect 213913 134058 213979 134061
rect 230749 134058 230815 134061
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 228968 134056 230815 134058
rect 228968 134000 230754 134056
rect 230810 134000 230815 134056
rect 268150 134028 268210 134134
rect 268510 134132 268516 134196
rect 268580 134132 268586 134196
rect 282729 134058 282795 134061
rect 279956 134056 282795 134058
rect 228968 133998 230815 134000
rect 279956 134000 282734 134056
rect 282790 134000 282795 134056
rect 279956 133998 282795 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 230749 133995 230815 133998
rect 282729 133995 282795 133998
rect 231301 133788 231367 133789
rect 231301 133786 231348 133788
rect 231256 133784 231348 133786
rect 231256 133728 231306 133784
rect 231256 133726 231348 133728
rect 231301 133724 231348 133726
rect 231412 133724 231418 133788
rect 264421 133786 264487 133789
rect 268510 133786 268516 133788
rect 264421 133784 268516 133786
rect 264421 133728 264426 133784
rect 264482 133728 268516 133784
rect 264421 133726 268516 133728
rect 231301 133723 231367 133724
rect 264421 133723 264487 133726
rect 268510 133724 268516 133726
rect 268580 133724 268586 133788
rect 231761 133514 231827 133517
rect 228968 133512 231827 133514
rect 228968 133456 231766 133512
rect 231822 133456 231827 133512
rect 228968 133454 231827 133456
rect 231761 133451 231827 133454
rect 170438 132772 170444 132836
rect 170508 132834 170514 132836
rect 217182 132834 217242 133348
rect 262070 133180 262076 133244
rect 262140 133242 262146 133244
rect 268150 133242 268210 133620
rect 281901 133242 281967 133245
rect 262140 133182 268210 133242
rect 279956 133240 281967 133242
rect 279956 133184 281906 133240
rect 281962 133184 281967 133240
rect 279956 133182 281967 133184
rect 262140 133180 262146 133182
rect 281901 133179 281967 133182
rect 231669 133106 231735 133109
rect 264237 133106 264303 133109
rect 228968 133104 231735 133106
rect 228968 133048 231674 133104
rect 231730 133048 231735 133104
rect 228968 133046 231735 133048
rect 231669 133043 231735 133046
rect 238710 133104 264303 133106
rect 238710 133048 264242 133104
rect 264298 133048 264303 133104
rect 238710 133046 264303 133048
rect 231158 132908 231164 132972
rect 231228 132970 231234 132972
rect 238710 132970 238770 133046
rect 264237 133043 264303 133046
rect 231228 132910 238770 132970
rect 231228 132908 231234 132910
rect 170508 132774 217242 132834
rect 265617 132834 265683 132837
rect 268150 132834 268210 133076
rect 265617 132832 268210 132834
rect 265617 132776 265622 132832
rect 265678 132776 268210 132832
rect 265617 132774 268210 132776
rect 170508 132772 170514 132774
rect 265617 132771 265683 132774
rect 214557 132562 214623 132565
rect 214557 132560 216874 132562
rect 214557 132504 214562 132560
rect 214618 132504 216874 132560
rect 214557 132502 216874 132504
rect 214557 132499 214623 132502
rect 216814 132426 216874 132502
rect 217366 132426 217426 132668
rect 231025 132562 231091 132565
rect 228968 132560 231091 132562
rect 228968 132504 231030 132560
rect 231086 132504 231091 132560
rect 228968 132502 231091 132504
rect 231025 132499 231091 132502
rect 264094 132500 264100 132564
rect 264164 132562 264170 132564
rect 264164 132502 267842 132562
rect 264164 132500 264170 132502
rect 216814 132366 217426 132426
rect 267782 132426 267842 132502
rect 268334 132426 268394 132668
rect 282729 132426 282795 132429
rect 267782 132366 268394 132426
rect 279956 132424 282795 132426
rect 279956 132368 282734 132424
rect 282790 132368 282795 132424
rect 279956 132366 282795 132368
rect 282729 132363 282795 132366
rect 230749 132154 230815 132157
rect 228968 132152 230815 132154
rect 228968 132096 230754 132152
rect 230810 132096 230815 132152
rect 228968 132094 230815 132096
rect 230749 132091 230815 132094
rect 265709 132018 265775 132021
rect 268150 132018 268210 132260
rect 265709 132016 268210 132018
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 265709 131960 265714 132016
rect 265770 131960 268210 132016
rect 265709 131958 268210 131960
rect 265709 131955 265775 131958
rect 231485 131610 231551 131613
rect 228968 131608 231551 131610
rect 228968 131552 231490 131608
rect 231546 131552 231551 131608
rect 228968 131550 231551 131552
rect 231485 131547 231551 131550
rect 258758 131548 258764 131612
rect 258828 131610 258834 131612
rect 268150 131610 268210 131852
rect 282821 131746 282887 131749
rect 279956 131744 282887 131746
rect 279956 131688 282826 131744
rect 282882 131688 282887 131744
rect 279956 131686 282887 131688
rect 282821 131683 282887 131686
rect 258828 131550 268210 131610
rect 258828 131548 258834 131550
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 214005 131411 214071 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 231761 131202 231827 131205
rect 228968 131200 231827 131202
rect 228968 131144 231766 131200
rect 231822 131144 231827 131200
rect 228968 131142 231827 131144
rect 231761 131139 231827 131142
rect 265617 131202 265683 131205
rect 268150 131202 268210 131444
rect 265617 131200 268210 131202
rect 265617 131144 265622 131200
rect 265678 131144 268210 131200
rect 265617 131142 268210 131144
rect 265617 131139 265683 131142
rect 216814 131006 217426 131066
rect 261293 130794 261359 130797
rect 268334 130794 268394 131036
rect 282269 130930 282335 130933
rect 279956 130928 282335 130930
rect 279956 130872 282274 130928
rect 282330 130872 282335 130928
rect 279956 130870 282335 130872
rect 282269 130867 282335 130870
rect 261293 130792 268394 130794
rect 261293 130736 261298 130792
rect 261354 130736 268394 130792
rect 261293 130734 268394 130736
rect 261293 130731 261359 130734
rect 231761 130658 231827 130661
rect 228968 130656 231827 130658
rect 213913 130114 213979 130117
rect 217182 130114 217242 130628
rect 228968 130600 231766 130656
rect 231822 130600 231827 130656
rect 228968 130598 231827 130600
rect 231761 130595 231827 130598
rect 264421 130658 264487 130661
rect 264421 130656 268210 130658
rect 264421 130600 264426 130656
rect 264482 130600 268210 130656
rect 264421 130598 268210 130600
rect 264421 130595 264487 130598
rect 268150 130492 268210 130598
rect 231485 130250 231551 130253
rect 228968 130248 231551 130250
rect 228968 130192 231490 130248
rect 231546 130192 231551 130248
rect 228968 130190 231551 130192
rect 231485 130187 231551 130190
rect 258574 130188 258580 130252
rect 258644 130250 258650 130252
rect 258644 130190 268210 130250
rect 258644 130188 258650 130190
rect 213913 130112 217242 130114
rect 213913 130056 213918 130112
rect 213974 130056 217242 130112
rect 268150 130084 268210 130190
rect 281717 130114 281783 130117
rect 279956 130112 281783 130114
rect 213913 130054 217242 130056
rect 279956 130056 281722 130112
rect 281778 130056 281783 130112
rect 279956 130054 281783 130056
rect 213913 130051 213979 130054
rect 281717 130051 281783 130054
rect 168966 129780 168972 129844
rect 169036 129842 169042 129844
rect 169036 129782 216874 129842
rect 169036 129780 169042 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 231393 129842 231459 129845
rect 228968 129840 231459 129842
rect 228968 129784 231398 129840
rect 231454 129784 231459 129840
rect 228968 129782 231459 129784
rect 231393 129779 231459 129782
rect 216814 129646 217426 129706
rect 268150 129434 268210 129676
rect 258030 129374 268210 129434
rect 67449 129298 67515 129301
rect 68142 129298 68816 129304
rect 231761 129298 231827 129301
rect 67449 129296 68816 129298
rect 67449 129240 67454 129296
rect 67510 129244 68816 129296
rect 228968 129296 231827 129298
rect 67510 129240 68202 129244
rect 67449 129238 68202 129240
rect 67449 129235 67515 129238
rect 217182 128890 217242 129268
rect 228968 129240 231766 129296
rect 231822 129240 231827 129296
rect 228968 129238 231827 129240
rect 231761 129235 231827 129238
rect 257286 128964 257292 129028
rect 257356 129026 257362 129028
rect 258030 129026 258090 129374
rect 257356 128966 258090 129026
rect 265341 129026 265407 129029
rect 268150 129026 268210 129268
rect 265341 129024 268210 129026
rect 265341 128968 265346 129024
rect 265402 128968 268210 129024
rect 265341 128966 268210 128968
rect 257356 128964 257362 128966
rect 265341 128963 265407 128966
rect 231669 128890 231735 128893
rect 200070 128830 217242 128890
rect 228968 128888 231735 128890
rect 228968 128832 231674 128888
rect 231730 128832 231735 128888
rect 228968 128830 231735 128832
rect 173198 128420 173204 128484
rect 173268 128482 173274 128484
rect 200070 128482 200130 128830
rect 231669 128827 231735 128830
rect 173268 128422 200130 128482
rect 213913 128482 213979 128485
rect 217182 128482 217242 128724
rect 265801 128618 265867 128621
rect 268518 128620 268578 128860
rect 279926 128754 279986 129404
rect 287278 128754 287284 128756
rect 279926 128694 287284 128754
rect 287278 128692 287284 128694
rect 287348 128692 287354 128756
rect 265801 128616 268210 128618
rect 265801 128560 265806 128616
rect 265862 128560 268210 128616
rect 265801 128558 268210 128560
rect 265801 128555 265867 128558
rect 213913 128480 217242 128482
rect 213913 128424 213918 128480
rect 213974 128424 217242 128480
rect 268150 128452 268210 128558
rect 268510 128556 268516 128620
rect 268580 128556 268586 128620
rect 282821 128618 282887 128621
rect 279956 128616 282887 128618
rect 279956 128560 282826 128616
rect 282882 128560 282887 128616
rect 279956 128558 282887 128560
rect 282821 128555 282887 128558
rect 213913 128422 217242 128424
rect 173268 128420 173274 128422
rect 213913 128419 213979 128422
rect 231761 128346 231827 128349
rect 228968 128344 231827 128346
rect 228968 128288 231766 128344
rect 231822 128288 231827 128344
rect 228968 128286 231827 128288
rect 231761 128283 231827 128286
rect 264421 128210 264487 128213
rect 268510 128210 268516 128212
rect 264421 128208 268516 128210
rect 264421 128152 264426 128208
rect 264482 128152 268516 128208
rect 264421 128150 268516 128152
rect 264421 128147 264487 128150
rect 268510 128148 268516 128150
rect 268580 128148 268586 128212
rect 66161 128074 66227 128077
rect 68142 128074 68816 128080
rect 66161 128072 68816 128074
rect 66161 128016 66166 128072
rect 66222 128020 68816 128072
rect 66222 128016 68202 128020
rect 66161 128014 68202 128016
rect 66161 128011 66227 128014
rect 213913 127530 213979 127533
rect 217182 127530 217242 128044
rect 230749 127938 230815 127941
rect 228968 127936 230815 127938
rect 228968 127880 230754 127936
rect 230810 127880 230815 127936
rect 228968 127878 230815 127880
rect 230749 127875 230815 127878
rect 265341 127666 265407 127669
rect 268150 127666 268210 127908
rect 281901 127802 281967 127805
rect 279956 127800 281967 127802
rect 279956 127744 281906 127800
rect 281962 127744 281967 127800
rect 279956 127742 281967 127744
rect 281901 127739 281967 127742
rect 265341 127664 268210 127666
rect 265341 127608 265346 127664
rect 265402 127608 268210 127664
rect 265341 127606 268210 127608
rect 265341 127603 265407 127606
rect 213913 127528 217242 127530
rect 213913 127472 213918 127528
rect 213974 127472 217242 127528
rect 213913 127470 217242 127472
rect 213913 127467 213979 127470
rect 231669 127394 231735 127397
rect 228968 127392 231735 127394
rect 169150 127196 169156 127260
rect 169220 127258 169226 127260
rect 169220 127198 200130 127258
rect 169220 127196 169226 127198
rect 200070 127122 200130 127198
rect 217366 127122 217426 127364
rect 228968 127336 231674 127392
rect 231730 127336 231735 127392
rect 228968 127334 231735 127336
rect 231669 127331 231735 127334
rect 268518 127260 268578 127500
rect 258030 127198 268210 127258
rect 200070 127062 217426 127122
rect 255814 127060 255820 127124
rect 255884 127122 255890 127124
rect 258030 127122 258090 127198
rect 255884 127062 258090 127122
rect 268150 127092 268210 127198
rect 268510 127196 268516 127260
rect 268580 127196 268586 127260
rect 288566 127122 288572 127124
rect 279956 127062 288572 127122
rect 255884 127060 255890 127062
rect 288566 127060 288572 127062
rect 288636 127060 288642 127124
rect 231577 126986 231643 126989
rect 228968 126984 231643 126986
rect 228968 126928 231582 126984
rect 231638 126928 231643 126984
rect 228968 126926 231643 126928
rect 231577 126923 231643 126926
rect 264421 126850 264487 126853
rect 268510 126850 268516 126852
rect 264421 126848 268516 126850
rect 264421 126792 264426 126848
rect 264482 126792 268516 126848
rect 264421 126790 268516 126792
rect 264421 126787 264487 126790
rect 268510 126788 268516 126790
rect 268580 126788 268586 126852
rect 67541 126306 67607 126309
rect 68142 126306 68816 126312
rect 67541 126304 68816 126306
rect 67541 126248 67546 126304
rect 67602 126252 68816 126304
rect 67602 126248 68202 126252
rect 67541 126246 68202 126248
rect 67541 126243 67607 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 231761 126442 231827 126445
rect 228968 126440 231827 126442
rect 228968 126384 231766 126440
rect 231822 126384 231827 126440
rect 228968 126382 231827 126384
rect 231761 126379 231827 126382
rect 265801 126442 265867 126445
rect 268150 126442 268210 126684
rect 265801 126440 268210 126442
rect 265801 126384 265806 126440
rect 265862 126384 268210 126440
rect 265801 126382 268210 126384
rect 265801 126379 265867 126382
rect 231710 126244 231716 126308
rect 231780 126306 231786 126308
rect 253473 126306 253539 126309
rect 282821 126306 282887 126309
rect 231780 126304 253539 126306
rect 231780 126248 253478 126304
rect 253534 126248 253539 126304
rect 279956 126304 282887 126306
rect 231780 126246 253539 126248
rect 231780 126244 231786 126246
rect 253473 126243 253539 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 230974 126034 230980 126036
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 228968 125974 230980 126034
rect 230974 125972 230980 125974
rect 231044 125972 231050 126036
rect 265617 126034 265683 126037
rect 268150 126034 268210 126276
rect 279956 126248 282826 126304
rect 282882 126248 282887 126304
rect 279956 126246 282887 126248
rect 282821 126243 282887 126246
rect 265617 126032 268210 126034
rect 265617 125976 265622 126032
rect 265678 125976 268210 126032
rect 265617 125974 268210 125976
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 265617 125971 265683 125974
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 213913 125699 213979 125702
rect 265709 125626 265775 125629
rect 268334 125626 268394 125868
rect 265709 125624 268394 125626
rect 265709 125568 265714 125624
rect 265770 125568 268394 125624
rect 265709 125566 268394 125568
rect 265709 125563 265775 125566
rect 231710 125490 231716 125492
rect 228968 125430 231716 125490
rect 231710 125428 231716 125430
rect 231780 125428 231786 125492
rect 282821 125490 282887 125493
rect 279956 125488 282887 125490
rect 279956 125432 282826 125488
rect 282882 125432 282887 125488
rect 279956 125430 282887 125432
rect 282821 125427 282887 125430
rect 65517 125218 65583 125221
rect 68142 125218 68816 125224
rect 65517 125216 68816 125218
rect 65517 125160 65522 125216
rect 65578 125164 68816 125216
rect 65578 125160 68202 125164
rect 65517 125158 68202 125160
rect 65517 125155 65583 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 230422 125292 230428 125356
rect 230492 125354 230498 125356
rect 231301 125354 231367 125357
rect 230492 125352 231367 125354
rect 230492 125296 231306 125352
rect 231362 125296 231367 125352
rect 230492 125294 231367 125296
rect 230492 125292 230498 125294
rect 231301 125291 231367 125294
rect 231761 125082 231827 125085
rect 228968 125080 231827 125082
rect 228968 125024 231766 125080
rect 231822 125024 231827 125080
rect 228968 125022 231827 125024
rect 231761 125019 231827 125022
rect 265801 125082 265867 125085
rect 268150 125082 268210 125324
rect 265801 125080 268210 125082
rect 265801 125024 265806 125080
rect 265862 125024 268210 125080
rect 265801 125022 268210 125024
rect 265801 125019 265867 125022
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 214005 124747 214071 124750
rect 265893 124674 265959 124677
rect 268150 124674 268210 124916
rect 282729 124810 282795 124813
rect 279956 124808 282795 124810
rect 279956 124752 282734 124808
rect 282790 124752 282795 124808
rect 279956 124750 282795 124752
rect 282729 124747 282795 124750
rect 265893 124672 268210 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 265893 124616 265898 124672
rect 265954 124616 268210 124672
rect 265893 124614 268210 124616
rect 265893 124611 265959 124614
rect 231485 124538 231551 124541
rect 228968 124536 231551 124538
rect 228968 124480 231490 124536
rect 231546 124480 231551 124536
rect 228968 124478 231551 124480
rect 231485 124475 231551 124478
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 213913 124339 213979 124342
rect 265525 124266 265591 124269
rect 268334 124266 268394 124508
rect 265525 124264 268394 124266
rect 265525 124208 265530 124264
rect 265586 124208 268394 124264
rect 265525 124206 268394 124208
rect 265525 124203 265591 124206
rect 231761 124130 231827 124133
rect 228968 124128 231827 124130
rect -960 123572 480 123812
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 228968 124072 231766 124128
rect 231822 124072 231827 124128
rect 228968 124070 231827 124072
rect 231761 124067 231827 124070
rect 267181 123858 267247 123861
rect 268150 123858 268210 124100
rect 281993 123994 282059 123997
rect 279956 123992 282059 123994
rect 279956 123936 281998 123992
rect 282054 123936 282059 123992
rect 279956 123934 282059 123936
rect 281993 123931 282059 123934
rect 267181 123856 268210 123858
rect 267181 123800 267186 123856
rect 267242 123800 268210 123856
rect 267181 123798 268210 123800
rect 267181 123795 267247 123798
rect 231158 123586 231164 123588
rect 214005 123584 217242 123586
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 228968 123526 231164 123586
rect 66069 123523 66135 123526
rect 214005 123523 214071 123526
rect 231158 123524 231164 123526
rect 231228 123524 231234 123588
rect 265893 123450 265959 123453
rect 268150 123450 268210 123692
rect 265893 123448 268210 123450
rect 213913 122906 213979 122909
rect 217182 122906 217242 123420
rect 265893 123392 265898 123448
rect 265954 123392 268210 123448
rect 265893 123390 268210 123392
rect 265893 123387 265959 123390
rect 231577 123178 231643 123181
rect 228968 123176 231643 123178
rect 228968 123120 231582 123176
rect 231638 123120 231643 123176
rect 228968 123118 231643 123120
rect 231577 123115 231643 123118
rect 265801 123042 265867 123045
rect 268518 123044 268578 123284
rect 282177 123178 282243 123181
rect 279956 123176 282243 123178
rect 279956 123120 282182 123176
rect 282238 123120 282243 123176
rect 279956 123118 282243 123120
rect 282177 123115 282243 123118
rect 265801 123040 268210 123042
rect 265801 122984 265806 123040
rect 265862 122984 268210 123040
rect 265801 122982 268210 122984
rect 265801 122979 265867 122982
rect 213913 122904 217242 122906
rect 213913 122848 213918 122904
rect 213974 122848 217242 122904
rect 268150 122876 268210 122982
rect 268510 122980 268516 123044
rect 268580 122980 268586 123044
rect 213913 122846 217242 122848
rect 213913 122843 213979 122846
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 66069 122571 66135 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 231761 122634 231827 122637
rect 228968 122632 231827 122634
rect 228968 122576 231766 122632
rect 231822 122576 231827 122632
rect 228968 122574 231827 122576
rect 231761 122571 231827 122574
rect 264421 122634 264487 122637
rect 268510 122634 268516 122636
rect 264421 122632 268516 122634
rect 264421 122576 264426 122632
rect 264482 122576 268516 122632
rect 264421 122574 268516 122576
rect 264421 122571 264487 122574
rect 268510 122572 268516 122574
rect 268580 122572 268586 122636
rect 282085 122498 282151 122501
rect 279956 122496 282151 122498
rect 279956 122440 282090 122496
rect 282146 122440 282151 122496
rect 279956 122438 282151 122440
rect 282085 122435 282151 122438
rect 230933 122226 230999 122229
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 228968 122224 230999 122226
rect 228968 122168 230938 122224
rect 230994 122168 230999 122224
rect 228968 122166 230999 122168
rect 214005 122163 214071 122166
rect 230933 122163 230999 122166
rect 265893 122090 265959 122093
rect 268150 122090 268210 122332
rect 265893 122088 268210 122090
rect 213913 121546 213979 121549
rect 217182 121546 217242 122060
rect 265893 122032 265898 122088
rect 265954 122032 268210 122088
rect 265893 122030 268210 122032
rect 265893 122027 265959 122030
rect 231485 121682 231551 121685
rect 228968 121680 231551 121682
rect 228968 121624 231490 121680
rect 231546 121624 231551 121680
rect 228968 121622 231551 121624
rect 231485 121619 231551 121622
rect 265801 121682 265867 121685
rect 268518 121684 268578 121924
rect 265801 121680 268210 121682
rect 265801 121624 265806 121680
rect 265862 121624 268210 121680
rect 265801 121622 268210 121624
rect 265801 121619 265867 121622
rect 213913 121544 217242 121546
rect 213913 121488 213918 121544
rect 213974 121488 217242 121544
rect 268150 121516 268210 121622
rect 268510 121620 268516 121684
rect 268580 121620 268586 121684
rect 282821 121682 282887 121685
rect 279956 121680 282887 121682
rect 279956 121624 282826 121680
rect 282882 121624 282887 121680
rect 279956 121622 282887 121624
rect 282821 121619 282887 121622
rect 213913 121486 217242 121488
rect 213913 121483 213979 121486
rect 67357 120866 67423 120869
rect 68142 120866 68816 120872
rect 67357 120864 68816 120866
rect 67357 120808 67362 120864
rect 67418 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 231761 121274 231827 121277
rect 228968 121272 231827 121274
rect 228968 121216 231766 121272
rect 231822 121216 231827 121272
rect 228968 121214 231827 121216
rect 231761 121211 231827 121214
rect 264421 121274 264487 121277
rect 268510 121274 268516 121276
rect 264421 121272 268516 121274
rect 264421 121216 264426 121272
rect 264482 121216 268516 121272
rect 264421 121214 268516 121216
rect 264421 121211 264487 121214
rect 268510 121212 268516 121214
rect 268580 121212 268586 121276
rect 214005 120864 217242 120866
rect 67418 120808 68202 120812
rect 67357 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 265985 120866 266051 120869
rect 268150 120866 268210 121108
rect 282821 120866 282887 120869
rect 265985 120864 268210 120866
rect 265985 120808 265990 120864
rect 266046 120808 268210 120864
rect 265985 120806 268210 120808
rect 279956 120864 282887 120866
rect 279956 120808 282826 120864
rect 282882 120808 282887 120864
rect 279956 120806 282887 120808
rect 67357 120803 67423 120806
rect 214005 120803 214071 120806
rect 265985 120803 266051 120806
rect 282821 120803 282887 120806
rect 231301 120730 231367 120733
rect 228968 120728 231367 120730
rect 213913 120186 213979 120189
rect 217182 120186 217242 120700
rect 228968 120672 231306 120728
rect 231362 120672 231367 120728
rect 228968 120670 231367 120672
rect 231301 120667 231367 120670
rect 265893 120458 265959 120461
rect 268150 120458 268210 120700
rect 265893 120456 268210 120458
rect 265893 120400 265898 120456
rect 265954 120400 268210 120456
rect 265893 120398 268210 120400
rect 265893 120395 265959 120398
rect 231485 120322 231551 120325
rect 228968 120320 231551 120322
rect 228968 120264 231490 120320
rect 231546 120264 231551 120320
rect 228968 120262 231551 120264
rect 231485 120259 231551 120262
rect 213913 120184 217242 120186
rect 213913 120128 213918 120184
rect 213974 120128 217242 120184
rect 213913 120126 217242 120128
rect 265801 120186 265867 120189
rect 265801 120184 267842 120186
rect 265801 120128 265806 120184
rect 265862 120128 267842 120184
rect 265801 120126 267842 120128
rect 213913 120123 213979 120126
rect 265801 120123 265867 120126
rect 267782 120050 267842 120126
rect 268334 120050 268394 120292
rect 282729 120186 282795 120189
rect 279956 120184 282795 120186
rect 279956 120128 282734 120184
rect 282790 120128 282795 120184
rect 279956 120126 282795 120128
rect 282729 120123 282795 120126
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 267782 119990 268394 120050
rect 231761 119778 231827 119781
rect 228968 119776 231827 119778
rect 228968 119720 231766 119776
rect 231822 119720 231827 119776
rect 228968 119718 231827 119720
rect 231761 119715 231827 119718
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 214005 119579 214071 119582
rect 265617 119506 265683 119509
rect 268150 119506 268210 119748
rect 265617 119504 268210 119506
rect 173014 119308 173020 119372
rect 173084 119370 173090 119372
rect 204989 119370 205055 119373
rect 173084 119368 205055 119370
rect 173084 119312 204994 119368
rect 205050 119312 205055 119368
rect 173084 119310 205055 119312
rect 173084 119308 173090 119310
rect 204989 119307 205055 119310
rect 213361 119098 213427 119101
rect 217182 119098 217242 119476
rect 265617 119448 265622 119504
rect 265678 119448 268210 119504
rect 265617 119446 268210 119448
rect 265617 119443 265683 119446
rect 231301 119370 231367 119373
rect 282821 119370 282887 119373
rect 228968 119368 231367 119370
rect 228968 119312 231306 119368
rect 231362 119312 231367 119368
rect 279956 119368 282887 119370
rect 228968 119310 231367 119312
rect 231301 119307 231367 119310
rect 213361 119096 217242 119098
rect 213361 119040 213366 119096
rect 213422 119040 217242 119096
rect 213361 119038 217242 119040
rect 264237 119098 264303 119101
rect 268150 119098 268210 119340
rect 279956 119312 282826 119368
rect 282882 119312 282887 119368
rect 279956 119310 282887 119312
rect 282821 119307 282887 119310
rect 264237 119096 268210 119098
rect 264237 119040 264242 119096
rect 264298 119040 268210 119096
rect 264237 119038 268210 119040
rect 213361 119035 213427 119038
rect 264237 119035 264303 119038
rect 213913 118962 213979 118965
rect 230657 118962 230723 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 228968 118960 230723 118962
rect 228968 118904 230662 118960
rect 230718 118904 230723 118960
rect 228968 118902 230723 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 230657 118899 230723 118902
rect 265525 118826 265591 118829
rect 265525 118824 267842 118826
rect 265525 118768 265530 118824
rect 265586 118768 267842 118824
rect 265525 118766 267842 118768
rect 265525 118763 265591 118766
rect 267782 118690 267842 118766
rect 268334 118690 268394 118932
rect 267782 118630 268394 118690
rect 281901 118554 281967 118557
rect 279956 118552 281967 118554
rect 237966 118418 237972 118420
rect 228968 118358 237972 118418
rect 237966 118356 237972 118358
rect 238036 118356 238042 118420
rect 265157 118282 265223 118285
rect 268150 118282 268210 118524
rect 279956 118496 281906 118552
rect 281962 118496 281967 118552
rect 279956 118494 281967 118496
rect 281901 118491 281967 118494
rect 265157 118280 268210 118282
rect 265157 118224 265162 118280
rect 265218 118224 268210 118280
rect 265157 118222 268210 118224
rect 265157 118219 265223 118222
rect 168230 117948 168236 118012
rect 168300 118010 168306 118012
rect 214741 118010 214807 118013
rect 168300 118008 214807 118010
rect 168300 117952 214746 118008
rect 214802 117952 214807 118008
rect 168300 117950 214807 117952
rect 168300 117948 168306 117950
rect 214741 117947 214807 117950
rect 213913 117602 213979 117605
rect 217182 117602 217242 118116
rect 231393 118010 231459 118013
rect 228968 118008 231459 118010
rect 228968 117952 231398 118008
rect 231454 117952 231459 118008
rect 228968 117950 231459 117952
rect 231393 117947 231459 117950
rect 265985 117874 266051 117877
rect 268150 117874 268210 118116
rect 282821 117874 282887 117877
rect 265985 117872 268210 117874
rect 265985 117816 265990 117872
rect 266046 117816 268210 117872
rect 265985 117814 268210 117816
rect 279956 117872 282887 117874
rect 279956 117816 282826 117872
rect 282882 117816 282887 117872
rect 279956 117814 282887 117816
rect 265985 117811 266051 117814
rect 282821 117811 282887 117814
rect 213913 117600 217242 117602
rect 213913 117544 213918 117600
rect 213974 117544 217242 117600
rect 213913 117542 217242 117544
rect 213913 117539 213979 117542
rect 231117 117466 231183 117469
rect 228968 117464 231183 117466
rect 214005 117330 214071 117333
rect 214005 117328 216874 117330
rect 214005 117272 214010 117328
rect 214066 117272 216874 117328
rect 214005 117270 216874 117272
rect 214005 117267 214071 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 228968 117408 231122 117464
rect 231178 117408 231183 117464
rect 228968 117406 231183 117408
rect 231117 117403 231183 117406
rect 265893 117466 265959 117469
rect 268150 117466 268210 117708
rect 265893 117464 268210 117466
rect 265893 117408 265898 117464
rect 265954 117408 268210 117464
rect 265893 117406 268210 117408
rect 265893 117403 265959 117406
rect 264421 117330 264487 117333
rect 268510 117330 268516 117332
rect 264421 117328 268516 117330
rect 264421 117272 264426 117328
rect 264482 117272 268516 117328
rect 264421 117270 268516 117272
rect 264421 117267 264487 117270
rect 268510 117268 268516 117270
rect 268580 117268 268586 117332
rect 216814 117134 217426 117194
rect 230657 117058 230723 117061
rect 228968 117056 230723 117058
rect 228968 117000 230662 117056
rect 230718 117000 230723 117056
rect 228968 116998 230723 117000
rect 230657 116995 230723 116998
rect 265525 116922 265591 116925
rect 268150 116922 268210 117164
rect 282821 117058 282887 117061
rect 279956 117056 282887 117058
rect 279956 117000 282826 117056
rect 282882 117000 282887 117056
rect 279956 116998 282887 117000
rect 282821 116995 282887 116998
rect 265525 116920 268210 116922
rect 265525 116864 265530 116920
rect 265586 116864 268210 116920
rect 265525 116862 268210 116864
rect 265525 116859 265591 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 231485 116514 231551 116517
rect 228968 116512 231551 116514
rect 228968 116456 231490 116512
rect 231546 116456 231551 116512
rect 228968 116454 231551 116456
rect 231485 116451 231551 116454
rect 265617 116514 265683 116517
rect 268150 116514 268210 116756
rect 265617 116512 268210 116514
rect 265617 116456 265622 116512
rect 265678 116456 268210 116512
rect 265617 116454 268210 116456
rect 265617 116451 265683 116454
rect 268510 116452 268516 116516
rect 268580 116452 268586 116516
rect 268518 116348 268578 116452
rect 282177 116378 282243 116381
rect 279956 116376 282243 116378
rect 279956 116320 282182 116376
rect 282238 116320 282243 116376
rect 279956 116318 282243 116320
rect 282177 116315 282243 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 214005 116179 214071 116182
rect 231209 116106 231275 116109
rect 228968 116104 231275 116106
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 228968 116048 231214 116104
rect 231270 116048 231275 116104
rect 228968 116046 231275 116048
rect 231209 116043 231275 116046
rect 266077 116106 266143 116109
rect 266077 116104 268210 116106
rect 266077 116048 266082 116104
rect 266138 116048 268210 116104
rect 266077 116046 268210 116048
rect 266077 116043 266143 116046
rect 268150 115940 268210 116046
rect 216814 115774 217426 115834
rect 240726 115562 240732 115564
rect 228968 115502 240732 115562
rect 240726 115500 240732 115502
rect 240796 115500 240802 115564
rect 282085 115562 282151 115565
rect 279956 115560 282151 115562
rect 213913 115018 213979 115021
rect 217182 115018 217242 115396
rect 265617 115290 265683 115293
rect 268150 115290 268210 115532
rect 279956 115504 282090 115560
rect 282146 115504 282151 115560
rect 279956 115502 282151 115504
rect 282085 115499 282151 115502
rect 265617 115288 268210 115290
rect 265617 115232 265622 115288
rect 265678 115232 268210 115288
rect 265617 115230 268210 115232
rect 265617 115227 265683 115230
rect 231209 115154 231275 115157
rect 228968 115152 231275 115154
rect 228968 115096 231214 115152
rect 231270 115096 231275 115152
rect 228968 115094 231275 115096
rect 231209 115091 231275 115094
rect 213913 115016 217242 115018
rect 213913 114960 213918 115016
rect 213974 114960 217242 115016
rect 213913 114958 217242 114960
rect 213913 114955 213979 114958
rect 265433 114882 265499 114885
rect 268150 114882 268210 115124
rect 265433 114880 268210 114882
rect 213453 114610 213519 114613
rect 217182 114610 217242 114852
rect 265433 114824 265438 114880
rect 265494 114824 268210 114880
rect 265433 114822 268210 114824
rect 265433 114819 265499 114822
rect 281717 114746 281783 114749
rect 258030 114686 268210 114746
rect 279956 114744 281783 114746
rect 279956 114688 281722 114744
rect 281778 114688 281783 114744
rect 279956 114686 281783 114688
rect 231117 114610 231183 114613
rect 213453 114608 217242 114610
rect 213453 114552 213458 114608
rect 213514 114552 217242 114608
rect 213453 114550 217242 114552
rect 228968 114608 231183 114610
rect 228968 114552 231122 114608
rect 231178 114552 231183 114608
rect 228968 114550 231183 114552
rect 213453 114547 213519 114550
rect 231117 114547 231183 114550
rect 254526 114548 254532 114612
rect 254596 114610 254602 114612
rect 258030 114610 258090 114686
rect 254596 114550 258090 114610
rect 268150 114580 268210 114686
rect 281717 114683 281783 114686
rect 254596 114548 254602 114550
rect 231761 114202 231827 114205
rect 228968 114200 231827 114202
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 228968 114144 231766 114200
rect 231822 114144 231827 114200
rect 228968 114142 231827 114144
rect 231761 114139 231827 114142
rect 265525 113930 265591 113933
rect 268150 113930 268210 114172
rect 282269 114066 282335 114069
rect 279956 114064 282335 114066
rect 279956 114008 282274 114064
rect 282330 114008 282335 114064
rect 279956 114006 282335 114008
rect 282269 114003 282335 114006
rect 265525 113928 268210 113930
rect 265525 113872 265530 113928
rect 265586 113872 268210 113928
rect 265525 113870 268210 113872
rect 265525 113867 265591 113870
rect 231301 113658 231367 113661
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 228968 113656 231367 113658
rect 228968 113600 231306 113656
rect 231362 113600 231367 113656
rect 228968 113598 231367 113600
rect 214005 113595 214071 113598
rect 231301 113595 231367 113598
rect 265433 113522 265499 113525
rect 268150 113522 268210 113764
rect 265433 113520 268210 113522
rect 213913 113250 213979 113253
rect 217366 113250 217426 113492
rect 265433 113464 265438 113520
rect 265494 113464 268210 113520
rect 265433 113462 268210 113464
rect 265433 113459 265499 113462
rect 231485 113250 231551 113253
rect 213913 113248 217426 113250
rect 213913 113192 213918 113248
rect 213974 113192 217426 113248
rect 213913 113190 217426 113192
rect 228968 113248 231551 113250
rect 228968 113192 231490 113248
rect 231546 113192 231551 113248
rect 228968 113190 231551 113192
rect 213913 113187 213979 113190
rect 231485 113187 231551 113190
rect 265893 113250 265959 113253
rect 265893 113248 267842 113250
rect 265893 113192 265898 113248
rect 265954 113192 267842 113248
rect 265893 113190 267842 113192
rect 265893 113187 265959 113190
rect 267782 113114 267842 113190
rect 268334 113114 268394 113356
rect 282637 113250 282703 113253
rect 279956 113248 282703 113250
rect 279956 113192 282642 113248
rect 282698 113192 282703 113248
rect 279956 113190 282703 113192
rect 282637 113187 282703 113190
rect 267782 113054 268394 113114
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 231669 112706 231735 112709
rect 228968 112704 231735 112706
rect 228968 112648 231674 112704
rect 231730 112648 231735 112704
rect 228968 112646 231735 112648
rect 231669 112643 231735 112646
rect 265525 112706 265591 112709
rect 268150 112706 268210 112948
rect 582649 112842 582715 112845
rect 583520 112842 584960 112932
rect 582649 112840 584960 112842
rect 582649 112784 582654 112840
rect 582710 112784 584960 112840
rect 582649 112782 584960 112784
rect 582649 112779 582715 112782
rect 265525 112704 268210 112706
rect 265525 112648 265530 112704
rect 265586 112648 268210 112704
rect 583520 112692 584960 112782
rect 265525 112646 268210 112648
rect 265525 112643 265591 112646
rect 231761 112298 231827 112301
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 228968 112296 231827 112298
rect 228968 112240 231766 112296
rect 231822 112240 231827 112296
rect 228968 112238 231827 112240
rect 214005 112235 214071 112238
rect 231761 112235 231827 112238
rect 265617 112298 265683 112301
rect 268150 112298 268210 112540
rect 282085 112434 282151 112437
rect 279956 112432 282151 112434
rect 279956 112376 282090 112432
rect 282146 112376 282151 112432
rect 279956 112374 282151 112376
rect 282085 112371 282151 112374
rect 265617 112296 268210 112298
rect 265617 112240 265622 112296
rect 265678 112240 268210 112296
rect 265617 112238 268210 112240
rect 265617 112235 265683 112238
rect 265893 112162 265959 112165
rect 265893 112160 268210 112162
rect 213913 111890 213979 111893
rect 217182 111890 217242 112132
rect 265893 112104 265898 112160
rect 265954 112104 268210 112160
rect 265893 112102 268210 112104
rect 265893 112099 265959 112102
rect 268150 111996 268210 112102
rect 213913 111888 217242 111890
rect 213913 111832 213918 111888
rect 213974 111832 217242 111888
rect 213913 111830 217242 111832
rect 213913 111827 213979 111830
rect 168281 111754 168347 111757
rect 231669 111754 231735 111757
rect 164694 111752 168347 111754
rect 164694 111696 168286 111752
rect 168342 111696 168347 111752
rect 164694 111694 168347 111696
rect 228968 111752 231735 111754
rect 228968 111696 231674 111752
rect 231730 111696 231735 111752
rect 228968 111694 231735 111696
rect 168281 111691 168347 111694
rect 231669 111691 231735 111694
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 231761 111346 231827 111349
rect 228968 111344 231827 111346
rect 228968 111288 231766 111344
rect 231822 111288 231827 111344
rect 228968 111286 231827 111288
rect 231761 111283 231827 111286
rect 264421 111346 264487 111349
rect 268150 111346 268210 111588
rect 264421 111344 268210 111346
rect 264421 111288 264426 111344
rect 264482 111288 268210 111344
rect 264421 111286 268210 111288
rect 264421 111283 264487 111286
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 265157 110938 265223 110941
rect 268150 110938 268210 111180
rect 279926 111074 279986 111724
rect 279926 111014 287070 111074
rect 282821 110938 282887 110941
rect 265157 110936 268210 110938
rect 265157 110880 265162 110936
rect 265218 110880 268210 110936
rect 265157 110878 268210 110880
rect 279956 110936 282887 110938
rect 279956 110880 282826 110936
rect 282882 110880 282887 110936
rect 279956 110878 282887 110880
rect 214005 110875 214071 110878
rect 265157 110875 265223 110878
rect 282821 110875 282887 110878
rect 230933 110802 230999 110805
rect 228968 110800 230999 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217182 110530 217242 110772
rect 228968 110744 230938 110800
rect 230994 110744 230999 110800
rect 228968 110742 230999 110744
rect 230933 110739 230999 110742
rect 213913 110528 217242 110530
rect 213913 110472 213918 110528
rect 213974 110472 217242 110528
rect 213913 110470 217242 110472
rect 265893 110530 265959 110533
rect 268334 110530 268394 110772
rect 265893 110528 268394 110530
rect 265893 110472 265898 110528
rect 265954 110472 268394 110528
rect 265893 110470 268394 110472
rect 287010 110530 287070 111014
rect 294270 110530 294276 110532
rect 287010 110470 294276 110530
rect 213913 110467 213979 110470
rect 265893 110467 265959 110470
rect 294270 110468 294276 110470
rect 294340 110468 294346 110532
rect 231761 110394 231827 110397
rect 228968 110392 231827 110394
rect 228968 110336 231766 110392
rect 231822 110336 231827 110392
rect 228968 110334 231827 110336
rect 231761 110331 231827 110334
rect 168189 110122 168255 110125
rect 164694 110120 168255 110122
rect 164694 110064 168194 110120
rect 168250 110064 168255 110120
rect 164694 110062 168255 110064
rect 168189 110059 168255 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 265525 110122 265591 110125
rect 268150 110122 268210 110364
rect 265525 110120 268210 110122
rect 265525 110064 265530 110120
rect 265586 110064 268210 110120
rect 265525 110062 268210 110064
rect 265525 110059 265591 110062
rect 231669 109850 231735 109853
rect 228968 109848 231735 109850
rect 228968 109792 231674 109848
rect 231730 109792 231735 109848
rect 228968 109790 231735 109792
rect 231669 109787 231735 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 265985 109714 266051 109717
rect 268150 109714 268210 109956
rect 265985 109712 268210 109714
rect 265985 109656 265990 109712
rect 266046 109656 268210 109712
rect 265985 109654 268210 109656
rect 214005 109651 214071 109654
rect 265985 109651 266051 109654
rect 279926 109578 279986 110092
rect 213913 109170 213979 109173
rect 217182 109170 217242 109548
rect 231669 109442 231735 109445
rect 228968 109440 231735 109442
rect 228968 109384 231674 109440
rect 231730 109384 231735 109440
rect 228968 109382 231735 109384
rect 231669 109379 231735 109382
rect 213913 109168 217242 109170
rect 213913 109112 213918 109168
rect 213974 109112 217242 109168
rect 213913 109110 217242 109112
rect 265893 109170 265959 109173
rect 268150 109170 268210 109548
rect 279926 109518 287070 109578
rect 282821 109442 282887 109445
rect 279956 109440 282887 109442
rect 279956 109384 282826 109440
rect 282882 109384 282887 109440
rect 279956 109382 282887 109384
rect 282821 109379 282887 109382
rect 265893 109168 268210 109170
rect 265893 109112 265898 109168
rect 265954 109112 268210 109168
rect 265893 109110 268210 109112
rect 287010 109170 287070 109518
rect 290590 109170 290596 109172
rect 287010 109110 290596 109170
rect 213913 109107 213979 109110
rect 265893 109107 265959 109110
rect 290590 109108 290596 109110
rect 290660 109108 290666 109172
rect 231761 108898 231827 108901
rect 228968 108896 231827 108898
rect 167913 108762 167979 108765
rect 164694 108760 167979 108762
rect 164694 108704 167918 108760
rect 167974 108704 167979 108760
rect 164694 108702 167979 108704
rect 167913 108699 167979 108702
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 228968 108840 231766 108896
rect 231822 108840 231827 108896
rect 228968 108838 231827 108840
rect 231761 108835 231827 108838
rect 265985 108762 266051 108765
rect 268150 108762 268210 109004
rect 265985 108760 268210 108762
rect 265985 108704 265990 108760
rect 266046 108704 268210 108760
rect 265985 108702 268210 108704
rect 265985 108699 266051 108702
rect 282821 108626 282887 108629
rect 279956 108624 282887 108626
rect 231669 108490 231735 108493
rect 228968 108488 231735 108490
rect 228968 108432 231674 108488
rect 231730 108432 231735 108488
rect 228968 108430 231735 108432
rect 231669 108427 231735 108430
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 265341 108354 265407 108357
rect 268150 108354 268210 108596
rect 279956 108568 282826 108624
rect 282882 108568 282887 108624
rect 279956 108566 282887 108568
rect 282821 108563 282887 108566
rect 265341 108352 268210 108354
rect 265341 108296 265346 108352
rect 265402 108296 268210 108352
rect 265341 108294 268210 108296
rect 214005 108291 214071 108294
rect 265341 108291 265407 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 230565 107946 230631 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 228968 107944 230631 107946
rect 228968 107888 230570 107944
rect 230626 107888 230631 107944
rect 228968 107886 230631 107888
rect 213913 107883 213979 107886
rect 230565 107883 230631 107886
rect 265893 107946 265959 107949
rect 268518 107948 268578 108188
rect 265893 107944 268210 107946
rect 265893 107888 265898 107944
rect 265954 107888 268210 107944
rect 265893 107886 268210 107888
rect 265893 107883 265959 107886
rect 268150 107780 268210 107886
rect 268510 107884 268516 107948
rect 268580 107884 268586 107948
rect 280245 107810 280311 107813
rect 279956 107808 280311 107810
rect 279956 107752 280250 107808
rect 280306 107752 280311 107808
rect 279956 107750 280311 107752
rect 280245 107747 280311 107750
rect 231761 107538 231827 107541
rect 228968 107536 231827 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 228968 107480 231766 107536
rect 231822 107480 231827 107536
rect 228968 107478 231827 107480
rect 231761 107475 231827 107478
rect 264513 107538 264579 107541
rect 268510 107538 268516 107540
rect 264513 107536 268516 107538
rect 264513 107480 264518 107536
rect 264574 107480 268516 107536
rect 264513 107478 268516 107480
rect 264513 107475 264579 107478
rect 268510 107476 268516 107478
rect 268580 107476 268586 107540
rect 231485 107130 231551 107133
rect 228968 107128 231551 107130
rect 228968 107072 231490 107128
rect 231546 107072 231551 107128
rect 228968 107070 231551 107072
rect 231485 107067 231551 107070
rect 264513 107130 264579 107133
rect 268150 107130 268210 107372
rect 264513 107128 268210 107130
rect 264513 107072 264518 107128
rect 264574 107072 268210 107128
rect 264513 107070 268210 107072
rect 264513 107067 264579 107070
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 214005 106931 214071 106934
rect 213913 106586 213979 106589
rect 217182 106586 217242 106828
rect 265985 106722 266051 106725
rect 268150 106722 268210 106964
rect 265985 106720 268210 106722
rect 265985 106664 265990 106720
rect 266046 106664 268210 106720
rect 265985 106662 268210 106664
rect 265985 106659 266051 106662
rect 230749 106586 230815 106589
rect 213913 106584 217242 106586
rect 213913 106528 213918 106584
rect 213974 106528 217242 106584
rect 213913 106526 217242 106528
rect 228968 106584 230815 106586
rect 228968 106528 230754 106584
rect 230810 106528 230815 106584
rect 228968 106526 230815 106528
rect 213913 106523 213979 106526
rect 230749 106523 230815 106526
rect 265893 106586 265959 106589
rect 265893 106584 268210 106586
rect 265893 106528 265898 106584
rect 265954 106528 268210 106584
rect 265893 106526 268210 106528
rect 265893 106523 265959 106526
rect 268150 106420 268210 106526
rect 279926 106450 279986 107100
rect 287094 106450 287100 106452
rect 279926 106390 287100 106450
rect 287094 106388 287100 106390
rect 287164 106388 287170 106452
rect 285622 106314 285628 106316
rect 279956 106254 285628 106314
rect 285622 106252 285628 106254
rect 285692 106252 285698 106316
rect 233918 106178 233924 106180
rect 213913 105770 213979 105773
rect 217182 105770 217242 106148
rect 228968 106118 233924 106178
rect 233918 106116 233924 106118
rect 233988 106116 233994 106180
rect 213913 105768 217242 105770
rect 213913 105712 213918 105768
rect 213974 105712 217242 105768
rect 213913 105710 217242 105712
rect 265249 105770 265315 105773
rect 268150 105770 268210 106012
rect 265249 105768 268210 105770
rect 265249 105712 265254 105768
rect 265310 105712 268210 105768
rect 265249 105710 268210 105712
rect 213913 105707 213979 105710
rect 265249 105707 265315 105710
rect 231761 105634 231827 105637
rect 228968 105632 231827 105634
rect 214414 105300 214420 105364
rect 214484 105362 214490 105364
rect 217182 105362 217242 105604
rect 228968 105576 231766 105632
rect 231822 105576 231827 105632
rect 228968 105574 231827 105576
rect 231761 105571 231827 105574
rect 214484 105302 217242 105362
rect 265893 105362 265959 105365
rect 268150 105362 268210 105604
rect 282821 105498 282887 105501
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 282821 105435 282887 105438
rect 265893 105360 268210 105362
rect 265893 105304 265898 105360
rect 265954 105304 268210 105360
rect 265893 105302 268210 105304
rect 214484 105300 214490 105302
rect 265893 105299 265959 105302
rect 214005 105226 214071 105229
rect 231485 105226 231551 105229
rect 214005 105224 217426 105226
rect 214005 105168 214010 105224
rect 214066 105168 217426 105224
rect 214005 105166 217426 105168
rect 228968 105224 231551 105226
rect 228968 105168 231490 105224
rect 231546 105168 231551 105224
rect 228968 105166 231551 105168
rect 214005 105163 214071 105166
rect 217366 104924 217426 105166
rect 231485 105163 231551 105166
rect 265617 104954 265683 104957
rect 268150 104954 268210 105196
rect 265617 104952 268210 104954
rect 265617 104896 265622 104952
rect 265678 104896 268210 104952
rect 265617 104894 268210 104896
rect 265617 104891 265683 104894
rect 281717 104818 281783 104821
rect 279956 104816 281783 104818
rect 231393 104682 231459 104685
rect 228968 104680 231459 104682
rect 228968 104624 231398 104680
rect 231454 104624 231459 104680
rect 228968 104622 231459 104624
rect 231393 104619 231459 104622
rect 265617 104546 265683 104549
rect 268150 104546 268210 104788
rect 279956 104760 281722 104816
rect 281778 104760 281783 104816
rect 279956 104758 281783 104760
rect 281717 104755 281783 104758
rect 265617 104544 268210 104546
rect 265617 104488 265622 104544
rect 265678 104488 268210 104544
rect 265617 104486 268210 104488
rect 265617 104483 265683 104486
rect 230565 104274 230631 104277
rect 228968 104272 230631 104274
rect 214649 103866 214715 103869
rect 217182 103866 217242 104244
rect 228968 104216 230570 104272
rect 230626 104216 230631 104272
rect 228968 104214 230631 104216
rect 230565 104211 230631 104214
rect 265985 104002 266051 104005
rect 268150 104002 268210 104380
rect 280245 104002 280311 104005
rect 265985 104000 268210 104002
rect 265985 103944 265990 104000
rect 266046 103944 268210 104000
rect 265985 103942 268210 103944
rect 279956 104000 280311 104002
rect 279956 103944 280250 104000
rect 280306 103944 280311 104000
rect 279956 103942 280311 103944
rect 265985 103939 266051 103942
rect 280245 103939 280311 103942
rect 214649 103864 217242 103866
rect 214649 103808 214654 103864
rect 214710 103808 217242 103864
rect 214649 103806 217242 103808
rect 214649 103803 214715 103806
rect 213913 103730 213979 103733
rect 231577 103730 231643 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 228968 103728 231643 103730
rect 228968 103672 231582 103728
rect 231638 103672 231643 103728
rect 228968 103670 231643 103672
rect 213913 103667 213979 103670
rect 217182 103564 217242 103670
rect 231577 103667 231643 103670
rect 265893 103594 265959 103597
rect 268150 103594 268210 103836
rect 265893 103592 268210 103594
rect 265893 103536 265898 103592
rect 265954 103536 268210 103592
rect 265893 103534 268210 103536
rect 265893 103531 265959 103534
rect 231117 103322 231183 103325
rect 228968 103320 231183 103322
rect 228968 103264 231122 103320
rect 231178 103264 231183 103320
rect 228968 103262 231183 103264
rect 231117 103259 231183 103262
rect 265525 103186 265591 103189
rect 268150 103186 268210 103428
rect 285806 103186 285812 103188
rect 265525 103184 268210 103186
rect 265525 103128 265530 103184
rect 265586 103128 268210 103184
rect 265525 103126 268210 103128
rect 279956 103126 285812 103186
rect 265525 103123 265591 103126
rect 285806 103124 285812 103126
rect 285876 103124 285882 103188
rect 213913 102506 213979 102509
rect 217182 102506 217242 102884
rect 230473 102778 230539 102781
rect 228968 102776 230539 102778
rect 228968 102720 230478 102776
rect 230534 102720 230539 102776
rect 228968 102718 230539 102720
rect 230473 102715 230539 102718
rect 265617 102778 265683 102781
rect 268150 102778 268210 103020
rect 265617 102776 268210 102778
rect 265617 102720 265622 102776
rect 265678 102720 268210 102776
rect 265617 102718 268210 102720
rect 265617 102715 265683 102718
rect 213913 102504 217242 102506
rect 213913 102448 213918 102504
rect 213974 102448 217242 102504
rect 213913 102446 217242 102448
rect 213913 102443 213979 102446
rect 67633 102370 67699 102373
rect 68142 102370 68816 102376
rect 230422 102370 230428 102372
rect 67633 102368 68816 102370
rect 67633 102312 67638 102368
rect 67694 102316 68816 102368
rect 67694 102312 68202 102316
rect 67633 102310 68202 102312
rect 200070 102310 217242 102370
rect 228968 102310 230428 102370
rect 67633 102307 67699 102310
rect 172094 102172 172100 102236
rect 172164 102234 172170 102236
rect 200070 102234 200130 102310
rect 172164 102174 200130 102234
rect 217182 102204 217242 102310
rect 230422 102308 230428 102310
rect 230492 102308 230498 102372
rect 265341 102370 265407 102373
rect 268518 102372 268578 102612
rect 281625 102506 281691 102509
rect 279956 102504 281691 102506
rect 279956 102448 281630 102504
rect 281686 102448 281691 102504
rect 279956 102446 281691 102448
rect 281625 102443 281691 102446
rect 265341 102368 268210 102370
rect 265341 102312 265346 102368
rect 265402 102312 268210 102368
rect 265341 102310 268210 102312
rect 265341 102307 265407 102310
rect 233734 102234 233740 102236
rect 231350 102174 233740 102234
rect 172164 102172 172170 102174
rect 231350 101826 231410 102174
rect 233734 102172 233740 102174
rect 233804 102172 233810 102236
rect 268150 102204 268210 102310
rect 268510 102308 268516 102372
rect 268580 102308 268586 102372
rect 264329 101962 264395 101965
rect 264329 101960 268210 101962
rect 264329 101904 264334 101960
rect 264390 101904 268210 101960
rect 264329 101902 268210 101904
rect 264329 101899 264395 101902
rect 228968 101766 231410 101826
rect 268150 101796 268210 101902
rect 265985 101554 266051 101557
rect 265985 101552 268394 101554
rect 214005 101146 214071 101149
rect 217182 101146 217242 101524
rect 265985 101496 265990 101552
rect 266046 101496 268394 101552
rect 265985 101494 268394 101496
rect 265985 101491 266051 101494
rect 230749 101418 230815 101421
rect 228968 101416 230815 101418
rect 228968 101360 230754 101416
rect 230810 101360 230815 101416
rect 228968 101358 230815 101360
rect 230749 101355 230815 101358
rect 268334 101252 268394 101494
rect 214005 101144 217242 101146
rect 214005 101088 214010 101144
rect 214066 101088 217242 101144
rect 214005 101086 217242 101088
rect 214005 101083 214071 101086
rect 265893 101010 265959 101013
rect 279926 101010 279986 101660
rect 291326 101010 291332 101012
rect 265893 101008 268210 101010
rect 213913 100874 213979 100877
rect 213913 100872 216874 100874
rect 213913 100816 213918 100872
rect 213974 100816 216874 100872
rect 213913 100814 216874 100816
rect 213913 100811 213979 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 216814 100738 216874 100814
rect 217366 100738 217426 100980
rect 265893 100952 265898 101008
rect 265954 100952 268210 101008
rect 265893 100950 268210 100952
rect 279926 100950 291332 101010
rect 265893 100947 265959 100950
rect 230565 100874 230631 100877
rect 228968 100872 230631 100874
rect 228968 100816 230570 100872
rect 230626 100816 230631 100872
rect 268150 100844 268210 100950
rect 291326 100948 291332 100950
rect 291396 100948 291402 101012
rect 280153 100874 280219 100877
rect 279956 100872 280219 100874
rect 228968 100814 230631 100816
rect 279956 100816 280158 100872
rect 280214 100816 280219 100872
rect 279956 100814 280219 100816
rect 230565 100811 230631 100814
rect 280153 100811 280219 100814
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 216814 100678 217426 100738
rect 67725 100675 67791 100678
rect 261569 100602 261635 100605
rect 268510 100602 268516 100604
rect 261569 100600 268516 100602
rect 261569 100544 261574 100600
rect 261630 100544 268516 100600
rect 261569 100542 268516 100544
rect 261569 100539 261635 100542
rect 268510 100540 268516 100542
rect 268580 100540 268586 100604
rect 231669 100466 231735 100469
rect 228968 100464 231735 100466
rect 228968 100408 231674 100464
rect 231730 100408 231735 100464
rect 228968 100406 231735 100408
rect 231669 100403 231735 100406
rect 213913 99786 213979 99789
rect 217182 99786 217242 100300
rect 265893 100194 265959 100197
rect 268150 100194 268210 100436
rect 281533 100194 281599 100197
rect 265893 100192 268210 100194
rect 265893 100136 265898 100192
rect 265954 100136 268210 100192
rect 265893 100134 268210 100136
rect 279956 100192 281599 100194
rect 279956 100136 281538 100192
rect 281594 100136 281599 100192
rect 279956 100134 281599 100136
rect 265893 100131 265959 100134
rect 281533 100131 281599 100134
rect 231485 99922 231551 99925
rect 228968 99920 231551 99922
rect 228968 99864 231490 99920
rect 231546 99864 231551 99920
rect 228968 99862 231551 99864
rect 231485 99859 231551 99862
rect 213913 99784 217242 99786
rect 213913 99728 213918 99784
rect 213974 99728 217242 99784
rect 213913 99726 217242 99728
rect 265157 99786 265223 99789
rect 268150 99786 268210 100028
rect 265157 99784 268210 99786
rect 265157 99728 265162 99784
rect 265218 99728 268210 99784
rect 265157 99726 268210 99728
rect 213913 99723 213979 99726
rect 265157 99723 265223 99726
rect 214833 99514 214899 99517
rect 214833 99512 216874 99514
rect 214833 99456 214838 99512
rect 214894 99456 216874 99512
rect 214833 99454 216874 99456
rect 214833 99451 214899 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 231761 99514 231827 99517
rect 228968 99512 231827 99514
rect 228968 99456 231766 99512
rect 231822 99456 231827 99512
rect 228968 99454 231827 99456
rect 231761 99451 231827 99454
rect 265617 99514 265683 99517
rect 265617 99512 267842 99514
rect 265617 99456 265622 99512
rect 265678 99456 267842 99512
rect 265617 99454 267842 99456
rect 265617 99451 265683 99454
rect 216814 99318 217426 99378
rect 267782 99378 267842 99454
rect 268334 99378 268394 99620
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 281574 99378 281580 99380
rect 267782 99318 268394 99378
rect 279956 99318 281580 99378
rect 281574 99316 281580 99318
rect 281644 99316 281650 99380
rect 583520 99364 584960 99454
rect 231761 99106 231827 99109
rect 229142 99104 231827 99106
rect 229142 99048 231766 99104
rect 231822 99048 231827 99104
rect 229142 99046 231827 99048
rect 229142 98970 229202 99046
rect 231761 99043 231827 99046
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 228968 98910 229202 98970
rect 229318 98908 229324 98972
rect 229388 98970 229394 98972
rect 261201 98970 261267 98973
rect 268334 98970 268394 99212
rect 229388 98910 258090 98970
rect 229388 98908 229394 98910
rect 231485 98562 231551 98565
rect 228968 98560 231551 98562
rect 228968 98504 231490 98560
rect 231546 98504 231551 98560
rect 228968 98502 231551 98504
rect 231485 98499 231551 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 258030 98426 258090 98910
rect 261201 98968 268394 98970
rect 261201 98912 261206 98968
rect 261262 98912 268394 98968
rect 261201 98910 268394 98912
rect 261201 98907 261267 98910
rect 264605 98834 264671 98837
rect 264605 98832 268210 98834
rect 264605 98776 264610 98832
rect 264666 98776 268210 98832
rect 264605 98774 268210 98776
rect 264605 98771 264671 98774
rect 268150 98668 268210 98774
rect 258030 98366 268210 98426
rect 214005 98363 214071 98366
rect 268150 98260 268210 98366
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 230933 98018 230999 98021
rect 279374 98020 279434 98532
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 228968 98016 230999 98018
rect 228968 97960 230938 98016
rect 230994 97960 230999 98016
rect 228968 97958 230999 97960
rect 213913 97955 213979 97958
rect 230933 97955 230999 97958
rect 265750 97956 265756 98020
rect 265820 98018 265826 98020
rect 268510 98018 268516 98020
rect 265820 97958 268516 98018
rect 265820 97956 265826 97958
rect 268510 97956 268516 97958
rect 268580 97956 268586 98020
rect 279366 97956 279372 98020
rect 279436 97956 279442 98020
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect 231577 97610 231643 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 228968 97608 231643 97610
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 216213 97066 216279 97069
rect 217182 97066 217242 97580
rect 228968 97552 231582 97608
rect 231638 97552 231643 97608
rect 228968 97550 231643 97552
rect 231577 97547 231643 97550
rect 265617 97610 265683 97613
rect 268150 97610 268210 97852
rect 265617 97608 268210 97610
rect 265617 97552 265622 97608
rect 265678 97552 268210 97608
rect 265617 97550 268210 97552
rect 265617 97547 265683 97550
rect 265341 97202 265407 97205
rect 268150 97202 268210 97444
rect 279374 97341 279434 97852
rect 279374 97336 279483 97341
rect 279374 97280 279422 97336
rect 279478 97280 279483 97336
rect 279374 97278 279483 97280
rect 279417 97275 279483 97278
rect 265341 97200 268210 97202
rect 265341 97144 265346 97200
rect 265402 97144 268210 97200
rect 265341 97142 268210 97144
rect 265341 97139 265407 97142
rect 268510 97140 268516 97204
rect 268580 97140 268586 97204
rect 229134 97066 229140 97068
rect 216213 97064 217242 97066
rect 216213 97008 216218 97064
rect 216274 97008 217242 97064
rect 216213 97006 217242 97008
rect 228968 97006 229140 97066
rect 216213 97003 216279 97006
rect 229134 97004 229140 97006
rect 229204 97066 229210 97068
rect 231761 97066 231827 97069
rect 229204 97064 231827 97066
rect 229204 97008 231766 97064
rect 231822 97008 231827 97064
rect 268518 97036 268578 97140
rect 229204 97006 231827 97008
rect 229204 97004 229210 97006
rect 231761 97003 231827 97006
rect 214741 96658 214807 96661
rect 217182 96658 217242 96900
rect 265985 96794 266051 96797
rect 265985 96792 268210 96794
rect 265985 96736 265990 96792
rect 266046 96736 268210 96792
rect 265985 96734 268210 96736
rect 265985 96731 266051 96734
rect 229093 96658 229159 96661
rect 214741 96656 217242 96658
rect 214741 96600 214746 96656
rect 214802 96600 217242 96656
rect 214741 96598 217242 96600
rect 228968 96656 229159 96658
rect 228968 96600 229098 96656
rect 229154 96600 229159 96656
rect 268150 96628 268210 96734
rect 279374 96661 279434 97036
rect 279325 96656 279434 96661
rect 228968 96598 229159 96600
rect 214741 96595 214807 96598
rect 229093 96595 229159 96598
rect 279325 96600 279330 96656
rect 279386 96600 279434 96656
rect 279325 96598 279434 96600
rect 279325 96595 279391 96598
rect 216673 95842 216739 95845
rect 217182 95842 217242 96356
rect 216673 95840 217242 95842
rect 216673 95784 216678 95840
rect 216734 95784 217242 95840
rect 216673 95782 217242 95784
rect 216673 95779 216739 95782
rect 228774 95706 228834 96220
rect 230473 95706 230539 95709
rect 228774 95704 230539 95706
rect 228774 95648 230478 95704
rect 230534 95648 230539 95704
rect 228774 95646 230539 95648
rect 230473 95643 230539 95646
rect 265525 95706 265591 95709
rect 268150 95706 268210 96220
rect 265525 95704 268210 95706
rect 265525 95648 265530 95704
rect 265586 95648 268210 95704
rect 265525 95646 268210 95648
rect 265525 95643 265591 95646
rect 227662 95372 227668 95436
rect 227732 95434 227738 95436
rect 228950 95434 228956 95436
rect 227732 95374 228956 95434
rect 227732 95372 227738 95374
rect 228950 95372 228956 95374
rect 229020 95372 229026 95436
rect 250294 95372 250300 95436
rect 250364 95434 250370 95436
rect 279374 95434 279434 96356
rect 250364 95374 279434 95434
rect 250364 95372 250370 95374
rect 178677 95162 178743 95165
rect 279325 95162 279391 95165
rect 178677 95160 279391 95162
rect 178677 95104 178682 95160
rect 178738 95104 279330 95160
rect 279386 95104 279391 95160
rect 178677 95102 279391 95104
rect 178677 95099 178743 95102
rect 279325 95099 279391 95102
rect 185577 95026 185643 95029
rect 279366 95026 279372 95028
rect 185577 95024 279372 95026
rect 185577 94968 185582 95024
rect 185638 94968 279372 95024
rect 185577 94966 279372 94968
rect 185577 94963 185643 94966
rect 279366 94964 279372 94966
rect 279436 94964 279442 95028
rect 66161 94890 66227 94893
rect 210601 94890 210667 94893
rect 66161 94888 210667 94890
rect 66161 94832 66166 94888
rect 66222 94832 210606 94888
rect 210662 94832 210667 94888
rect 66161 94830 210667 94832
rect 66161 94827 66227 94830
rect 210601 94827 210667 94830
rect 94957 94756 95023 94757
rect 104341 94756 104407 94757
rect 94912 94692 94918 94756
rect 94982 94754 95023 94756
rect 94982 94752 95074 94754
rect 95018 94696 95074 94752
rect 94982 94694 95074 94696
rect 94982 94692 95023 94694
rect 104296 94692 104302 94756
rect 104366 94754 104407 94756
rect 116669 94756 116735 94757
rect 120625 94756 120691 94757
rect 133137 94756 133203 94757
rect 151721 94756 151787 94757
rect 116669 94754 116678 94756
rect 104366 94752 104458 94754
rect 104402 94696 104458 94752
rect 104366 94694 104458 94696
rect 116586 94752 116678 94754
rect 116586 94696 116674 94752
rect 116586 94694 116678 94696
rect 104366 94692 104407 94694
rect 94957 94691 95023 94692
rect 104341 94691 104407 94692
rect 116669 94692 116678 94694
rect 116742 94692 116748 94756
rect 120616 94692 120622 94756
rect 120686 94754 120692 94756
rect 120686 94694 120778 94754
rect 120686 94692 120692 94694
rect 133128 94692 133134 94756
rect 133198 94754 133204 94756
rect 151721 94754 151766 94756
rect 133198 94694 133290 94754
rect 151674 94752 151766 94754
rect 151674 94696 151726 94752
rect 151674 94694 151766 94696
rect 133198 94692 133204 94694
rect 151721 94692 151766 94694
rect 151830 94692 151836 94756
rect 116669 94691 116735 94692
rect 120625 94691 120691 94692
rect 133137 94691 133203 94692
rect 151721 94691 151787 94692
rect 67449 93802 67515 93805
rect 214414 93802 214420 93804
rect 67449 93800 214420 93802
rect 67449 93744 67454 93800
rect 67510 93744 214420 93800
rect 67449 93742 214420 93744
rect 67449 93739 67515 93742
rect 214414 93740 214420 93742
rect 214484 93740 214490 93804
rect 60641 93666 60707 93669
rect 206461 93666 206527 93669
rect 60641 93664 206527 93666
rect 60641 93608 60646 93664
rect 60702 93608 206466 93664
rect 206522 93608 206527 93664
rect 60641 93606 206527 93608
rect 60641 93603 60707 93606
rect 206461 93603 206527 93606
rect 85665 93532 85731 93533
rect 107745 93532 107811 93533
rect 115841 93532 115907 93533
rect 122097 93532 122163 93533
rect 85614 93530 85620 93532
rect 85574 93470 85620 93530
rect 85684 93528 85731 93532
rect 107694 93530 107700 93532
rect 85726 93472 85731 93528
rect 85614 93468 85620 93470
rect 85684 93468 85731 93472
rect 107654 93470 107700 93530
rect 107764 93528 107811 93532
rect 115790 93530 115796 93532
rect 107806 93472 107811 93528
rect 107694 93468 107700 93470
rect 107764 93468 107811 93472
rect 115750 93470 115796 93530
rect 115860 93528 115907 93532
rect 122046 93530 122052 93532
rect 115902 93472 115907 93528
rect 115790 93468 115796 93470
rect 115860 93468 115907 93472
rect 122006 93470 122052 93530
rect 122116 93528 122163 93532
rect 122158 93472 122163 93528
rect 122046 93468 122052 93470
rect 122116 93468 122163 93472
rect 85665 93467 85731 93468
rect 107745 93467 107811 93468
rect 115841 93467 115907 93468
rect 122097 93467 122163 93468
rect 196709 93530 196775 93533
rect 281574 93530 281580 93532
rect 196709 93528 281580 93530
rect 196709 93472 196714 93528
rect 196770 93472 281580 93528
rect 196709 93470 281580 93472
rect 196709 93467 196775 93470
rect 281574 93468 281580 93470
rect 281644 93468 281650 93532
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 110086 93196 110092 93260
rect 110156 93258 110162 93260
rect 110229 93258 110295 93261
rect 110156 93256 110295 93258
rect 110156 93200 110234 93256
rect 110290 93200 110295 93256
rect 110156 93198 110295 93200
rect 110156 93196 110162 93198
rect 110229 93195 110295 93198
rect 84326 92380 84332 92444
rect 84396 92442 84402 92444
rect 85113 92442 85179 92445
rect 88057 92444 88123 92445
rect 88006 92442 88012 92444
rect 84396 92440 85179 92442
rect 84396 92384 85118 92440
rect 85174 92384 85179 92440
rect 84396 92382 85179 92384
rect 87966 92382 88012 92442
rect 88076 92440 88123 92444
rect 88118 92384 88123 92440
rect 84396 92380 84402 92382
rect 85113 92379 85179 92382
rect 88006 92380 88012 92382
rect 88076 92380 88123 92384
rect 98126 92380 98132 92444
rect 98196 92442 98202 92444
rect 99281 92442 99347 92445
rect 100017 92444 100083 92445
rect 105721 92444 105787 92445
rect 106825 92444 106891 92445
rect 99966 92442 99972 92444
rect 98196 92440 99347 92442
rect 98196 92384 99286 92440
rect 99342 92384 99347 92440
rect 98196 92382 99347 92384
rect 99926 92382 99972 92442
rect 100036 92440 100083 92444
rect 105670 92442 105676 92444
rect 100078 92384 100083 92440
rect 98196 92380 98202 92382
rect 88057 92379 88123 92380
rect 99281 92379 99347 92382
rect 99966 92380 99972 92382
rect 100036 92380 100083 92384
rect 105630 92382 105676 92442
rect 105740 92440 105787 92444
rect 106774 92442 106780 92444
rect 105782 92384 105787 92440
rect 105670 92380 105676 92382
rect 105740 92380 105787 92384
rect 106734 92382 106780 92442
rect 106844 92440 106891 92444
rect 106886 92384 106891 92440
rect 106774 92380 106780 92382
rect 106844 92380 106891 92384
rect 113030 92380 113036 92444
rect 113100 92442 113106 92444
rect 114461 92442 114527 92445
rect 120257 92444 120323 92445
rect 123201 92444 123267 92445
rect 124121 92444 124187 92445
rect 125409 92444 125475 92445
rect 134425 92444 134491 92445
rect 151537 92444 151603 92445
rect 152089 92444 152155 92445
rect 120206 92442 120212 92444
rect 113100 92440 114527 92442
rect 113100 92384 114466 92440
rect 114522 92384 114527 92440
rect 113100 92382 114527 92384
rect 120166 92382 120212 92442
rect 120276 92440 120323 92444
rect 123150 92442 123156 92444
rect 120318 92384 120323 92440
rect 113100 92380 113106 92382
rect 100017 92379 100083 92380
rect 105721 92379 105787 92380
rect 106825 92379 106891 92380
rect 114461 92379 114527 92382
rect 120206 92380 120212 92382
rect 120276 92380 120323 92384
rect 123110 92382 123156 92442
rect 123220 92440 123267 92444
rect 124070 92442 124076 92444
rect 123262 92384 123267 92440
rect 123150 92380 123156 92382
rect 123220 92380 123267 92384
rect 124030 92382 124076 92442
rect 124140 92440 124187 92444
rect 125358 92442 125364 92444
rect 124182 92384 124187 92440
rect 124070 92380 124076 92382
rect 124140 92380 124187 92384
rect 125318 92382 125364 92442
rect 125428 92440 125475 92444
rect 134374 92442 134380 92444
rect 125470 92384 125475 92440
rect 125358 92380 125364 92382
rect 125428 92380 125475 92384
rect 134334 92382 134380 92442
rect 134444 92440 134491 92444
rect 151486 92442 151492 92444
rect 134486 92384 134491 92440
rect 134374 92380 134380 92382
rect 134444 92380 134491 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 152038 92442 152044 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 120257 92379 120323 92380
rect 123201 92379 123267 92380
rect 124121 92379 124187 92380
rect 125409 92379 125475 92380
rect 134425 92379 134491 92380
rect 151537 92379 151603 92380
rect 152089 92379 152155 92380
rect 109166 92244 109172 92308
rect 109236 92306 109242 92308
rect 109677 92306 109743 92309
rect 168230 92306 168236 92308
rect 109236 92304 109743 92306
rect 109236 92248 109682 92304
rect 109738 92248 109743 92304
rect 109236 92246 109743 92248
rect 109236 92244 109242 92246
rect 109677 92243 109743 92246
rect 122790 92246 168236 92306
rect 117998 92108 118004 92172
rect 118068 92170 118074 92172
rect 122790 92170 122850 92246
rect 168230 92244 168236 92246
rect 168300 92244 168306 92308
rect 118068 92110 122850 92170
rect 118068 92108 118074 92110
rect 101857 91764 101923 91765
rect 101806 91762 101812 91764
rect 101766 91702 101812 91762
rect 101876 91760 101923 91764
rect 101918 91704 101923 91760
rect 101806 91700 101812 91702
rect 101876 91700 101923 91704
rect 125726 91700 125732 91764
rect 125796 91762 125802 91764
rect 126881 91762 126947 91765
rect 125796 91760 126947 91762
rect 125796 91704 126886 91760
rect 126942 91704 126947 91760
rect 125796 91702 126947 91704
rect 125796 91700 125802 91702
rect 101857 91699 101923 91700
rect 126881 91699 126947 91702
rect 112294 91564 112300 91628
rect 112364 91626 112370 91628
rect 112713 91626 112779 91629
rect 112364 91624 112779 91626
rect 112364 91568 112718 91624
rect 112774 91568 112779 91624
rect 112364 91566 112779 91568
rect 112364 91564 112370 91566
rect 112713 91563 112779 91566
rect 119286 91564 119292 91628
rect 119356 91626 119362 91628
rect 119521 91626 119587 91629
rect 119356 91624 119587 91626
rect 119356 91568 119526 91624
rect 119582 91568 119587 91624
rect 119356 91566 119587 91568
rect 119356 91564 119362 91566
rect 119521 91563 119587 91566
rect 136030 91564 136036 91628
rect 136100 91626 136106 91628
rect 136265 91626 136331 91629
rect 136100 91624 136331 91626
rect 136100 91568 136270 91624
rect 136326 91568 136331 91624
rect 136100 91566 136331 91568
rect 136100 91564 136106 91566
rect 136265 91563 136331 91566
rect 122833 91492 122899 91493
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 122833 91427 122899 91428
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99097 91354 99163 91357
rect 98564 91352 99163 91354
rect 98564 91296 99102 91352
rect 99158 91296 99163 91352
rect 98564 91294 99163 91296
rect 98564 91292 98570 91294
rect 99097 91291 99163 91294
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 101949 91354 102015 91357
rect 100956 91352 102015 91354
rect 100956 91296 101954 91352
rect 102010 91296 102015 91352
rect 100956 91294 102015 91296
rect 100956 91292 100962 91294
rect 101949 91291 102015 91294
rect 113214 91292 113220 91356
rect 113284 91354 113290 91356
rect 114461 91354 114527 91357
rect 113284 91352 114527 91354
rect 113284 91296 114466 91352
rect 114522 91296 114527 91352
rect 113284 91294 114527 91296
rect 113284 91292 113290 91294
rect 114461 91291 114527 91294
rect 115422 91292 115428 91356
rect 115492 91354 115498 91356
rect 115841 91354 115907 91357
rect 115492 91352 115907 91354
rect 115492 91296 115846 91352
rect 115902 91296 115907 91352
rect 115492 91294 115907 91296
rect 115492 91292 115498 91294
rect 115841 91291 115907 91294
rect 126462 91292 126468 91356
rect 126532 91354 126538 91356
rect 126789 91354 126855 91357
rect 126532 91352 126855 91354
rect 126532 91296 126794 91352
rect 126850 91296 126855 91352
rect 126532 91294 126855 91296
rect 126532 91292 126538 91294
rect 126789 91291 126855 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75821 91218 75887 91221
rect 74828 91216 75887 91218
rect 74828 91160 75826 91216
rect 75882 91160 75887 91216
rect 74828 91158 75887 91160
rect 74828 91156 74834 91158
rect 75821 91155 75887 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89069 91218 89135 91221
rect 88996 91216 89135 91218
rect 88996 91160 89074 91216
rect 89130 91160 89135 91216
rect 88996 91158 89135 91160
rect 88996 91156 89002 91158
rect 89069 91155 89135 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90633 91218 90699 91221
rect 90284 91216 90699 91218
rect 90284 91160 90638 91216
rect 90694 91160 90699 91216
rect 90284 91158 90699 91160
rect 90284 91156 90290 91158
rect 90633 91155 90699 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 91921 91218 91987 91221
rect 91388 91216 91987 91218
rect 91388 91160 91926 91216
rect 91982 91160 91987 91216
rect 91388 91158 91987 91160
rect 91388 91156 91394 91158
rect 91921 91155 91987 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97073 91218 97139 91221
rect 96724 91216 97139 91218
rect 96724 91160 97078 91216
rect 97134 91160 97139 91216
rect 96724 91158 97139 91160
rect 96724 91156 96730 91158
rect 97073 91155 97139 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99189 91218 99255 91221
rect 100569 91220 100635 91221
rect 102041 91220 102107 91221
rect 100518 91218 100524 91220
rect 99116 91216 99255 91218
rect 99116 91160 99194 91216
rect 99250 91160 99255 91216
rect 99116 91158 99255 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 101990 91218 101996 91220
rect 100630 91160 100635 91216
rect 99116 91156 99122 91158
rect 99189 91155 99255 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 102102 91160 102107 91216
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103329 91218 103395 91221
rect 102796 91216 103395 91218
rect 102796 91160 103334 91216
rect 103390 91160 103395 91216
rect 102796 91158 103395 91160
rect 102796 91156 102802 91158
rect 100569 91155 100635 91156
rect 102041 91155 102107 91156
rect 103329 91155 103395 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 104636 91156 104642 91158
rect 104801 91155 104867 91158
rect 105486 91156 105492 91220
rect 105556 91218 105562 91220
rect 105721 91218 105787 91221
rect 105556 91216 105787 91218
rect 105556 91160 105726 91216
rect 105782 91160 105787 91216
rect 105556 91158 105787 91160
rect 105556 91156 105562 91158
rect 105721 91155 105787 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107101 91218 107167 91221
rect 106476 91216 107167 91218
rect 106476 91160 107106 91216
rect 107162 91160 107167 91216
rect 106476 91158 107167 91160
rect 106476 91156 106482 91158
rect 107101 91155 107167 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108757 91218 108823 91221
rect 108132 91216 108823 91218
rect 108132 91160 108762 91216
rect 108818 91160 108823 91216
rect 108132 91158 108823 91160
rect 108132 91156 108138 91158
rect 108757 91155 108823 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111057 91218 111123 91221
rect 110708 91216 111123 91218
rect 110708 91160 111062 91216
rect 111118 91160 111123 91216
rect 110708 91158 111123 91160
rect 110708 91156 110714 91158
rect 111057 91155 111123 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111701 91218 111767 91221
rect 111260 91216 111767 91218
rect 111260 91160 111706 91216
rect 111762 91160 111767 91216
rect 111260 91158 111767 91160
rect 111260 91156 111266 91158
rect 111701 91155 111767 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 114369 91220 114435 91221
rect 114318 91218 114324 91220
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 114278 91158 114324 91218
rect 114388 91216 114435 91220
rect 114430 91160 114435 91216
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 114318 91156 114324 91158
rect 114388 91156 114435 91160
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115749 91218 115815 91221
rect 114940 91216 115815 91218
rect 114940 91160 115754 91216
rect 115810 91160 115815 91216
rect 114940 91158 115815 91160
rect 114940 91156 114946 91158
rect 114369 91155 114435 91156
rect 115749 91155 115815 91158
rect 117078 91156 117084 91220
rect 117148 91218 117154 91220
rect 117221 91218 117287 91221
rect 118233 91220 118299 91221
rect 119705 91220 119771 91221
rect 118182 91218 118188 91220
rect 117148 91216 117287 91218
rect 117148 91160 117226 91216
rect 117282 91160 117287 91216
rect 117148 91158 117287 91160
rect 118142 91158 118188 91218
rect 118252 91216 118299 91220
rect 119654 91218 119660 91220
rect 118294 91160 118299 91216
rect 117148 91156 117154 91158
rect 117221 91155 117287 91158
rect 118182 91156 118188 91158
rect 118252 91156 118299 91160
rect 119614 91158 119660 91218
rect 119724 91216 119771 91220
rect 119766 91160 119771 91216
rect 119654 91156 119660 91158
rect 119724 91156 119771 91160
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 122281 91218 122347 91221
rect 121748 91216 122347 91218
rect 121748 91160 122286 91216
rect 122342 91160 122347 91216
rect 121748 91158 122347 91160
rect 121748 91156 121754 91158
rect 118233 91155 118299 91156
rect 119705 91155 119771 91156
rect 122281 91155 122347 91158
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 125501 91218 125567 91221
rect 126697 91220 126763 91221
rect 126646 91218 126652 91220
rect 124508 91216 125567 91218
rect 124508 91160 125506 91216
rect 125562 91160 125567 91216
rect 124508 91158 125567 91160
rect 126606 91158 126652 91218
rect 126716 91216 126763 91220
rect 126758 91160 126763 91216
rect 124508 91156 124514 91158
rect 125501 91155 125567 91158
rect 126646 91156 126652 91158
rect 126716 91156 126763 91160
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 129457 91220 129523 91221
rect 130745 91220 130811 91221
rect 132401 91220 132467 91221
rect 151721 91220 151787 91221
rect 129406 91218 129412 91220
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 129366 91158 129412 91218
rect 129476 91216 129523 91220
rect 130694 91218 130700 91220
rect 129518 91160 129523 91216
rect 127636 91156 127642 91158
rect 126697 91155 126763 91156
rect 128261 91155 128327 91158
rect 129406 91156 129412 91158
rect 129476 91156 129523 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 132350 91218 132356 91220
rect 130806 91160 130811 91216
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 151670 91218 151676 91220
rect 132462 91160 132467 91216
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 151630 91158 151676 91218
rect 151740 91216 151787 91220
rect 151782 91160 151787 91216
rect 151670 91156 151676 91158
rect 151740 91156 151787 91160
rect 129457 91155 129523 91156
rect 130745 91155 130811 91156
rect 132401 91155 132467 91156
rect 151721 91155 151787 91156
rect 66069 91082 66135 91085
rect 172094 91082 172100 91084
rect 66069 91080 172100 91082
rect 66069 91024 66074 91080
rect 66130 91024 172100 91080
rect 66069 91022 172100 91024
rect 66069 91019 66135 91022
rect 172094 91020 172100 91022
rect 172164 91020 172170 91084
rect 62021 89722 62087 89725
rect 211889 89722 211955 89725
rect 62021 89720 211955 89722
rect 62021 89664 62026 89720
rect 62082 89664 211894 89720
rect 211950 89664 211955 89720
rect 62021 89662 211955 89664
rect 62021 89659 62087 89662
rect 211889 89659 211955 89662
rect 97073 88226 97139 88229
rect 169150 88226 169156 88228
rect 97073 88224 169156 88226
rect 97073 88168 97078 88224
rect 97134 88168 169156 88224
rect 97073 88166 169156 88168
rect 97073 88163 97139 88166
rect 169150 88164 169156 88166
rect 169220 88164 169226 88228
rect 57830 86804 57836 86868
rect 57900 86866 57906 86868
rect 280153 86866 280219 86869
rect 57900 86864 280219 86866
rect 57900 86808 280158 86864
rect 280214 86808 280219 86864
rect 57900 86806 280219 86808
rect 57900 86804 57906 86806
rect 280153 86803 280219 86806
rect 108757 86730 108823 86733
rect 170438 86730 170444 86732
rect 108757 86728 170444 86730
rect 108757 86672 108762 86728
rect 108818 86672 170444 86728
rect 108757 86670 170444 86672
rect 108757 86667 108823 86670
rect 170438 86668 170444 86670
rect 170508 86668 170514 86732
rect 132401 86594 132467 86597
rect 166206 86594 166212 86596
rect 132401 86592 166212 86594
rect 132401 86536 132406 86592
rect 132462 86536 166212 86592
rect 132401 86534 166212 86536
rect 132401 86531 132467 86534
rect 166206 86532 166212 86534
rect 166276 86532 166282 86596
rect 582741 86186 582807 86189
rect 583520 86186 584960 86276
rect 582741 86184 584960 86186
rect 582741 86128 582746 86184
rect 582802 86128 584960 86184
rect 582741 86126 584960 86128
rect 582741 86123 582807 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 101949 84146 102015 84149
rect 173198 84146 173204 84148
rect 101949 84144 173204 84146
rect 101949 84088 101954 84144
rect 102010 84088 173204 84144
rect 101949 84086 173204 84088
rect 101949 84083 102015 84086
rect 173198 84084 173204 84086
rect 173268 84084 173274 84148
rect 114369 84010 114435 84013
rect 166390 84010 166396 84012
rect 114369 84008 166396 84010
rect 114369 83952 114374 84008
rect 114430 83952 166396 84008
rect 114369 83950 166396 83952
rect 114369 83947 114435 83950
rect 166390 83948 166396 83950
rect 166460 83948 166466 84012
rect 102041 78570 102107 78573
rect 168966 78570 168972 78572
rect 102041 78568 168972 78570
rect 102041 78512 102046 78568
rect 102102 78512 168972 78568
rect 102041 78510 168972 78512
rect 102041 78507 102107 78510
rect 168966 78508 168972 78510
rect 169036 78508 169042 78572
rect 115841 77210 115907 77213
rect 170254 77210 170260 77212
rect 115841 77208 170260 77210
rect 115841 77152 115846 77208
rect 115902 77152 170260 77208
rect 115841 77150 170260 77152
rect 115841 77147 115907 77150
rect 170254 77148 170260 77150
rect 170324 77148 170330 77212
rect 56593 73810 56659 73813
rect 258758 73810 258764 73812
rect 56593 73808 258764 73810
rect 56593 73752 56598 73808
rect 56654 73752 258764 73808
rect 56593 73750 258764 73752
rect 56593 73747 56659 73750
rect 258758 73748 258764 73750
rect 258828 73748 258834 73812
rect 582465 72994 582531 72997
rect 583520 72994 584960 73084
rect 582465 72992 584960 72994
rect 582465 72936 582470 72992
rect 582526 72936 584960 72992
rect 582465 72934 584960 72936
rect 582465 72931 582531 72934
rect 583520 72844 584960 72934
rect 63493 72450 63559 72453
rect 264094 72450 264100 72452
rect 63493 72448 264100 72450
rect 63493 72392 63498 72448
rect 63554 72392 264100 72448
rect 63493 72390 264100 72392
rect 63493 72387 63559 72390
rect 264094 72388 264100 72390
rect 264164 72388 264170 72452
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 62982 69532 62988 69596
rect 63052 69594 63058 69596
rect 332685 69594 332751 69597
rect 63052 69592 332751 69594
rect 63052 69536 332690 69592
rect 332746 69536 332751 69592
rect 63052 69534 332751 69536
rect 63052 69532 63058 69534
rect 332685 69531 332751 69534
rect 92473 64154 92539 64157
rect 239254 64154 239260 64156
rect 92473 64152 239260 64154
rect 92473 64096 92478 64152
rect 92534 64096 239260 64152
rect 92473 64094 239260 64096
rect 92473 64091 92539 64094
rect 239254 64092 239260 64094
rect 239324 64092 239330 64156
rect 13813 62794 13879 62797
rect 255814 62794 255820 62796
rect 13813 62792 255820 62794
rect 13813 62736 13818 62792
rect 13874 62736 255820 62792
rect 13813 62734 255820 62736
rect 13813 62731 13879 62734
rect 255814 62732 255820 62734
rect 255884 62732 255890 62796
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 27613 51778 27679 51781
rect 254526 51778 254532 51780
rect 27613 51776 254532 51778
rect 27613 51720 27618 51776
rect 27674 51720 254532 51776
rect 27613 51718 254532 51720
rect 27613 51715 27679 51718
rect 254526 51716 254532 51718
rect 254596 51716 254602 51780
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 98637 43482 98703 43485
rect 265750 43482 265756 43484
rect 98637 43480 265756 43482
rect 98637 43424 98642 43480
rect 98698 43424 265756 43480
rect 98637 43422 265756 43424
rect 98637 43419 98703 43422
rect 265750 43420 265756 43422
rect 265820 43420 265826 43484
rect 38653 40626 38719 40629
rect 257286 40626 257292 40628
rect 38653 40624 257292 40626
rect 38653 40568 38658 40624
rect 38714 40568 257292 40624
rect 38653 40566 257292 40568
rect 38653 40563 38719 40566
rect 257286 40564 257292 40566
rect 257356 40564 257362 40628
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 42793 30970 42859 30973
rect 258574 30970 258580 30972
rect 42793 30968 258580 30970
rect 42793 30912 42798 30968
rect 42854 30912 258580 30968
rect 42793 30910 258580 30912
rect 42793 30907 42859 30910
rect 258574 30908 258580 30910
rect 258644 30908 258650 30972
rect 2865 25530 2931 25533
rect 262806 25530 262812 25532
rect 2865 25528 262812 25530
rect 2865 25472 2870 25528
rect 2926 25472 262812 25528
rect 2865 25470 262812 25472
rect 2865 25467 2931 25470
rect 262806 25468 262812 25470
rect 262876 25468 262882 25532
rect 53925 24850 53991 24853
rect 55121 24850 55187 24853
rect 227662 24850 227668 24852
rect 53925 24848 227668 24850
rect 53925 24792 53930 24848
rect 53986 24792 55126 24848
rect 55182 24792 227668 24848
rect 53925 24790 227668 24792
rect 53925 24787 53991 24790
rect 55121 24787 55187 24790
rect 227662 24788 227668 24790
rect 227732 24788 227738 24852
rect 1393 24170 1459 24173
rect 53925 24170 53991 24173
rect 1393 24168 53991 24170
rect 1393 24112 1398 24168
rect 1454 24112 53930 24168
rect 53986 24112 53991 24168
rect 1393 24110 53991 24112
rect 1393 24107 1459 24110
rect 53925 24107 53991 24110
rect 70393 24170 70459 24173
rect 262070 24170 262076 24172
rect 70393 24168 262076 24170
rect 70393 24112 70398 24168
rect 70454 24112 262076 24168
rect 70393 24110 262076 24112
rect 70393 24107 70459 24110
rect 262070 24108 262076 24110
rect 262140 24108 262146 24172
rect 19425 19954 19491 19957
rect 228214 19954 228220 19956
rect 19425 19952 228220 19954
rect 19425 19896 19430 19952
rect 19486 19896 228220 19952
rect 19425 19894 228220 19896
rect 19425 19891 19491 19894
rect 228214 19892 228220 19894
rect 228284 19892 228290 19956
rect 582373 19818 582439 19821
rect 583520 19818 584960 19908
rect 582373 19816 584960 19818
rect 582373 19760 582378 19816
rect 582434 19760 584960 19816
rect 582373 19758 584960 19760
rect 582373 19755 582439 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 117313 11658 117379 11661
rect 232446 11658 232452 11660
rect 117313 11656 232452 11658
rect 117313 11600 117318 11656
rect 117374 11600 232452 11656
rect 117313 11598 232452 11600
rect 117313 11595 117379 11598
rect 232446 11596 232452 11598
rect 232516 11596 232522 11660
rect 582557 6626 582623 6629
rect 583520 6626 584960 6716
rect 582557 6624 584960 6626
rect -960 6490 480 6580
rect 582557 6568 582562 6624
rect 582618 6568 584960 6624
rect 582557 6566 584960 6568
rect 582557 6563 582623 6566
rect 2957 6490 3023 6493
rect -960 6488 3023 6490
rect -960 6432 2962 6488
rect 3018 6432 3023 6488
rect 583520 6476 584960 6566
rect -960 6430 3023 6432
rect -960 6340 480 6430
rect 2957 6427 3023 6430
rect 242014 4796 242020 4860
rect 242084 4858 242090 4860
rect 257061 4858 257127 4861
rect 242084 4856 257127 4858
rect 242084 4800 257066 4856
rect 257122 4800 257127 4856
rect 242084 4798 257127 4800
rect 242084 4796 242090 4798
rect 257061 4795 257127 4798
rect 295926 3844 295932 3908
rect 295996 3906 296002 3908
rect 298461 3906 298527 3909
rect 295996 3904 298527 3906
rect 295996 3848 298466 3904
rect 298522 3848 298527 3904
rect 295996 3846 298527 3848
rect 295996 3844 296002 3846
rect 298461 3843 298527 3846
rect 302734 3844 302740 3908
rect 302804 3906 302810 3908
rect 307937 3906 308003 3909
rect 302804 3904 308003 3906
rect 302804 3848 307942 3904
rect 307998 3848 308003 3904
rect 302804 3846 308003 3848
rect 302804 3844 302810 3846
rect 307937 3843 308003 3846
rect 298686 3572 298692 3636
rect 298756 3634 298762 3636
rect 303153 3634 303219 3637
rect 298756 3632 303219 3634
rect 298756 3576 303158 3632
rect 303214 3576 303219 3632
rect 298756 3574 303219 3576
rect 298756 3572 298762 3574
rect 303153 3571 303219 3574
rect 240358 3436 240364 3500
rect 240428 3498 240434 3500
rect 240501 3498 240567 3501
rect 240428 3496 240567 3498
rect 240428 3440 240506 3496
rect 240562 3440 240567 3496
rect 240428 3438 240567 3440
rect 240428 3436 240434 3438
rect 240501 3435 240567 3438
rect 244222 3436 244228 3500
rect 244292 3498 244298 3500
rect 245193 3498 245259 3501
rect 244292 3496 245259 3498
rect 244292 3440 245198 3496
rect 245254 3440 245259 3496
rect 244292 3438 245259 3440
rect 244292 3436 244298 3438
rect 245193 3435 245259 3438
rect 245694 3436 245700 3500
rect 245764 3498 245770 3500
rect 246389 3498 246455 3501
rect 245764 3496 246455 3498
rect 245764 3440 246394 3496
rect 246450 3440 246455 3496
rect 245764 3438 246455 3440
rect 245764 3436 245770 3438
rect 246389 3435 246455 3438
rect 248454 3436 248460 3500
rect 248524 3498 248530 3500
rect 248781 3498 248847 3501
rect 248524 3496 248847 3498
rect 248524 3440 248786 3496
rect 248842 3440 248847 3496
rect 248524 3438 248847 3440
rect 248524 3436 248530 3438
rect 248781 3435 248847 3438
rect 249742 3436 249748 3500
rect 249812 3498 249818 3500
rect 249977 3498 250043 3501
rect 249812 3496 250043 3498
rect 249812 3440 249982 3496
rect 250038 3440 250043 3496
rect 249812 3438 250043 3440
rect 249812 3436 249818 3438
rect 249977 3435 250043 3438
rect 251214 3436 251220 3500
rect 251284 3498 251290 3500
rect 252369 3498 252435 3501
rect 251284 3496 252435 3498
rect 251284 3440 252374 3496
rect 252430 3440 252435 3496
rect 251284 3438 252435 3440
rect 251284 3436 251290 3438
rect 252369 3435 252435 3438
rect 252502 3436 252508 3500
rect 252572 3498 252578 3500
rect 253473 3498 253539 3501
rect 252572 3496 253539 3498
rect 252572 3440 253478 3496
rect 253534 3440 253539 3496
rect 252572 3438 253539 3440
rect 252572 3436 252578 3438
rect 253473 3435 253539 3438
rect 255262 3436 255268 3500
rect 255332 3498 255338 3500
rect 255865 3498 255931 3501
rect 259453 3500 259519 3501
rect 259453 3498 259500 3500
rect 255332 3496 255931 3498
rect 255332 3440 255870 3496
rect 255926 3440 255931 3496
rect 255332 3438 255931 3440
rect 259408 3496 259500 3498
rect 259408 3440 259458 3496
rect 259408 3438 259500 3440
rect 255332 3436 255338 3438
rect 255865 3435 255931 3438
rect 259453 3436 259500 3438
rect 259564 3436 259570 3500
rect 288382 3436 288388 3500
rect 288452 3498 288458 3500
rect 288985 3498 289051 3501
rect 288452 3496 289051 3498
rect 288452 3440 288990 3496
rect 289046 3440 289051 3496
rect 288452 3438 289051 3440
rect 288452 3436 288458 3438
rect 259453 3435 259519 3436
rect 288985 3435 289051 3438
rect 291142 3436 291148 3500
rect 291212 3498 291218 3500
rect 291377 3498 291443 3501
rect 291212 3496 291443 3498
rect 291212 3440 291382 3496
rect 291438 3440 291443 3496
rect 291212 3438 291443 3440
rect 291212 3436 291218 3438
rect 291377 3435 291443 3438
rect 292614 3436 292620 3500
rect 292684 3498 292690 3500
rect 293677 3498 293743 3501
rect 292684 3496 293743 3498
rect 292684 3440 293682 3496
rect 293738 3440 293743 3496
rect 292684 3438 293743 3440
rect 292684 3436 292690 3438
rect 293677 3435 293743 3438
rect 295374 3436 295380 3500
rect 295444 3498 295450 3500
rect 296069 3498 296135 3501
rect 295444 3496 296135 3498
rect 295444 3440 296074 3496
rect 296130 3440 296135 3496
rect 295444 3438 296135 3440
rect 295444 3436 295450 3438
rect 296069 3435 296135 3438
rect 299606 3436 299612 3500
rect 299676 3498 299682 3500
rect 300761 3498 300827 3501
rect 299676 3496 300827 3498
rect 299676 3440 300766 3496
rect 300822 3440 300827 3496
rect 299676 3438 300827 3440
rect 299676 3436 299682 3438
rect 300761 3435 300827 3438
rect 304942 3436 304948 3500
rect 305012 3498 305018 3500
rect 305545 3498 305611 3501
rect 305012 3496 305611 3498
rect 305012 3440 305550 3496
rect 305606 3440 305611 3496
rect 305012 3438 305611 3440
rect 305012 3436 305018 3438
rect 305545 3435 305611 3438
rect 249006 3300 249012 3364
rect 249076 3362 249082 3364
rect 258257 3362 258323 3365
rect 249076 3360 258323 3362
rect 249076 3304 258262 3360
rect 258318 3304 258323 3360
rect 249076 3302 258323 3304
rect 249076 3300 249082 3302
rect 258257 3299 258323 3302
rect 268326 3300 268332 3364
rect 268396 3362 268402 3364
rect 279509 3362 279575 3365
rect 268396 3360 279575 3362
rect 268396 3304 279514 3360
rect 279570 3304 279575 3360
rect 268396 3302 279575 3304
rect 268396 3300 268402 3302
rect 279509 3299 279575 3302
<< via3 >>
rect 111012 702476 111076 702540
rect 57836 586332 57900 586396
rect 115980 584020 116044 584084
rect 114508 581708 114572 581772
rect 118740 578852 118804 578916
rect 111748 578232 111812 578236
rect 111748 578176 111762 578232
rect 111762 578176 111812 578232
rect 111748 578172 111812 578176
rect 66116 577084 66180 577148
rect 66668 571780 66732 571844
rect 68876 570284 68940 570348
rect 64644 565796 64708 565860
rect 106412 564436 106476 564500
rect 61884 561852 61948 561916
rect 105492 561852 105556 561916
rect 60596 560492 60660 560556
rect 107700 557636 107764 557700
rect 62988 547980 63052 548044
rect 107884 546756 107948 546820
rect 111012 540092 111076 540156
rect 70348 538732 70412 538796
rect 103652 538052 103716 538116
rect 57836 537508 57900 537572
rect 57836 537372 57900 537436
rect 98500 537372 98564 537436
rect 114508 536012 114572 536076
rect 53604 532204 53668 532268
rect 48084 532068 48148 532132
rect 44036 531932 44100 531996
rect 118740 495484 118804 495548
rect 118740 494940 118804 495004
rect 50844 494804 50908 494868
rect 124444 494668 124508 494732
rect 52316 492628 52380 492692
rect 53052 491948 53116 492012
rect 109540 491404 109604 491468
rect 111012 491268 111076 491332
rect 99420 490588 99484 490652
rect 59124 490452 59188 490516
rect 115980 490044 116044 490108
rect 98500 489908 98564 489972
rect 101996 489908 102060 489972
rect 122788 489908 122852 489972
rect 55076 489092 55140 489156
rect 115796 488412 115860 488476
rect 69060 486508 69124 486572
rect 118924 486372 118988 486436
rect 111748 485012 111812 485076
rect 115612 485012 115676 485076
rect 70348 484604 70412 484668
rect 68692 482564 68756 482628
rect 65932 480524 65996 480588
rect 112300 478892 112364 478956
rect 66116 478484 66180 478548
rect 106412 478076 106476 478140
rect 61700 477396 61764 477460
rect 117084 477396 117148 477460
rect 118740 475900 118804 475964
rect 66668 473996 66732 474060
rect 118004 473996 118068 474060
rect 66668 473724 66732 473788
rect 68876 471004 68940 471068
rect 104940 471140 105004 471204
rect 105492 467876 105556 467940
rect 64644 467740 64708 467804
rect 64644 467196 64708 467260
rect 99972 466244 100036 466308
rect 107700 465700 107764 465764
rect 61884 463524 61948 463588
rect 116532 463524 116596 463588
rect 102732 461484 102796 461548
rect 60596 460940 60660 461004
rect 115796 459580 115860 459644
rect 115612 458220 115676 458284
rect 107884 456044 107948 456108
rect 62988 447748 63052 447812
rect 103836 445708 103900 445772
rect 133092 445708 133156 445772
rect 103836 444348 103900 444412
rect 61884 442852 61948 442916
rect 61884 441628 61948 441692
rect 53604 441084 53668 441148
rect 99052 441084 99116 441148
rect 59124 440948 59188 441012
rect 65932 440328 65996 440332
rect 65932 440272 65982 440328
rect 65982 440272 65996 440328
rect 65932 440268 65996 440272
rect 102732 440132 102796 440196
rect 64644 439452 64708 439516
rect 69060 439452 69124 439516
rect 124260 439316 124324 439380
rect 99420 439044 99484 439108
rect 68692 438908 68756 438972
rect 55076 438772 55140 438836
rect 124444 438772 124508 438836
rect 125732 438772 125796 438836
rect 99972 438636 100036 438700
rect 70348 437684 70412 437748
rect 57836 437412 57900 437476
rect 105492 435916 105556 435980
rect 44036 434556 44100 434620
rect 48084 433196 48148 433260
rect 48084 430612 48148 430676
rect 128676 404908 128740 404972
rect 61700 401644 61764 401708
rect 109540 401236 109604 401300
rect 66116 400284 66180 400348
rect 53604 399604 53668 399668
rect 50844 399468 50908 399532
rect 129780 399468 129844 399532
rect 168420 398788 168484 398852
rect 52316 397972 52380 398036
rect 115980 394028 116044 394092
rect 173020 393892 173084 393956
rect 101996 393348 102060 393412
rect 133828 393348 133892 393412
rect 57836 391172 57900 391236
rect 121684 390628 121748 390692
rect 122604 389812 122668 389876
rect 59124 389132 59188 389196
rect 111012 389132 111076 389196
rect 122420 388860 122484 388924
rect 99052 388316 99116 388380
rect 123340 388316 123404 388380
rect 115428 387772 115492 387836
rect 120764 387772 120828 387836
rect 122604 387772 122668 387836
rect 70532 387636 70596 387700
rect 53052 387500 53116 387564
rect 251220 385596 251284 385660
rect 112300 385324 112364 385388
rect 66116 384780 66180 384844
rect 115428 384508 115492 384572
rect 69980 383148 70044 383212
rect 118924 381516 118988 381580
rect 118924 380972 118988 381036
rect 69060 380292 69124 380356
rect 52316 377708 52380 377772
rect 70532 377708 70596 377772
rect 62988 377300 63052 377364
rect 252508 377300 252572 377364
rect 68876 377164 68940 377228
rect 65380 375940 65444 376004
rect 255268 375940 255332 376004
rect 68876 372872 68940 372876
rect 68876 372816 68926 372872
rect 68926 372816 68940 372872
rect 68876 372812 68940 372816
rect 117084 372676 117148 372740
rect 118004 371316 118068 371380
rect 55076 370500 55140 370564
rect 122236 370500 122300 370564
rect 304948 370500 305012 370564
rect 299612 369004 299676 369068
rect 118740 368596 118804 368660
rect 259500 367644 259564 367708
rect 120764 366284 120828 366348
rect 302740 363564 302804 363628
rect 242020 362204 242084 362268
rect 123340 360844 123404 360908
rect 115980 357308 116044 357372
rect 124812 356084 124876 356148
rect 61700 355268 61764 355332
rect 70348 342892 70412 342956
rect 61884 342212 61948 342276
rect 124812 341396 124876 341460
rect 70532 340988 70596 341052
rect 48084 340776 48148 340780
rect 48084 340720 48098 340776
rect 48098 340720 48148 340776
rect 48084 340716 48148 340720
rect 64644 340716 64708 340780
rect 52316 339628 52380 339692
rect 44036 339356 44100 339420
rect 128676 337996 128740 338060
rect 57836 337860 57900 337924
rect 61332 337920 61396 337924
rect 61332 337864 61382 337920
rect 61382 337864 61396 337920
rect 61332 337860 61396 337864
rect 126100 337452 126164 337516
rect 124812 337316 124876 337380
rect 70532 336092 70596 336156
rect 292620 336092 292684 336156
rect 70348 335956 70412 336020
rect 248460 334732 248524 334796
rect 291148 334596 291212 334660
rect 53604 333916 53668 333980
rect 288388 333236 288452 333300
rect 125732 332480 125796 332484
rect 125732 332424 125782 332480
rect 125782 332424 125796 332480
rect 125732 332420 125796 332424
rect 244228 331740 244292 331804
rect 122604 331060 122668 331124
rect 55076 330380 55140 330444
rect 133092 329760 133156 329764
rect 133092 329704 133142 329760
rect 133142 329704 133156 329760
rect 133092 329700 133156 329704
rect 298692 329020 298756 329084
rect 129780 328400 129844 328404
rect 129780 328344 129830 328400
rect 129830 328344 129844 328400
rect 129780 328340 129844 328344
rect 124260 324320 124324 324324
rect 124260 324264 124310 324320
rect 124310 324264 124324 324320
rect 124260 324260 124324 324264
rect 61700 323716 61764 323780
rect 65380 323580 65444 323644
rect 245700 322084 245764 322148
rect 249748 320724 249812 320788
rect 68876 316644 68940 316708
rect 295932 316644 295996 316708
rect 240364 315284 240428 315348
rect 121684 314256 121748 314260
rect 121684 314200 121698 314256
rect 121698 314200 121748 314256
rect 121684 314196 121748 314200
rect 268332 306988 268396 307052
rect 69060 305628 69124 305692
rect 70900 304132 70964 304196
rect 249012 302772 249076 302836
rect 247724 298284 247788 298348
rect 227668 298148 227732 298212
rect 118740 295972 118804 296036
rect 123340 294204 123404 294268
rect 287100 293932 287164 293996
rect 250300 292708 250364 292772
rect 242940 289852 243004 289916
rect 70532 286724 70596 286788
rect 124812 283460 124876 283524
rect 241652 280196 241716 280260
rect 66116 276252 66180 276316
rect 119292 275572 119356 275636
rect 50844 265100 50908 265164
rect 123340 255852 123404 255916
rect 61516 253812 61580 253876
rect 126100 253132 126164 253196
rect 57836 251364 57900 251428
rect 65932 250412 65996 250476
rect 70532 248372 70596 248436
rect 120028 246468 120092 246532
rect 240548 245652 240612 245716
rect 59124 240348 59188 240412
rect 61332 238444 61396 238508
rect 119292 238444 119356 238508
rect 61516 235180 61580 235244
rect 288572 228244 288636 228308
rect 230428 227020 230492 227084
rect 285628 226884 285692 226948
rect 133828 226264 133892 226268
rect 133828 226208 133878 226264
rect 133878 226208 133892 226264
rect 133828 226204 133892 226208
rect 50844 225524 50908 225588
rect 291332 222804 291396 222868
rect 278820 213148 278884 213212
rect 285812 208932 285876 208996
rect 233188 197916 233252 197980
rect 236500 196692 236564 196756
rect 65932 196556 65996 196620
rect 280292 192476 280356 192540
rect 237604 190980 237668 191044
rect 287284 189620 287348 189684
rect 290596 187036 290660 187100
rect 237420 186900 237484 186964
rect 66116 184180 66180 184244
rect 245884 182820 245948 182884
rect 70900 180100 70964 180164
rect 166212 179420 166276 179484
rect 294276 178740 294340 178804
rect 295380 178604 295444 178668
rect 97028 177652 97092 177716
rect 98316 177652 98380 177716
rect 100708 177652 100772 177716
rect 104572 177652 104636 177716
rect 113220 177652 113284 177716
rect 114324 177652 114388 177716
rect 118372 177712 118436 177716
rect 118372 177656 118422 177712
rect 118422 177656 118436 177712
rect 118372 177652 118436 177656
rect 119476 177652 119540 177716
rect 121868 177652 121932 177716
rect 127020 177652 127084 177716
rect 129412 177712 129476 177716
rect 129412 177656 129462 177712
rect 129462 177656 129476 177712
rect 129412 177652 129476 177656
rect 234660 177516 234724 177580
rect 228956 177380 229020 177444
rect 238524 177244 238588 177308
rect 279372 177108 279436 177172
rect 109540 176972 109604 177036
rect 125732 176972 125796 177036
rect 133092 177032 133156 177036
rect 133092 176976 133142 177032
rect 133142 176976 133156 177032
rect 133092 176972 133156 176976
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 105676 176760 105740 176764
rect 105676 176704 105726 176760
rect 105726 176704 105740 176760
rect 105676 176700 105740 176704
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 123156 176700 123220 176764
rect 130700 176760 130764 176764
rect 130700 176704 130750 176760
rect 130750 176704 130764 176760
rect 130700 176700 130764 176704
rect 132356 176760 132420 176764
rect 132356 176704 132406 176760
rect 132406 176704 132420 176760
rect 132356 176700 132420 176704
rect 134380 176700 134444 176764
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 281580 176156 281644 176220
rect 229508 175884 229572 175948
rect 268516 175748 268580 175812
rect 116900 175536 116964 175540
rect 116900 175480 116950 175536
rect 116950 175480 116964 175536
rect 116900 175476 116964 175480
rect 120764 175536 120828 175540
rect 120764 175480 120814 175536
rect 120814 175480 120828 175536
rect 120764 175476 120828 175480
rect 124444 175536 124508 175540
rect 124444 175480 124494 175536
rect 124494 175480 124508 175536
rect 124444 175476 124508 175480
rect 158852 175536 158916 175540
rect 158852 175480 158902 175536
rect 158902 175480 158916 175536
rect 158852 175476 158916 175480
rect 110644 175400 110708 175404
rect 110644 175344 110694 175400
rect 110694 175344 110708 175400
rect 110644 175340 110708 175344
rect 112116 175340 112180 175404
rect 166396 175340 166460 175404
rect 229140 174932 229204 174996
rect 279372 175204 279436 175268
rect 268516 174932 268580 174996
rect 229140 174252 229204 174316
rect 281580 171668 281644 171732
rect 168420 168404 168484 168468
rect 238708 168328 238772 168332
rect 238708 168272 238758 168328
rect 238758 168272 238772 168328
rect 238708 168268 238772 168272
rect 237604 167588 237668 167652
rect 239076 167044 239140 167108
rect 268516 167180 268580 167244
rect 268516 166772 268580 166836
rect 166396 162828 166460 162892
rect 268516 162964 268580 163028
rect 166212 161604 166276 161668
rect 268516 159836 268580 159900
rect 237972 159020 238036 159084
rect 237420 158748 237484 158812
rect 229508 158068 229572 158132
rect 279372 156708 279436 156772
rect 247724 154804 247788 154868
rect 240548 153172 240612 153236
rect 240732 152356 240796 152420
rect 233188 148684 233252 148748
rect 230428 147732 230492 147796
rect 268516 147868 268580 147932
rect 230980 146100 231044 146164
rect 268516 146100 268580 146164
rect 166212 144876 166276 144940
rect 233740 143924 233804 143988
rect 242940 142972 243004 143036
rect 233924 142700 233988 142764
rect 245884 141612 245948 141676
rect 231348 141340 231412 141404
rect 241652 141068 241716 141132
rect 268516 140932 268580 140996
rect 268516 140524 268580 140588
rect 262812 140116 262876 140180
rect 232452 138348 232516 138412
rect 236500 138212 236564 138276
rect 234660 137804 234724 137868
rect 170260 136716 170324 136780
rect 280292 136988 280356 137052
rect 166396 135492 166460 135556
rect 239076 135764 239140 135828
rect 239260 135764 239324 135828
rect 268516 134132 268580 134196
rect 231348 133784 231412 133788
rect 231348 133728 231362 133784
rect 231362 133728 231412 133784
rect 231348 133724 231412 133728
rect 268516 133724 268580 133788
rect 170444 132772 170508 132836
rect 262076 133180 262140 133244
rect 231164 132908 231228 132972
rect 264100 132500 264164 132564
rect 258764 131548 258828 131612
rect 258580 130188 258644 130252
rect 168972 129780 169036 129844
rect 257292 128964 257356 129028
rect 173204 128420 173268 128484
rect 287284 128692 287348 128756
rect 268516 128556 268580 128620
rect 268516 128148 268580 128212
rect 169156 127196 169220 127260
rect 255820 127060 255884 127124
rect 268516 127196 268580 127260
rect 288572 127060 288636 127124
rect 268516 126788 268580 126852
rect 231716 126244 231780 126308
rect 230980 125972 231044 126036
rect 231716 125428 231780 125492
rect 230428 125292 230492 125356
rect 231164 123524 231228 123588
rect 268516 122980 268580 123044
rect 268516 122572 268580 122636
rect 268516 121620 268580 121684
rect 268516 121212 268580 121276
rect 173020 119308 173084 119372
rect 237972 118356 238036 118420
rect 168236 117948 168300 118012
rect 268516 117268 268580 117332
rect 268516 116452 268580 116516
rect 240732 115500 240796 115564
rect 254532 114548 254596 114612
rect 294276 110468 294340 110532
rect 290596 109108 290660 109172
rect 268516 107884 268580 107948
rect 268516 107476 268580 107540
rect 287100 106388 287164 106452
rect 285628 106252 285692 106316
rect 233924 106116 233988 106180
rect 214420 105300 214484 105364
rect 285812 103124 285876 103188
rect 172100 102172 172164 102236
rect 230428 102308 230492 102372
rect 233740 102172 233804 102236
rect 268516 102308 268580 102372
rect 291332 100948 291396 101012
rect 268516 100540 268580 100604
rect 281580 99316 281644 99380
rect 229324 98908 229388 98972
rect 265756 97956 265820 98020
rect 268516 97956 268580 98020
rect 279372 97956 279436 98020
rect 268516 97140 268580 97204
rect 229140 97004 229204 97068
rect 227668 95372 227732 95436
rect 228956 95372 229020 95436
rect 250300 95372 250364 95436
rect 279372 94964 279436 95028
rect 94918 94752 94982 94756
rect 94918 94696 94962 94752
rect 94962 94696 94982 94752
rect 94918 94692 94982 94696
rect 104302 94752 104366 94756
rect 104302 94696 104346 94752
rect 104346 94696 104366 94752
rect 104302 94692 104366 94696
rect 116678 94752 116742 94756
rect 116678 94696 116730 94752
rect 116730 94696 116742 94752
rect 116678 94692 116742 94696
rect 120622 94752 120686 94756
rect 120622 94696 120630 94752
rect 120630 94696 120686 94752
rect 120622 94692 120686 94696
rect 133134 94752 133198 94756
rect 133134 94696 133142 94752
rect 133142 94696 133198 94752
rect 133134 94692 133198 94696
rect 151766 94752 151830 94756
rect 151766 94696 151782 94752
rect 151782 94696 151830 94752
rect 151766 94692 151830 94696
rect 214420 93740 214484 93804
rect 85620 93528 85684 93532
rect 85620 93472 85670 93528
rect 85670 93472 85684 93528
rect 85620 93468 85684 93472
rect 107700 93528 107764 93532
rect 107700 93472 107750 93528
rect 107750 93472 107764 93528
rect 107700 93468 107764 93472
rect 115796 93528 115860 93532
rect 115796 93472 115846 93528
rect 115846 93472 115860 93528
rect 115796 93468 115860 93472
rect 122052 93528 122116 93532
rect 122052 93472 122102 93528
rect 122102 93472 122116 93528
rect 122052 93468 122116 93472
rect 281580 93468 281644 93532
rect 103284 93196 103348 93260
rect 110092 93196 110156 93260
rect 84332 92380 84396 92444
rect 88012 92440 88076 92444
rect 88012 92384 88062 92440
rect 88062 92384 88076 92440
rect 88012 92380 88076 92384
rect 98132 92380 98196 92444
rect 99972 92440 100036 92444
rect 99972 92384 100022 92440
rect 100022 92384 100036 92440
rect 99972 92380 100036 92384
rect 105676 92440 105740 92444
rect 105676 92384 105726 92440
rect 105726 92384 105740 92440
rect 105676 92380 105740 92384
rect 106780 92440 106844 92444
rect 106780 92384 106830 92440
rect 106830 92384 106844 92440
rect 106780 92380 106844 92384
rect 113036 92380 113100 92444
rect 120212 92440 120276 92444
rect 120212 92384 120262 92440
rect 120262 92384 120276 92440
rect 120212 92380 120276 92384
rect 123156 92440 123220 92444
rect 123156 92384 123206 92440
rect 123206 92384 123220 92440
rect 123156 92380 123220 92384
rect 124076 92440 124140 92444
rect 124076 92384 124126 92440
rect 124126 92384 124140 92440
rect 124076 92380 124140 92384
rect 125364 92440 125428 92444
rect 125364 92384 125414 92440
rect 125414 92384 125428 92440
rect 125364 92380 125428 92384
rect 134380 92440 134444 92444
rect 134380 92384 134430 92440
rect 134430 92384 134444 92440
rect 134380 92380 134444 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 109172 92244 109236 92308
rect 118004 92108 118068 92172
rect 168236 92244 168300 92308
rect 101812 91760 101876 91764
rect 101812 91704 101862 91760
rect 101862 91704 101876 91760
rect 101812 91700 101876 91704
rect 125732 91700 125796 91764
rect 112300 91564 112364 91628
rect 119292 91564 119356 91628
rect 136036 91564 136100 91628
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 98500 91292 98564 91356
rect 100892 91292 100956 91356
rect 113220 91292 113284 91356
rect 115428 91292 115492 91356
rect 126468 91292 126532 91356
rect 74764 91156 74828 91220
rect 86724 91156 86788 91220
rect 88932 91156 88996 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 93900 91156 93964 91220
rect 96292 91156 96356 91220
rect 96660 91156 96724 91220
rect 97212 91156 97276 91220
rect 99052 91156 99116 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 104572 91156 104636 91220
rect 105492 91156 105556 91220
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111196 91156 111260 91220
rect 111932 91156 111996 91220
rect 114324 91216 114388 91220
rect 114324 91160 114374 91216
rect 114374 91160 114388 91216
rect 114324 91156 114388 91160
rect 114876 91156 114940 91220
rect 117084 91156 117148 91220
rect 118188 91216 118252 91220
rect 118188 91160 118238 91216
rect 118238 91160 118252 91216
rect 118188 91156 118252 91160
rect 119660 91216 119724 91220
rect 119660 91160 119710 91216
rect 119710 91160 119724 91216
rect 119660 91156 119724 91160
rect 121684 91156 121748 91220
rect 124444 91156 124508 91220
rect 126652 91216 126716 91220
rect 126652 91160 126702 91216
rect 126702 91160 126716 91216
rect 126652 91156 126716 91160
rect 127572 91156 127636 91220
rect 129412 91216 129476 91220
rect 129412 91160 129462 91216
rect 129462 91160 129476 91216
rect 129412 91156 129476 91160
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 151676 91216 151740 91220
rect 151676 91160 151726 91216
rect 151726 91160 151740 91216
rect 151676 91156 151740 91160
rect 172100 91020 172164 91084
rect 169156 88164 169220 88228
rect 57836 86804 57900 86868
rect 170444 86668 170508 86732
rect 166212 86532 166276 86596
rect 173204 84084 173268 84148
rect 166396 83948 166460 84012
rect 168972 78508 169036 78572
rect 170260 77148 170324 77212
rect 258764 73748 258828 73812
rect 264100 72388 264164 72452
rect 62988 69532 63052 69596
rect 239260 64092 239324 64156
rect 255820 62732 255884 62796
rect 254532 51716 254596 51780
rect 265756 43420 265820 43484
rect 257292 40564 257356 40628
rect 258580 30908 258644 30972
rect 262812 25468 262876 25532
rect 227668 24788 227732 24852
rect 262076 24108 262140 24172
rect 228220 19892 228284 19956
rect 232452 11596 232516 11660
rect 242020 4796 242084 4860
rect 295932 3844 295996 3908
rect 302740 3844 302804 3908
rect 298692 3572 298756 3636
rect 240364 3436 240428 3500
rect 244228 3436 244292 3500
rect 245700 3436 245764 3500
rect 248460 3436 248524 3500
rect 249748 3436 249812 3500
rect 251220 3436 251284 3500
rect 252508 3436 252572 3500
rect 255268 3436 255332 3500
rect 259500 3496 259564 3500
rect 259500 3440 259514 3496
rect 259514 3440 259564 3496
rect 259500 3436 259564 3440
rect 288388 3436 288452 3500
rect 291148 3436 291212 3500
rect 292620 3436 292684 3500
rect 295380 3436 295444 3500
rect 299612 3436 299676 3500
rect 304948 3436 305012 3500
rect 249012 3300 249076 3364
rect 268332 3300 268396 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 44035 531996 44101 531997
rect 44035 531932 44036 531996
rect 44100 531932 44101 531996
rect 44035 531931 44101 531932
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 44038 434621 44098 531931
rect 45234 514894 45854 550338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48083 532132 48149 532133
rect 48083 532068 48084 532132
rect 48148 532068 48149 532132
rect 48083 532067 48149 532068
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 44035 434620 44101 434621
rect 44035 434556 44036 434620
rect 44100 434556 44101 434620
rect 44035 434555 44101 434556
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 44038 339421 44098 434555
rect 45234 406894 45854 442338
rect 48086 433261 48146 532067
rect 48954 518614 49574 554058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 57835 586396 57901 586397
rect 57835 586332 57836 586396
rect 57900 586332 57901 586396
rect 57835 586331 57901 586332
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 53603 532268 53669 532269
rect 53603 532204 53604 532268
rect 53668 532204 53669 532268
rect 53603 532203 53669 532204
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 50843 494868 50909 494869
rect 50843 494804 50844 494868
rect 50908 494804 50909 494868
rect 50843 494803 50909 494804
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48083 433260 48149 433261
rect 48083 433196 48084 433260
rect 48148 433196 48149 433260
rect 48083 433195 48149 433196
rect 48083 430676 48149 430677
rect 48083 430612 48084 430676
rect 48148 430612 48149 430676
rect 48083 430611 48149 430612
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 44035 339420 44101 339421
rect 44035 339356 44036 339420
rect 44100 339356 44101 339420
rect 44035 339355 44101 339356
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 334894 45854 370338
rect 48086 340781 48146 430611
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 50846 399533 50906 494803
rect 52315 492692 52381 492693
rect 52315 492628 52316 492692
rect 52380 492628 52381 492692
rect 52315 492627 52381 492628
rect 50843 399532 50909 399533
rect 50843 399468 50844 399532
rect 50908 399468 50909 399532
rect 50843 399467 50909 399468
rect 52318 398037 52378 492627
rect 53051 492012 53117 492013
rect 53051 491948 53052 492012
rect 53116 491948 53117 492012
rect 53051 491947 53117 491948
rect 52315 398036 52381 398037
rect 52315 397972 52316 398036
rect 52380 397972 52381 398036
rect 52315 397971 52381 397972
rect 53054 387565 53114 491947
rect 53606 441149 53666 532203
rect 55794 525454 56414 560898
rect 57838 537573 57898 586331
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 57835 537572 57901 537573
rect 57835 537508 57836 537572
rect 57900 537508 57901 537572
rect 57835 537507 57901 537508
rect 57835 537436 57901 537437
rect 57835 537372 57836 537436
rect 57900 537372 57901 537436
rect 57835 537371 57901 537372
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55075 489156 55141 489157
rect 55075 489092 55076 489156
rect 55140 489092 55141 489156
rect 55075 489091 55141 489092
rect 55794 489134 56414 489218
rect 53603 441148 53669 441149
rect 53603 441084 53604 441148
rect 53668 441084 53669 441148
rect 53603 441083 53669 441084
rect 55078 438837 55138 489091
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55075 438836 55141 438837
rect 55075 438772 55076 438836
rect 55140 438772 55141 438836
rect 55075 438771 55141 438772
rect 55794 417454 56414 452898
rect 57838 437477 57898 537371
rect 59514 529174 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66115 577148 66181 577149
rect 66115 577084 66116 577148
rect 66180 577084 66181 577148
rect 66115 577083 66181 577084
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 61883 561916 61949 561917
rect 61883 561852 61884 561916
rect 61948 561852 61949 561916
rect 61883 561851 61949 561852
rect 60595 560556 60661 560557
rect 60595 560492 60596 560556
rect 60660 560492 60661 560556
rect 60595 560491 60661 560492
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59123 490516 59189 490517
rect 59123 490452 59124 490516
rect 59188 490452 59189 490516
rect 59123 490451 59189 490452
rect 59126 441013 59186 490451
rect 59514 457174 60134 492618
rect 60598 461005 60658 560491
rect 61699 477460 61765 477461
rect 61699 477396 61700 477460
rect 61764 477396 61765 477460
rect 61699 477395 61765 477396
rect 60595 461004 60661 461005
rect 60595 460940 60596 461004
rect 60660 460940 60661 461004
rect 60595 460939 60661 460940
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59123 441012 59189 441013
rect 59123 440948 59124 441012
rect 59188 440948 59189 441012
rect 59123 440947 59189 440948
rect 57835 437476 57901 437477
rect 57835 437412 57836 437476
rect 57900 437412 57901 437476
rect 57835 437411 57901 437412
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 53603 399668 53669 399669
rect 53603 399604 53604 399668
rect 53668 399604 53669 399668
rect 53603 399603 53669 399604
rect 53051 387564 53117 387565
rect 53051 387500 53052 387564
rect 53116 387500 53117 387564
rect 53051 387499 53117 387500
rect 52315 377772 52381 377773
rect 52315 377708 52316 377772
rect 52380 377708 52381 377772
rect 52315 377707 52381 377708
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48083 340780 48149 340781
rect 48083 340716 48084 340780
rect 48148 340716 48149 340780
rect 48083 340715 48149 340716
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 338614 49574 374058
rect 52318 339693 52378 377707
rect 52315 339692 52381 339693
rect 52315 339628 52316 339692
rect 52380 339628 52381 339692
rect 52315 339627 52381 339628
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 53606 333981 53666 399603
rect 55794 381454 56414 416898
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 57835 391236 57901 391237
rect 57835 391172 57836 391236
rect 57900 391172 57901 391236
rect 57835 391171 57901 391172
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55075 370564 55141 370565
rect 55075 370500 55076 370564
rect 55140 370500 55141 370564
rect 55075 370499 55141 370500
rect 53603 333980 53669 333981
rect 53603 333916 53604 333980
rect 53668 333916 53669 333980
rect 53603 333915 53669 333916
rect 55078 330445 55138 370499
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55075 330444 55141 330445
rect 55075 330380 55076 330444
rect 55140 330380 55141 330444
rect 55075 330379 55141 330380
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 55794 309454 56414 344898
rect 57838 337925 57898 391171
rect 59123 389196 59189 389197
rect 59123 389132 59124 389196
rect 59188 389132 59189 389196
rect 59123 389131 59189 389132
rect 57835 337924 57901 337925
rect 57835 337860 57836 337924
rect 57900 337860 57901 337924
rect 57835 337859 57901 337860
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 50843 265164 50909 265165
rect 50843 265100 50844 265164
rect 50908 265100 50909 265164
rect 50843 265099 50909 265100
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 50846 225589 50906 265099
rect 55794 237454 56414 272898
rect 57835 251428 57901 251429
rect 57835 251364 57836 251428
rect 57900 251364 57901 251428
rect 57835 251363 57901 251364
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 50843 225588 50909 225589
rect 50843 225524 50844 225588
rect 50908 225524 50909 225588
rect 50843 225523 50909 225524
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 57838 86869 57898 251363
rect 59126 240413 59186 389131
rect 59514 385174 60134 420618
rect 61702 401709 61762 477395
rect 61886 463589 61946 561851
rect 62987 548044 63053 548045
rect 62987 547980 62988 548044
rect 63052 547980 63053 548044
rect 62987 547979 63053 547980
rect 61883 463588 61949 463589
rect 61883 463524 61884 463588
rect 61948 463524 61949 463588
rect 61883 463523 61949 463524
rect 62990 447813 63050 547979
rect 63234 532894 63854 568338
rect 64643 565860 64709 565861
rect 64643 565796 64644 565860
rect 64708 565796 64709 565860
rect 64643 565795 64709 565796
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 64646 467805 64706 565795
rect 65931 480588 65997 480589
rect 65931 480524 65932 480588
rect 65996 480524 65997 480588
rect 65931 480523 65997 480524
rect 64643 467804 64709 467805
rect 64643 467740 64644 467804
rect 64708 467740 64709 467804
rect 64643 467739 64709 467740
rect 64646 467261 64706 467739
rect 64643 467260 64709 467261
rect 64643 467196 64644 467260
rect 64708 467196 64709 467260
rect 64643 467195 64709 467196
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 62987 447812 63053 447813
rect 62987 447748 62988 447812
rect 63052 447748 63053 447812
rect 62987 447747 63053 447748
rect 61883 442916 61949 442917
rect 61883 442852 61884 442916
rect 61948 442852 61949 442916
rect 61883 442851 61949 442852
rect 61886 441693 61946 442851
rect 61883 441692 61949 441693
rect 61883 441628 61884 441692
rect 61948 441628 61949 441692
rect 61883 441627 61949 441628
rect 61699 401708 61765 401709
rect 61699 401644 61700 401708
rect 61764 401644 61765 401708
rect 61699 401643 61765 401644
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 61699 355332 61765 355333
rect 61699 355268 61700 355332
rect 61764 355268 61765 355332
rect 61699 355267 61765 355268
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 61331 337924 61397 337925
rect 61331 337860 61332 337924
rect 61396 337860 61397 337924
rect 61331 337859 61397 337860
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59123 240412 59189 240413
rect 59123 240348 59124 240412
rect 59188 240348 59189 240412
rect 59123 240347 59189 240348
rect 59514 205174 60134 240618
rect 61334 238509 61394 337859
rect 61702 323781 61762 355267
rect 61886 342277 61946 441627
rect 63234 424894 63854 460338
rect 65934 440333 65994 480523
rect 66118 478549 66178 577083
rect 66954 572614 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 584000 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 584000 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 584000 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 584000 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 584000 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 584000 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 584000 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 584000 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 111011 702540 111077 702541
rect 111011 702476 111012 702540
rect 111076 702476 111077 702540
rect 111011 702475 111077 702476
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 76576 579454 76896 579486
rect 76576 579218 76618 579454
rect 76854 579218 76896 579454
rect 76576 579134 76896 579218
rect 76576 578898 76618 579134
rect 76854 578898 76896 579134
rect 76576 578866 76896 578898
rect 87840 579454 88160 579486
rect 87840 579218 87882 579454
rect 88118 579218 88160 579454
rect 87840 579134 88160 579218
rect 87840 578898 87882 579134
rect 88118 578898 88160 579134
rect 87840 578866 88160 578898
rect 99104 579454 99424 579486
rect 99104 579218 99146 579454
rect 99382 579218 99424 579454
rect 99104 579134 99424 579218
rect 99104 578898 99146 579134
rect 99382 578898 99424 579134
rect 99104 578866 99424 578898
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66667 571844 66733 571845
rect 66667 571780 66668 571844
rect 66732 571780 66733 571844
rect 66667 571779 66733 571780
rect 66115 478548 66181 478549
rect 66115 478484 66116 478548
rect 66180 478484 66181 478548
rect 66115 478483 66181 478484
rect 65931 440332 65997 440333
rect 65931 440268 65932 440332
rect 65996 440268 65997 440332
rect 65931 440267 65997 440268
rect 64643 439516 64709 439517
rect 64643 439452 64644 439516
rect 64708 439452 64709 439516
rect 64643 439451 64709 439452
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 62987 377364 63053 377365
rect 62987 377300 62988 377364
rect 63052 377300 63053 377364
rect 62987 377299 63053 377300
rect 61883 342276 61949 342277
rect 61883 342212 61884 342276
rect 61948 342212 61949 342276
rect 61883 342211 61949 342212
rect 61699 323780 61765 323781
rect 61699 323716 61700 323780
rect 61764 323716 61765 323780
rect 61699 323715 61765 323716
rect 61515 253876 61581 253877
rect 61515 253812 61516 253876
rect 61580 253812 61581 253876
rect 61515 253811 61581 253812
rect 61331 238508 61397 238509
rect 61331 238444 61332 238508
rect 61396 238444 61397 238508
rect 61331 238443 61397 238444
rect 61518 235245 61578 253811
rect 61515 235244 61581 235245
rect 61515 235180 61516 235244
rect 61580 235180 61581 235244
rect 61515 235179 61581 235180
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 57835 86868 57901 86869
rect 57835 86804 57836 86868
rect 57900 86804 57901 86868
rect 57835 86803 57901 86804
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 61174 60134 96618
rect 62990 69597 63050 377299
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 64646 340781 64706 439451
rect 66118 400349 66178 478483
rect 66670 474061 66730 571779
rect 66954 536614 67574 572058
rect 68875 570348 68941 570349
rect 68875 570284 68876 570348
rect 68940 570284 68941 570348
rect 68875 570283 68941 570284
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66667 474060 66733 474061
rect 66667 473996 66668 474060
rect 66732 473996 66733 474060
rect 66667 473995 66733 473996
rect 66670 473789 66730 473995
rect 66667 473788 66733 473789
rect 66667 473724 66668 473788
rect 66732 473724 66733 473788
rect 66667 473723 66733 473724
rect 66954 464614 67574 500058
rect 68691 482628 68757 482629
rect 68691 482564 68692 482628
rect 68756 482564 68757 482628
rect 68691 482563 68757 482564
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 68694 438973 68754 482563
rect 68878 471069 68938 570283
rect 106411 564500 106477 564501
rect 106411 564436 106412 564500
rect 106476 564436 106477 564500
rect 106411 564435 106477 564436
rect 105491 561916 105557 561917
rect 105491 561852 105492 561916
rect 105556 561852 105557 561916
rect 105491 561851 105557 561852
rect 82208 561454 82528 561486
rect 82208 561218 82250 561454
rect 82486 561218 82528 561454
rect 82208 561134 82528 561218
rect 82208 560898 82250 561134
rect 82486 560898 82528 561134
rect 82208 560866 82528 560898
rect 93472 561454 93792 561486
rect 93472 561218 93514 561454
rect 93750 561218 93792 561454
rect 93472 561134 93792 561218
rect 93472 560898 93514 561134
rect 93750 560898 93792 561134
rect 93472 560866 93792 560898
rect 105494 547890 105554 561851
rect 104942 547830 105554 547890
rect 76576 543454 76896 543486
rect 76576 543218 76618 543454
rect 76854 543218 76896 543454
rect 76576 543134 76896 543218
rect 76576 542898 76618 543134
rect 76854 542898 76896 543134
rect 76576 542866 76896 542898
rect 87840 543454 88160 543486
rect 87840 543218 87882 543454
rect 88118 543218 88160 543454
rect 87840 543134 88160 543218
rect 87840 542898 87882 543134
rect 88118 542898 88160 543134
rect 87840 542866 88160 542898
rect 99104 543454 99424 543486
rect 99104 543218 99146 543454
rect 99382 543218 99424 543454
rect 99104 543134 99424 543218
rect 99104 542898 99146 543134
rect 99382 542898 99424 543134
rect 99104 542866 99424 542898
rect 70347 538796 70413 538797
rect 70347 538732 70348 538796
rect 70412 538732 70413 538796
rect 70347 538731 70413 538732
rect 69059 486572 69125 486573
rect 69059 486508 69060 486572
rect 69124 486508 69125 486572
rect 69059 486507 69125 486508
rect 68875 471068 68941 471069
rect 68875 471004 68876 471068
rect 68940 471004 68941 471068
rect 68875 471003 68941 471004
rect 68691 438972 68757 438973
rect 68691 438908 68692 438972
rect 68756 438908 68757 438972
rect 68691 438907 68757 438908
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66115 400348 66181 400349
rect 66115 400284 66116 400348
rect 66180 400284 66181 400348
rect 66115 400283 66181 400284
rect 66118 384845 66178 400283
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66115 384844 66181 384845
rect 66115 384780 66116 384844
rect 66180 384780 66181 384844
rect 66115 384779 66181 384780
rect 65379 376004 65445 376005
rect 65379 375940 65380 376004
rect 65444 375940 65445 376004
rect 65379 375939 65445 375940
rect 64643 340780 64709 340781
rect 64643 340716 64644 340780
rect 64708 340716 64709 340780
rect 64643 340715 64709 340716
rect 65382 323645 65442 375939
rect 66954 356614 67574 392058
rect 68878 377229 68938 471003
rect 69062 439517 69122 486507
rect 70350 484669 70410 538731
rect 103651 538116 103717 538117
rect 103651 538052 103652 538116
rect 103716 538052 103717 538116
rect 103651 538051 103717 538052
rect 73794 507454 74414 538000
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 492000 74414 506898
rect 77514 511174 78134 538000
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 492000 78134 510618
rect 81234 514894 81854 538000
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 492000 81854 514338
rect 84954 518614 85574 538000
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 492000 85574 518058
rect 91794 525454 92414 538000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 492000 92414 524898
rect 95514 529174 96134 538000
rect 98499 537436 98565 537437
rect 98499 537372 98500 537436
rect 98564 537372 98565 537436
rect 98499 537371 98565 537372
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 492000 96134 492618
rect 98502 489973 98562 537371
rect 99234 532894 99854 538000
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 492000 99854 496338
rect 102954 536614 103574 538000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 99419 490652 99485 490653
rect 99419 490588 99420 490652
rect 99484 490588 99485 490652
rect 99419 490587 99485 490588
rect 98499 489972 98565 489973
rect 98499 489908 98500 489972
rect 98564 489908 98565 489972
rect 98499 489907 98565 489908
rect 70347 484668 70413 484669
rect 70347 484604 70348 484668
rect 70412 484604 70413 484668
rect 70347 484603 70413 484604
rect 75576 471454 75896 471486
rect 75576 471218 75618 471454
rect 75854 471218 75896 471454
rect 75576 471134 75896 471218
rect 75576 470898 75618 471134
rect 75854 470898 75896 471134
rect 75576 470866 75896 470898
rect 84840 471454 85160 471486
rect 84840 471218 84882 471454
rect 85118 471218 85160 471454
rect 84840 471134 85160 471218
rect 84840 470898 84882 471134
rect 85118 470898 85160 471134
rect 84840 470866 85160 470898
rect 94104 471454 94424 471486
rect 94104 471218 94146 471454
rect 94382 471218 94424 471454
rect 94104 471134 94424 471218
rect 94104 470898 94146 471134
rect 94382 470898 94424 471134
rect 94104 470866 94424 470898
rect 80208 453454 80528 453486
rect 80208 453218 80250 453454
rect 80486 453218 80528 453454
rect 80208 453134 80528 453218
rect 80208 452898 80250 453134
rect 80486 452898 80528 453134
rect 80208 452866 80528 452898
rect 89472 453454 89792 453486
rect 89472 453218 89514 453454
rect 89750 453218 89792 453454
rect 89472 453134 89792 453218
rect 89472 452898 89514 453134
rect 89750 452898 89792 453134
rect 89472 452866 89792 452898
rect 99051 441148 99117 441149
rect 99051 441084 99052 441148
rect 99116 441084 99117 441148
rect 99051 441083 99117 441084
rect 69059 439516 69125 439517
rect 69059 439452 69060 439516
rect 69124 439452 69125 439516
rect 69059 439451 69125 439452
rect 70347 437748 70413 437749
rect 70347 437684 70348 437748
rect 70412 437684 70413 437748
rect 70347 437683 70413 437684
rect 69979 383212 70045 383213
rect 69979 383148 69980 383212
rect 70044 383210 70045 383212
rect 70350 383210 70410 437683
rect 73794 435454 74414 438000
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 388000 74414 398898
rect 77514 403174 78134 438000
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 388000 78134 402618
rect 81234 406894 81854 438000
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 388000 81854 406338
rect 84954 410614 85574 438000
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 388000 85574 410058
rect 91794 417454 92414 438000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 388000 92414 416898
rect 95514 421174 96134 438000
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 388000 96134 420618
rect 99054 388381 99114 441083
rect 99422 439109 99482 490587
rect 101995 489972 102061 489973
rect 101995 489908 101996 489972
rect 102060 489908 102061 489972
rect 101995 489907 102061 489908
rect 99971 466308 100037 466309
rect 99971 466244 99972 466308
rect 100036 466244 100037 466308
rect 99971 466243 100037 466244
rect 99419 439108 99485 439109
rect 99419 439044 99420 439108
rect 99484 439044 99485 439108
rect 99419 439043 99485 439044
rect 99974 438701 100034 466243
rect 99971 438700 100037 438701
rect 99971 438636 99972 438700
rect 100036 438636 100037 438700
rect 99971 438635 100037 438636
rect 99234 424894 99854 438000
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 101998 393413 102058 489907
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102731 461548 102797 461549
rect 102731 461484 102732 461548
rect 102796 461484 102797 461548
rect 102731 461483 102797 461484
rect 102734 440197 102794 461483
rect 102731 440196 102797 440197
rect 102731 440132 102732 440196
rect 102796 440132 102797 440196
rect 102731 440131 102797 440132
rect 102954 428614 103574 464058
rect 103654 460950 103714 538051
rect 104942 471205 105002 547830
rect 106414 478141 106474 564435
rect 107699 557700 107765 557701
rect 107699 557636 107700 557700
rect 107764 557636 107765 557700
rect 107699 557635 107765 557636
rect 106411 478140 106477 478141
rect 106411 478076 106412 478140
rect 106476 478076 106477 478140
rect 106411 478075 106477 478076
rect 104939 471204 105005 471205
rect 104939 471140 104940 471204
rect 105004 471140 105005 471204
rect 104939 471139 105005 471140
rect 105491 467940 105557 467941
rect 105491 467876 105492 467940
rect 105556 467876 105557 467940
rect 105491 467875 105557 467876
rect 103654 460890 103898 460950
rect 103838 445773 103898 460890
rect 103835 445772 103901 445773
rect 103835 445708 103836 445772
rect 103900 445708 103901 445772
rect 103835 445707 103901 445708
rect 103838 444413 103898 445707
rect 103835 444412 103901 444413
rect 103835 444348 103836 444412
rect 103900 444348 103901 444412
rect 103835 444347 103901 444348
rect 105494 435981 105554 467875
rect 107702 465765 107762 557635
rect 107883 546820 107949 546821
rect 107883 546756 107884 546820
rect 107948 546756 107949 546820
rect 107883 546755 107949 546756
rect 107699 465764 107765 465765
rect 107699 465700 107700 465764
rect 107764 465700 107765 465764
rect 107699 465699 107765 465700
rect 107886 456109 107946 546755
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 111014 540157 111074 702475
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 115979 584084 116045 584085
rect 115979 584020 115980 584084
rect 116044 584020 116045 584084
rect 115979 584019 116045 584020
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111747 578236 111813 578237
rect 111747 578172 111748 578236
rect 111812 578172 111813 578236
rect 111747 578171 111813 578172
rect 111011 540156 111077 540157
rect 111011 540092 111012 540156
rect 111076 540092 111077 540156
rect 111011 540091 111077 540092
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109539 491468 109605 491469
rect 109539 491404 109540 491468
rect 109604 491404 109605 491468
rect 109539 491403 109605 491404
rect 107883 456108 107949 456109
rect 107883 456044 107884 456108
rect 107948 456044 107949 456108
rect 107883 456043 107949 456044
rect 105491 435980 105557 435981
rect 105491 435916 105492 435980
rect 105556 435916 105557 435980
rect 105491 435915 105557 435916
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 101995 393412 102061 393413
rect 101995 393348 101996 393412
rect 102060 393348 102061 393412
rect 101995 393347 102061 393348
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99051 388380 99117 388381
rect 99051 388316 99052 388380
rect 99116 388316 99117 388380
rect 99051 388315 99117 388316
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 388000 99854 388338
rect 102954 392614 103574 428058
rect 109542 401301 109602 491403
rect 109794 471454 110414 506898
rect 111011 491332 111077 491333
rect 111011 491268 111012 491332
rect 111076 491268 111077 491332
rect 111011 491267 111077 491268
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109539 401300 109605 401301
rect 109539 401236 109540 401300
rect 109604 401236 109605 401300
rect 109539 401235 109605 401236
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 388000 103574 392058
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 388000 110414 398898
rect 111014 389197 111074 491267
rect 111750 485077 111810 578171
rect 113514 547174 114134 582618
rect 114507 581772 114573 581773
rect 114507 581708 114508 581772
rect 114572 581708 114573 581772
rect 114507 581707 114573 581708
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 114510 536077 114570 581707
rect 114507 536076 114573 536077
rect 114507 536012 114508 536076
rect 114572 536012 114573 536076
rect 114507 536011 114573 536012
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111747 485076 111813 485077
rect 111747 485012 111748 485076
rect 111812 485012 111813 485076
rect 111747 485011 111813 485012
rect 112299 478956 112365 478957
rect 112299 478892 112300 478956
rect 112364 478892 112365 478956
rect 112299 478891 112365 478892
rect 111011 389196 111077 389197
rect 111011 389132 111012 389196
rect 111076 389132 111077 389196
rect 111011 389131 111077 389132
rect 70531 387700 70597 387701
rect 70531 387636 70532 387700
rect 70596 387636 70597 387700
rect 70531 387635 70597 387636
rect 70044 383150 70410 383210
rect 70044 383148 70045 383150
rect 69979 383147 70045 383148
rect 69059 380356 69125 380357
rect 69059 380292 69060 380356
rect 69124 380292 69125 380356
rect 69059 380291 69125 380292
rect 68875 377228 68941 377229
rect 68875 377164 68876 377228
rect 68940 377164 68941 377228
rect 68875 377163 68941 377164
rect 68875 372876 68941 372877
rect 68875 372812 68876 372876
rect 68940 372812 68941 372876
rect 68875 372811 68941 372812
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 65379 323644 65445 323645
rect 65379 323580 65380 323644
rect 65444 323580 65445 323644
rect 65379 323579 65445 323580
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 68878 316709 68938 372811
rect 68875 316708 68941 316709
rect 68875 316644 68876 316708
rect 68940 316644 68941 316708
rect 68875 316643 68941 316644
rect 69062 305693 69122 380291
rect 70534 377773 70594 387635
rect 112302 385389 112362 478891
rect 113514 475174 114134 510618
rect 115982 490109 116042 584019
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 118739 578916 118805 578917
rect 118739 578852 118740 578916
rect 118804 578852 118805 578916
rect 118739 578851 118805 578852
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 115979 490108 116045 490109
rect 115979 490044 115980 490108
rect 116044 490044 116045 490108
rect 115979 490043 116045 490044
rect 115982 489930 116042 490043
rect 115982 489870 116594 489930
rect 115795 488476 115861 488477
rect 115795 488412 115796 488476
rect 115860 488412 115861 488476
rect 115795 488411 115861 488412
rect 115611 485076 115677 485077
rect 115611 485012 115612 485076
rect 115676 485012 115677 485076
rect 115611 485011 115677 485012
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 115614 458285 115674 485011
rect 115798 459645 115858 488411
rect 116534 463589 116594 489870
rect 117234 478894 117854 514338
rect 118742 495549 118802 578851
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118739 495548 118805 495549
rect 118739 495484 118740 495548
rect 118804 495484 118805 495548
rect 118739 495483 118805 495484
rect 118742 495005 118802 495483
rect 118739 495004 118805 495005
rect 118739 494940 118740 495004
rect 118804 494940 118805 495004
rect 118739 494939 118805 494940
rect 118923 486436 118989 486437
rect 118923 486372 118924 486436
rect 118988 486372 118989 486436
rect 118923 486371 118989 486372
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117083 477460 117149 477461
rect 117083 477396 117084 477460
rect 117148 477396 117149 477460
rect 117083 477395 117149 477396
rect 116531 463588 116597 463589
rect 116531 463524 116532 463588
rect 116596 463524 116597 463588
rect 116531 463523 116597 463524
rect 115795 459644 115861 459645
rect 115795 459580 115796 459644
rect 115860 459580 115861 459644
rect 115795 459579 115861 459580
rect 115611 458284 115677 458285
rect 115611 458220 115612 458284
rect 115676 458220 115677 458284
rect 115611 458219 115677 458220
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 388000 114134 402618
rect 115979 394092 116045 394093
rect 115979 394028 115980 394092
rect 116044 394028 116045 394092
rect 115979 394027 116045 394028
rect 115427 387836 115493 387837
rect 115427 387772 115428 387836
rect 115492 387772 115493 387836
rect 115427 387771 115493 387772
rect 112299 385388 112365 385389
rect 112299 385324 112300 385388
rect 112364 385324 112365 385388
rect 112299 385323 112365 385324
rect 115430 384573 115490 387771
rect 115427 384572 115493 384573
rect 115427 384508 115428 384572
rect 115492 384508 115493 384572
rect 115427 384507 115493 384508
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 70531 377772 70597 377773
rect 70531 377708 70532 377772
rect 70596 377708 70597 377772
rect 70531 377707 70597 377708
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 115982 357373 116042 394027
rect 117086 372741 117146 477395
rect 117234 442894 117854 478338
rect 118739 475964 118805 475965
rect 118739 475900 118740 475964
rect 118804 475900 118805 475964
rect 118739 475899 118805 475900
rect 118003 474060 118069 474061
rect 118003 473996 118004 474060
rect 118068 473996 118069 474060
rect 118003 473995 118069 473996
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 388000 117854 406338
rect 117083 372740 117149 372741
rect 117083 372676 117084 372740
rect 117148 372676 117149 372740
rect 117083 372675 117149 372676
rect 118006 371381 118066 473995
rect 118003 371380 118069 371381
rect 118003 371316 118004 371380
rect 118068 371316 118069 371380
rect 118003 371315 118069 371316
rect 118742 368661 118802 475899
rect 118926 381581 118986 486371
rect 120954 482614 121574 518058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 124443 494732 124509 494733
rect 124443 494668 124444 494732
rect 124508 494668 124509 494732
rect 124443 494667 124509 494668
rect 122787 489972 122853 489973
rect 122787 489970 122788 489972
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120763 387836 120829 387837
rect 120763 387772 120764 387836
rect 120828 387772 120829 387836
rect 120763 387771 120829 387772
rect 118923 381580 118989 381581
rect 118923 381516 118924 381580
rect 118988 381516 118989 381580
rect 118923 381515 118989 381516
rect 118926 381037 118986 381515
rect 118923 381036 118989 381037
rect 118923 380972 118924 381036
rect 118988 380972 118989 381036
rect 118923 380971 118989 380972
rect 118739 368660 118805 368661
rect 118739 368596 118740 368660
rect 118804 368596 118805 368660
rect 118739 368595 118805 368596
rect 120766 366349 120826 387771
rect 120954 374614 121574 410058
rect 122606 489910 122788 489970
rect 121683 390692 121749 390693
rect 121683 390628 121684 390692
rect 121748 390628 121749 390692
rect 121683 390627 121749 390628
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120763 366348 120829 366349
rect 120763 366284 120764 366348
rect 120828 366284 120829 366348
rect 120763 366283 120829 366284
rect 115979 357372 116045 357373
rect 115979 357308 115980 357372
rect 116044 357308 116045 357372
rect 115979 357307 116045 357308
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 70347 342956 70413 342957
rect 70347 342892 70348 342956
rect 70412 342892 70413 342956
rect 70347 342891 70413 342892
rect 70350 336021 70410 342891
rect 70531 341052 70597 341053
rect 70531 340988 70532 341052
rect 70596 340988 70597 341052
rect 70531 340987 70597 340988
rect 70534 336157 70594 340987
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 70531 336156 70597 336157
rect 70531 336092 70532 336156
rect 70596 336092 70597 336156
rect 70531 336091 70597 336092
rect 70347 336020 70413 336021
rect 70347 335956 70348 336020
rect 70412 335956 70413 336020
rect 70347 335955 70413 335956
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 69059 305692 69125 305693
rect 69059 305628 69060 305692
rect 69124 305628 69125 305692
rect 69059 305627 69125 305628
rect 70899 304196 70965 304197
rect 70899 304132 70900 304196
rect 70964 304132 70965 304196
rect 70899 304131 70965 304132
rect 70902 287070 70962 304131
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 331174 114134 338000
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 334894 117854 338000
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 120954 302614 121574 338058
rect 121686 314261 121746 390627
rect 122606 389877 122666 489910
rect 122787 489908 122788 489910
rect 122852 489908 122853 489972
rect 122787 489907 122853 489908
rect 124259 439380 124325 439381
rect 124259 439316 124260 439380
rect 124324 439316 124325 439380
rect 124259 439315 124325 439316
rect 122603 389876 122669 389877
rect 122603 389812 122604 389876
rect 122668 389812 122669 389876
rect 122603 389811 122669 389812
rect 122419 388924 122485 388925
rect 122419 388860 122420 388924
rect 122484 388860 122485 388924
rect 122419 388859 122485 388860
rect 122422 374010 122482 388859
rect 123339 388380 123405 388381
rect 123339 388316 123340 388380
rect 123404 388316 123405 388380
rect 123339 388315 123405 388316
rect 122603 387836 122669 387837
rect 122603 387772 122604 387836
rect 122668 387772 122669 387836
rect 122603 387771 122669 387772
rect 122606 383890 122666 387771
rect 122606 383830 122850 383890
rect 122790 383670 122850 383830
rect 122238 373950 122482 374010
rect 122606 383610 122850 383670
rect 122606 374010 122666 383610
rect 122606 373950 123034 374010
rect 122238 370565 122298 373950
rect 122974 373010 123034 373950
rect 122606 372950 123034 373010
rect 122235 370564 122301 370565
rect 122235 370500 122236 370564
rect 122300 370500 122301 370564
rect 122235 370499 122301 370500
rect 122606 331125 122666 372950
rect 123342 360909 123402 388315
rect 123339 360908 123405 360909
rect 123339 360844 123340 360908
rect 123404 360844 123405 360908
rect 123339 360843 123405 360844
rect 122603 331124 122669 331125
rect 122603 331060 122604 331124
rect 122668 331060 122669 331124
rect 122603 331059 122669 331060
rect 124262 324325 124322 439315
rect 124446 438837 124506 494667
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 124443 438836 124509 438837
rect 124443 438772 124444 438836
rect 124508 438772 124509 438836
rect 124443 438771 124509 438772
rect 125731 438836 125797 438837
rect 125731 438772 125732 438836
rect 125796 438772 125797 438836
rect 125731 438771 125797 438772
rect 124811 356148 124877 356149
rect 124811 356084 124812 356148
rect 124876 356084 124877 356148
rect 124811 356083 124877 356084
rect 124814 341461 124874 356083
rect 124811 341460 124877 341461
rect 124811 341396 124812 341460
rect 124876 341396 124877 341460
rect 124811 341395 124877 341396
rect 124811 337380 124877 337381
rect 124811 337316 124812 337380
rect 124876 337316 124877 337380
rect 124811 337315 124877 337316
rect 124259 324324 124325 324325
rect 124259 324260 124260 324324
rect 124324 324260 124325 324324
rect 124259 324259 124325 324260
rect 121683 314260 121749 314261
rect 121683 314196 121684 314260
rect 121748 314196 121749 314260
rect 121683 314195 121749 314196
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 118739 296036 118805 296037
rect 118739 295972 118740 296036
rect 118804 295972 118805 296036
rect 118739 295971 118805 295972
rect 70534 287010 70962 287070
rect 118742 287070 118802 295971
rect 120954 294000 121574 302058
rect 123339 294268 123405 294269
rect 123339 294204 123340 294268
rect 123404 294204 123405 294268
rect 123339 294203 123405 294204
rect 118742 287010 119354 287070
rect 70534 286789 70594 287010
rect 70531 286788 70597 286789
rect 70531 286724 70532 286788
rect 70596 286724 70597 286788
rect 70531 286723 70597 286724
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66115 276316 66181 276317
rect 66115 276252 66116 276316
rect 66180 276252 66181 276316
rect 66115 276251 66181 276252
rect 65931 250476 65997 250477
rect 65931 250412 65932 250476
rect 65996 250412 65997 250476
rect 65931 250411 65997 250412
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 65934 196621 65994 250411
rect 65931 196620 65997 196621
rect 65931 196556 65932 196620
rect 65996 196556 65997 196620
rect 65931 196555 65997 196556
rect 66118 184245 66178 276251
rect 66954 248614 67574 284058
rect 119294 275637 119354 287010
rect 119291 275636 119357 275637
rect 119291 275572 119292 275636
rect 119356 275572 119357 275636
rect 119291 275571 119357 275572
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 123342 255917 123402 294203
rect 124814 283525 124874 337315
rect 125734 332485 125794 438771
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 133091 445772 133157 445773
rect 133091 445708 133092 445772
rect 133156 445708 133157 445772
rect 133091 445707 133157 445708
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 128675 404972 128741 404973
rect 128675 404970 128676 404972
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 128494 404910 128676 404970
rect 128494 345030 128554 404910
rect 128675 404908 128676 404910
rect 128740 404908 128741 404972
rect 128675 404907 128741 404908
rect 129779 399532 129845 399533
rect 129779 399468 129780 399532
rect 129844 399468 129845 399532
rect 129779 399467 129845 399468
rect 128494 344970 128738 345030
rect 126099 337516 126165 337517
rect 126099 337452 126100 337516
rect 126164 337452 126165 337516
rect 126099 337451 126165 337452
rect 125731 332484 125797 332485
rect 125731 332420 125732 332484
rect 125796 332420 125797 332484
rect 125731 332419 125797 332420
rect 124811 283524 124877 283525
rect 124811 283460 124812 283524
rect 124876 283460 124877 283524
rect 124811 283459 124877 283460
rect 123339 255916 123405 255917
rect 123339 255852 123340 255916
rect 123404 255852 123405 255916
rect 123339 255851 123405 255852
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 126102 253197 126162 337451
rect 127794 309454 128414 344898
rect 128678 338061 128738 344970
rect 128675 338060 128741 338061
rect 128675 337996 128676 338060
rect 128740 337996 128741 338060
rect 128675 337995 128741 337996
rect 129782 328405 129842 399467
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 129779 328404 129845 328405
rect 129779 328340 129780 328404
rect 129844 328340 129845 328404
rect 129779 328339 129845 328340
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 126099 253196 126165 253197
rect 126099 253132 126100 253196
rect 126164 253132 126165 253196
rect 126099 253131 126165 253132
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 70531 248436 70597 248437
rect 70531 248372 70532 248436
rect 70596 248372 70597 248436
rect 70531 248371 70597 248372
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 70534 238770 70594 248371
rect 120027 246532 120093 246533
rect 120027 246468 120028 246532
rect 120092 246468 120093 246532
rect 120027 246467 120093 246468
rect 120030 238770 120090 246467
rect 70534 238710 70962 238770
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66115 184244 66181 184245
rect 66115 184180 66116 184244
rect 66180 184180 66181 184244
rect 66115 184179 66181 184180
rect 66954 176600 67574 212058
rect 70902 180165 70962 238710
rect 119294 238710 120090 238770
rect 119294 238509 119354 238710
rect 119291 238508 119357 238509
rect 119291 238444 119292 238508
rect 119356 238444 119357 238508
rect 119291 238443 119357 238444
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 70899 180164 70965 180165
rect 70899 180100 70900 180164
rect 70964 180100 70965 180164
rect 70899 180099 70965 180100
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177716 97093 177717
rect 97027 177652 97028 177716
rect 97092 177652 97093 177716
rect 97027 177651 97093 177652
rect 98315 177716 98381 177717
rect 98315 177652 98316 177716
rect 98380 177652 98381 177716
rect 98315 177651 98381 177652
rect 97030 175130 97090 177651
rect 96960 175070 97090 175130
rect 98318 175130 98378 177651
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177716 100773 177717
rect 100707 177652 100708 177716
rect 100772 177652 100773 177716
rect 100707 177651 100773 177652
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177651
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 101998 175130 102058 176699
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 104571 177716 104637 177717
rect 104571 177652 104572 177716
rect 104636 177652 104637 177716
rect 104571 177651 104637 177652
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177651
rect 109539 177036 109605 177037
rect 109539 176972 109540 177036
rect 109604 176972 109605 177036
rect 109539 176971 109605 176972
rect 105675 176764 105741 176765
rect 105675 176700 105676 176764
rect 105740 176700 105741 176764
rect 105675 176699 105741 176700
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 105678 175130 105738 176699
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176699
rect 109542 175130 109602 176971
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113219 177716 113285 177717
rect 113219 177652 113220 177716
rect 113284 177652 113285 177716
rect 113219 177651 113285 177652
rect 110643 175404 110709 175405
rect 110643 175340 110644 175404
rect 110708 175340 110709 175404
rect 110643 175339 110709 175340
rect 112115 175404 112181 175405
rect 112115 175340 112116 175404
rect 112180 175340 112181 175404
rect 112115 175339 112181 175340
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 175339
rect 112118 175130 112178 175339
rect 113222 175130 113282 177651
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177716 114389 177717
rect 114323 177652 114324 177716
rect 114388 177652 114389 177716
rect 114323 177651 114389 177652
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177651
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 115798 175130 115858 176699
rect 117234 176600 117854 190338
rect 120954 230614 121574 238000
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177716 118437 177717
rect 118371 177652 118372 177716
rect 118436 177652 118437 177716
rect 118371 177651 118437 177652
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 116899 175540 116965 175541
rect 116899 175476 116900 175540
rect 116964 175476 116965 175540
rect 116899 175475 116965 175476
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175475
rect 118374 175130 118434 177651
rect 119478 175130 119538 177651
rect 120954 176600 121574 194058
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 177716 121933 177717
rect 121867 177652 121868 177716
rect 121932 177652 121933 177716
rect 121867 177651 121933 177652
rect 127019 177716 127085 177717
rect 127019 177652 127020 177716
rect 127084 177652 127085 177716
rect 127019 177651 127085 177652
rect 120763 175540 120829 175541
rect 120763 175476 120764 175540
rect 120828 175476 120829 175540
rect 120763 175475 120829 175476
rect 120766 175130 120826 175475
rect 121870 175130 121930 177651
rect 125731 177036 125797 177037
rect 125731 176972 125732 177036
rect 125796 176972 125797 177036
rect 125731 176971 125797 176972
rect 123155 176764 123221 176765
rect 123155 176700 123156 176764
rect 123220 176700 123221 176764
rect 123155 176699 123221 176700
rect 123158 175130 123218 176699
rect 124443 175540 124509 175541
rect 124443 175476 124444 175540
rect 124508 175476 124509 175540
rect 124443 175475 124509 175476
rect 124446 175130 124506 175475
rect 125734 175130 125794 176971
rect 127022 175130 127082 177651
rect 127794 176600 128414 200898
rect 131514 313174 132134 348618
rect 133094 329765 133154 445707
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 133827 393412 133893 393413
rect 133827 393348 133828 393412
rect 133892 393348 133893 393412
rect 133827 393347 133893 393348
rect 133091 329764 133157 329765
rect 133091 329700 133092 329764
rect 133156 329700 133157 329764
rect 133091 329699 133157 329700
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 133830 226269 133890 393347
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 133827 226268 133893 226269
rect 133827 226204 133828 226268
rect 133892 226204 133893 226268
rect 133827 226203 133893 226204
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 130702 175130 130762 176699
rect 131514 176600 132134 204618
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 133091 177036 133157 177037
rect 133091 176972 133092 177036
rect 133156 176972 133157 177036
rect 133091 176971 133157 176972
rect 132355 176764 132421 176765
rect 132355 176700 132356 176764
rect 132420 176700 132421 176764
rect 132355 176699 132421 176700
rect 132358 175130 132418 176699
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 176971
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 168419 398852 168485 398853
rect 168419 398788 168420 398852
rect 168484 398788 168485 398852
rect 168419 398787 168485 398788
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 179484 166277 179485
rect 166211 179420 166212 179484
rect 166276 179420 166277 179484
rect 166211 179419 166277 179420
rect 158851 175540 158917 175541
rect 158851 175476 158852 175540
rect 158916 175476 158917 175540
rect 158851 175475 158917 175476
rect 158854 175130 158914 175475
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 161669 166274 179419
rect 166395 175404 166461 175405
rect 166395 175340 166396 175404
rect 166460 175340 166461 175404
rect 166395 175339 166461 175340
rect 166398 162893 166458 175339
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166395 162892 166461 162893
rect 166395 162828 166396 162892
rect 166460 162828 166461 162892
rect 166395 162827 166461 162828
rect 166211 161668 166277 161669
rect 166211 161604 166212 161668
rect 166276 161604 166277 161668
rect 166211 161603 166277 161604
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166211 144940 166277 144941
rect 166211 144876 166212 144940
rect 166276 144876 166277 144940
rect 166211 144875 166277 144876
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 62987 69596 63053 69597
rect 62987 69532 62988 69596
rect 63052 69532 63053 69596
rect 62987 69531 63053 69532
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 85622 93533 85682 94830
rect 85619 93532 85685 93533
rect 85619 93468 85620 93532
rect 85684 93468 85685 93532
rect 85619 93467 85685 93468
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 86726 91221 86786 94830
rect 88014 92445 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88934 91221 88994 94830
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91221 93962 94830
rect 94920 94757 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 96008 94830 96354 94890
rect 94917 94756 94983 94757
rect 94917 94692 94918 94756
rect 94982 94692 94983 94756
rect 94917 94691 94983 94692
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91221 96722 94830
rect 97214 91221 97274 94830
rect 98134 92445 98194 94830
rect 98131 92444 98197 92445
rect 98131 92380 98132 92444
rect 98196 92380 98197 92444
rect 98131 92379 98197 92380
rect 98502 91357 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 92445 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 92444 100037 92445
rect 99971 92380 99972 92444
rect 100036 92380 100037 92444
rect 99971 92379 100037 92380
rect 100526 91221 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91765 101874 94830
rect 101811 91764 101877 91765
rect 101811 91700 101812 91764
rect 101876 91700 101877 91764
rect 101811 91699 101877 91700
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 91221 102794 93810
rect 103286 93261 103346 94830
rect 104304 94757 104364 95200
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 104301 94756 104367 94757
rect 104301 94692 104302 94756
rect 104366 94692 104367 94756
rect 104301 94691 104367 94692
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 92445 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106414 91221 106474 94830
rect 106782 92445 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 93533 107762 94830
rect 107699 93532 107765 93533
rect 107699 93468 107700 93532
rect 107764 93468 107765 93532
rect 107699 93467 107765 93468
rect 106779 92444 106845 92445
rect 106779 92380 106780 92444
rect 106844 92380 106845 92444
rect 106779 92379 106845 92380
rect 108070 91221 108130 94830
rect 109174 92309 109234 94830
rect 109171 92308 109237 92309
rect 109171 92244 109172 92308
rect 109236 92244 109237 92308
rect 109171 92243 109237 92244
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91221 111258 94830
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113038 94830 113204 94890
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 112302 91629 112362 94830
rect 113038 92445 113098 94830
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113035 92444 113101 92445
rect 113035 92380 113036 92444
rect 113100 92380 113101 92444
rect 113035 92379 113101 92380
rect 112299 91628 112365 91629
rect 112299 91564 112300 91628
rect 112364 91564 112365 91628
rect 112299 91563 112365 91564
rect 113222 91357 113282 93810
rect 113219 91356 113285 91357
rect 113219 91292 113220 91356
rect 113284 91292 113285 91356
rect 113219 91291 113285 91292
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 115430 91357 115490 94830
rect 115798 93533 115858 94830
rect 116680 94757 116740 95200
rect 117088 94890 117148 95200
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116677 94756 116743 94757
rect 116677 94692 116678 94756
rect 116742 94692 116743 94756
rect 116677 94691 116743 94692
rect 115795 93532 115861 93533
rect 115795 93468 115796 93532
rect 115860 93468 115861 93532
rect 115795 93467 115861 93468
rect 115427 91356 115493 91357
rect 115427 91292 115428 91356
rect 115492 91292 115493 91356
rect 115427 91291 115493 91292
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92173 118066 94830
rect 118003 92172 118069 92173
rect 118003 92108 118004 92172
rect 118068 92108 118069 92172
rect 118003 92107 118069 92108
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 119536 94830 119722 94890
rect 119294 91629 119354 94830
rect 119291 91628 119357 91629
rect 119291 91564 119292 91628
rect 119356 91564 119357 91628
rect 119291 91563 119357 91564
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120214 92445 120274 94830
rect 120624 94757 120684 95200
rect 121712 94890 121772 95200
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120621 94756 120687 94757
rect 120621 94692 120622 94756
rect 120686 94692 120687 94756
rect 120621 94691 120687 94692
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91221 121746 94830
rect 122054 93533 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122051 93532 122117 93533
rect 122051 93468 122052 93532
rect 122116 93468 122117 93532
rect 122051 93467 122117 93468
rect 122606 91490 122666 93810
rect 123158 92445 123218 94830
rect 124078 92445 124138 94830
rect 123155 92444 123221 92445
rect 123155 92380 123156 92444
rect 123220 92380 123221 92444
rect 123155 92379 123221 92380
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 124446 91221 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 92445 125426 94830
rect 125363 92444 125429 92445
rect 125363 92380 125364 92444
rect 125428 92380 125429 92444
rect 125363 92379 125429 92380
rect 125734 91765 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 91764 125797 91765
rect 125731 91700 125732 91764
rect 125796 91700 125797 91764
rect 125731 91699 125797 91700
rect 126470 91357 126530 94830
rect 126467 91356 126533 91357
rect 126467 91292 126468 91356
rect 126532 91292 126533 91356
rect 126467 91291 126533 91292
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 127574 91221 127634 94830
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133136 94757 133196 95200
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133133 94756 133199 94757
rect 133133 94692 133134 94756
rect 133198 94692 133199 94756
rect 133133 94691 133199 94692
rect 134382 92445 134442 94830
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 91629 136098 94830
rect 151496 94754 151556 95200
rect 151494 94694 151556 94754
rect 136035 91628 136101 91629
rect 136035 91564 136036 91628
rect 136100 91564 136101 91628
rect 136035 91563 136101 91564
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151494 92445 151554 94694
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151904 94754 151964 95200
rect 151904 94694 152106 94754
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 151678 91221 151738 94150
rect 152046 92445 152106 94694
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151675 91220 151741 91221
rect 151675 91156 151676 91220
rect 151740 91156 151741 91220
rect 151675 91155 151741 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 86597 166274 144875
rect 166395 135556 166461 135557
rect 166395 135492 166396 135556
rect 166460 135492 166461 135556
rect 166395 135491 166461 135492
rect 166211 86596 166277 86597
rect 166211 86532 166212 86596
rect 166276 86532 166277 86596
rect 166211 86531 166277 86532
rect 166398 84013 166458 135491
rect 167514 133174 168134 168618
rect 168422 168469 168482 398787
rect 171234 388894 171854 424338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 173019 393956 173085 393957
rect 173019 393892 173020 393956
rect 173084 393892 173085 393956
rect 173019 393891 173085 393892
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 168419 168468 168485 168469
rect 168419 168404 168420 168468
rect 168484 168404 168485 168468
rect 168419 168403 168485 168404
rect 171234 136894 171854 172338
rect 170259 136780 170325 136781
rect 170259 136716 170260 136780
rect 170324 136716 170325 136780
rect 170259 136715 170325 136716
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 168971 129844 169037 129845
rect 168971 129780 168972 129844
rect 169036 129780 169037 129844
rect 168971 129779 169037 129780
rect 168235 118012 168301 118013
rect 168235 117948 168236 118012
rect 168300 117948 168301 118012
rect 168235 117947 168301 117948
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 84012 166461 84013
rect 166395 83948 166396 84012
rect 166460 83948 166461 84012
rect 166395 83947 166461 83948
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 92309 168298 117947
rect 168235 92308 168301 92309
rect 168235 92244 168236 92308
rect 168300 92244 168301 92308
rect 168235 92243 168301 92244
rect 168974 78573 169034 129779
rect 169155 127260 169221 127261
rect 169155 127196 169156 127260
rect 169220 127196 169221 127260
rect 169155 127195 169221 127196
rect 169158 88229 169218 127195
rect 169155 88228 169221 88229
rect 169155 88164 169156 88228
rect 169220 88164 169221 88228
rect 169155 88163 169221 88164
rect 168971 78572 169037 78573
rect 168971 78508 168972 78572
rect 169036 78508 169037 78572
rect 168971 78507 169037 78508
rect 170262 77213 170322 136715
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170443 132836 170509 132837
rect 170443 132772 170444 132836
rect 170508 132772 170509 132836
rect 170443 132771 170509 132772
rect 170446 86733 170506 132771
rect 171234 100894 171854 136338
rect 173022 119373 173082 393891
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 173203 128484 173269 128485
rect 173203 128420 173204 128484
rect 173268 128420 173269 128484
rect 173203 128419 173269 128420
rect 173019 119372 173085 119373
rect 173019 119308 173020 119372
rect 173084 119308 173085 119372
rect 173019 119307 173085 119308
rect 172099 102236 172165 102237
rect 172099 102172 172100 102236
rect 172164 102172 172165 102236
rect 172099 102171 172165 102172
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 86732 170509 86733
rect 170443 86668 170444 86732
rect 170508 86668 170509 86732
rect 170443 86667 170509 86668
rect 170259 77212 170325 77213
rect 170259 77148 170260 77212
rect 170324 77148 170325 77212
rect 170259 77147 170325 77148
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 172102 91085 172162 102171
rect 172099 91084 172165 91085
rect 172099 91020 172100 91084
rect 172164 91020 172165 91084
rect 172099 91019 172165 91020
rect 173206 84149 173266 128419
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173203 84148 173269 84149
rect 173203 84084 173204 84148
rect 173268 84084 173269 84148
rect 173203 84083 173269 84084
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 227667 298212 227733 298213
rect 227667 298148 227668 298212
rect 227732 298148 227733 298212
rect 227667 298147 227733 298148
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 227670 174450 227730 298147
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 230427 227084 230493 227085
rect 230427 227020 230428 227084
rect 230492 227020 230493 227084
rect 230427 227019 230493 227020
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 228955 177444 229021 177445
rect 228955 177380 228956 177444
rect 229020 177380 229021 177444
rect 228955 177379 229021 177380
rect 228958 175130 229018 177379
rect 229507 175948 229573 175949
rect 229507 175884 229508 175948
rect 229572 175884 229573 175948
rect 229507 175883 229573 175884
rect 228958 175070 229202 175130
rect 229142 174997 229202 175070
rect 229139 174996 229205 174997
rect 229139 174932 229140 174996
rect 229204 174932 229205 174996
rect 229139 174931 229205 174932
rect 227670 174390 229202 174450
rect 229142 174317 229202 174390
rect 229139 174316 229205 174317
rect 229139 174252 229140 174316
rect 229204 174252 229205 174316
rect 229139 174251 229205 174252
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 229510 158133 229570 175883
rect 229507 158132 229573 158133
rect 229507 158068 229508 158132
rect 229572 158068 229573 158132
rect 229507 158067 229573 158068
rect 230430 147797 230490 227019
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 233187 197980 233253 197981
rect 233187 197916 233188 197980
rect 233252 197916 233253 197980
rect 233187 197915 233253 197916
rect 233190 148749 233250 197915
rect 234659 177580 234725 177581
rect 234659 177516 234660 177580
rect 234724 177516 234725 177580
rect 234659 177515 234725 177516
rect 233187 148748 233253 148749
rect 233187 148684 233188 148748
rect 233252 148684 233253 148748
rect 233187 148683 233253 148684
rect 230427 147796 230493 147797
rect 230427 147732 230428 147796
rect 230492 147732 230493 147796
rect 230427 147731 230493 147732
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 230979 146164 231045 146165
rect 230979 146100 230980 146164
rect 231044 146100 231045 146164
rect 230979 146099 231045 146100
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 230982 126037 231042 146099
rect 233739 143988 233805 143989
rect 233739 143924 233740 143988
rect 233804 143924 233805 143988
rect 233739 143923 233805 143924
rect 231347 141404 231413 141405
rect 231347 141340 231348 141404
rect 231412 141340 231413 141404
rect 231347 141339 231413 141340
rect 231350 133789 231410 141339
rect 232451 138412 232517 138413
rect 232451 138348 232452 138412
rect 232516 138348 232517 138412
rect 232451 138347 232517 138348
rect 231347 133788 231413 133789
rect 231347 133724 231348 133788
rect 231412 133724 231413 133788
rect 231347 133723 231413 133724
rect 231163 132972 231229 132973
rect 231163 132908 231164 132972
rect 231228 132908 231229 132972
rect 231163 132907 231229 132908
rect 230979 126036 231045 126037
rect 230979 125972 230980 126036
rect 231044 125972 231045 126036
rect 230979 125971 231045 125972
rect 230427 125356 230493 125357
rect 230427 125292 230428 125356
rect 230492 125292 230493 125356
rect 230427 125291 230493 125292
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 214419 105364 214485 105365
rect 214419 105300 214420 105364
rect 214484 105300 214485 105364
rect 214419 105299 214485 105300
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214422 93805 214482 105299
rect 230430 102373 230490 125291
rect 231166 123589 231226 132907
rect 231715 126308 231781 126309
rect 231715 126244 231716 126308
rect 231780 126244 231781 126308
rect 231715 126243 231781 126244
rect 231718 125493 231778 126243
rect 231715 125492 231781 125493
rect 231715 125428 231716 125492
rect 231780 125428 231781 125492
rect 231715 125427 231781 125428
rect 231163 123588 231229 123589
rect 231163 123524 231164 123588
rect 231228 123524 231229 123588
rect 231163 123523 231229 123524
rect 230427 102372 230493 102373
rect 230427 102308 230428 102372
rect 230492 102308 230493 102372
rect 230427 102307 230493 102308
rect 229323 98972 229389 98973
rect 229323 98970 229324 98972
rect 228958 98910 229324 98970
rect 228958 97066 229018 98910
rect 229323 98908 229324 98910
rect 229388 98908 229389 98972
rect 229323 98907 229389 98908
rect 228774 97006 229018 97066
rect 229139 97068 229205 97069
rect 227667 95436 227733 95437
rect 227667 95372 227668 95436
rect 227732 95372 227733 95436
rect 227667 95371 227733 95372
rect 214419 93804 214485 93805
rect 214419 93740 214420 93804
rect 214484 93740 214485 93804
rect 214419 93739 214485 93740
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 227670 24853 227730 95371
rect 228774 84210 228834 97006
rect 229139 97004 229140 97068
rect 229204 97004 229205 97068
rect 229139 97003 229205 97004
rect 229142 96930 229202 97003
rect 228958 96870 229202 96930
rect 228958 95437 229018 96870
rect 228955 95436 229021 95437
rect 228955 95372 228956 95436
rect 229020 95372 229021 95436
rect 228955 95371 229021 95372
rect 228222 84150 228834 84210
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 227667 24852 227733 24853
rect 227667 24788 227668 24852
rect 227732 24788 227733 24852
rect 227667 24787 227733 24788
rect 228222 19957 228282 84150
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228219 19956 228285 19957
rect 228219 19892 228220 19956
rect 228284 19892 228285 19956
rect 228219 19891 228285 19892
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 232454 11661 232514 138347
rect 233742 102237 233802 143923
rect 233923 142764 233989 142765
rect 233923 142700 233924 142764
rect 233988 142700 233989 142764
rect 233923 142699 233989 142700
rect 233926 106181 233986 142699
rect 234662 137869 234722 177515
rect 235794 165454 236414 200898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 242019 362268 242085 362269
rect 242019 362204 242020 362268
rect 242084 362204 242085 362268
rect 242019 362203 242085 362204
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 240363 315348 240429 315349
rect 240363 315284 240364 315348
rect 240428 315284 240429 315348
rect 240363 315283 240429 315284
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 236499 196756 236565 196757
rect 236499 196692 236500 196756
rect 236564 196692 236565 196756
rect 236499 196691 236565 196692
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 137868 234725 137869
rect 234659 137804 234660 137868
rect 234724 137804 234725 137868
rect 234659 137803 234725 137804
rect 235794 129454 236414 164898
rect 236502 138277 236562 196691
rect 237603 191044 237669 191045
rect 237603 190980 237604 191044
rect 237668 190980 237669 191044
rect 237603 190979 237669 190980
rect 237419 186964 237485 186965
rect 237419 186900 237420 186964
rect 237484 186900 237485 186964
rect 237419 186899 237485 186900
rect 237422 158813 237482 186899
rect 237606 167653 237666 190979
rect 238523 177308 238589 177309
rect 238523 177244 238524 177308
rect 238588 177244 238589 177308
rect 238523 177243 238589 177244
rect 238526 168330 238586 177243
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238707 168332 238773 168333
rect 238707 168330 238708 168332
rect 238526 168270 238708 168330
rect 238707 168268 238708 168270
rect 238772 168268 238773 168332
rect 238707 168267 238773 168268
rect 237603 167652 237669 167653
rect 237603 167588 237604 167652
rect 237668 167588 237669 167652
rect 237603 167587 237669 167588
rect 239075 167108 239141 167109
rect 239075 167044 239076 167108
rect 239140 167044 239141 167108
rect 239075 167043 239141 167044
rect 237971 159084 238037 159085
rect 237971 159020 237972 159084
rect 238036 159020 238037 159084
rect 237971 159019 238037 159020
rect 237419 158812 237485 158813
rect 237419 158748 237420 158812
rect 237484 158748 237485 158812
rect 237419 158747 237485 158748
rect 236499 138276 236565 138277
rect 236499 138212 236500 138276
rect 236564 138212 236565 138276
rect 236499 138211 236565 138212
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233923 106180 233989 106181
rect 233923 106116 233924 106180
rect 233988 106116 233989 106180
rect 233923 106115 233989 106116
rect 233739 102236 233805 102237
rect 233739 102172 233740 102236
rect 233804 102172 233805 102236
rect 233739 102171 233805 102172
rect 235794 93454 236414 128898
rect 237974 118421 238034 159019
rect 239078 135829 239138 167043
rect 239075 135828 239141 135829
rect 239075 135764 239076 135828
rect 239140 135764 239141 135828
rect 239075 135763 239141 135764
rect 239259 135828 239325 135829
rect 239259 135764 239260 135828
rect 239324 135764 239325 135828
rect 239259 135763 239325 135764
rect 237971 118420 238037 118421
rect 237971 118356 237972 118420
rect 238036 118356 238037 118420
rect 237971 118355 238037 118356
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 239262 64157 239322 135763
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239259 64156 239325 64157
rect 239259 64092 239260 64156
rect 239324 64092 239325 64156
rect 239259 64091 239325 64092
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 232451 11660 232517 11661
rect 232451 11596 232452 11660
rect 232516 11596 232517 11660
rect 232451 11595 232517 11596
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 240366 3501 240426 315283
rect 241651 280260 241717 280261
rect 241651 280196 241652 280260
rect 241716 280196 241717 280260
rect 241651 280195 241717 280196
rect 240547 245716 240613 245717
rect 240547 245652 240548 245716
rect 240612 245652 240613 245716
rect 240547 245651 240613 245652
rect 240550 153237 240610 245651
rect 240547 153236 240613 153237
rect 240547 153172 240548 153236
rect 240612 153172 240613 153236
rect 240547 153171 240613 153172
rect 240731 152420 240797 152421
rect 240731 152356 240732 152420
rect 240796 152356 240797 152420
rect 240731 152355 240797 152356
rect 240734 115565 240794 152355
rect 241654 141133 241714 280195
rect 241651 141132 241717 141133
rect 241651 141068 241652 141132
rect 241716 141068 241717 141132
rect 241651 141067 241717 141068
rect 240731 115564 240797 115565
rect 240731 115500 240732 115564
rect 240796 115500 240797 115564
rect 240731 115499 240797 115500
rect 242022 4861 242082 362203
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 251219 385660 251285 385661
rect 251219 385596 251220 385660
rect 251284 385596 251285 385660
rect 251219 385595 251285 385596
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 244227 331804 244293 331805
rect 244227 331740 244228 331804
rect 244292 331740 244293 331804
rect 244227 331739 244293 331740
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 289916 243005 289917
rect 242939 289852 242940 289916
rect 243004 289852 243005 289916
rect 242939 289851 243005 289852
rect 242942 143037 243002 289851
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242939 143036 243005 143037
rect 242939 142972 242940 143036
rect 243004 142972 243005 143036
rect 242939 142971 243005 142972
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 242019 4860 242085 4861
rect 242019 4796 242020 4860
rect 242084 4796 242085 4860
rect 242019 4795 242085 4796
rect 240363 3500 240429 3501
rect 240363 3436 240364 3500
rect 240428 3436 240429 3500
rect 240363 3435 240429 3436
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 244230 3501 244290 331739
rect 245699 322148 245765 322149
rect 245699 322084 245700 322148
rect 245764 322084 245765 322148
rect 245699 322083 245765 322084
rect 245702 3501 245762 322083
rect 246954 320614 247574 356058
rect 248459 334796 248525 334797
rect 248459 334732 248460 334796
rect 248524 334732 248525 334796
rect 248459 334731 248525 334732
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 247723 298348 247789 298349
rect 247723 298284 247724 298348
rect 247788 298284 247789 298348
rect 247723 298283 247789 298284
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 245883 182884 245949 182885
rect 245883 182820 245884 182884
rect 245948 182820 245949 182884
rect 245883 182819 245949 182820
rect 245886 141677 245946 182819
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 245883 141676 245949 141677
rect 245883 141612 245884 141676
rect 245948 141612 245949 141676
rect 245883 141611 245949 141612
rect 246954 140614 247574 176058
rect 247726 154869 247786 298283
rect 247723 154868 247789 154869
rect 247723 154804 247724 154868
rect 247788 154804 247789 154868
rect 247723 154803 247789 154804
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 244227 3500 244293 3501
rect 244227 3436 244228 3500
rect 244292 3436 244293 3500
rect 244227 3435 244293 3436
rect 245699 3500 245765 3501
rect 245699 3436 245700 3500
rect 245764 3436 245765 3500
rect 245699 3435 245765 3436
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 248462 3501 248522 334731
rect 249747 320788 249813 320789
rect 249747 320724 249748 320788
rect 249812 320724 249813 320788
rect 249747 320723 249813 320724
rect 249011 302836 249077 302837
rect 249011 302772 249012 302836
rect 249076 302772 249077 302836
rect 249011 302771 249077 302772
rect 248459 3500 248525 3501
rect 248459 3436 248460 3500
rect 248524 3436 248525 3500
rect 248459 3435 248525 3436
rect 249014 3365 249074 302771
rect 249750 3501 249810 320723
rect 250299 292772 250365 292773
rect 250299 292708 250300 292772
rect 250364 292708 250365 292772
rect 250299 292707 250365 292708
rect 250302 95437 250362 292707
rect 250299 95436 250365 95437
rect 250299 95372 250300 95436
rect 250364 95372 250365 95436
rect 250299 95371 250365 95372
rect 251222 3501 251282 385595
rect 252507 377364 252573 377365
rect 252507 377300 252508 377364
rect 252572 377300 252573 377364
rect 252507 377299 252573 377300
rect 252510 3501 252570 377299
rect 253794 363454 254414 398898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 255267 376004 255333 376005
rect 255267 375940 255268 376004
rect 255332 375940 255333 376004
rect 255267 375939 255333 375940
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 254531 114612 254597 114613
rect 254531 114548 254532 114612
rect 254596 114548 254597 114612
rect 254531 114547 254597 114548
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 254534 51781 254594 114547
rect 254531 51780 254597 51781
rect 254531 51716 254532 51780
rect 254596 51716 254597 51780
rect 254531 51715 254597 51716
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 249747 3500 249813 3501
rect 249747 3436 249748 3500
rect 249812 3436 249813 3500
rect 249747 3435 249813 3436
rect 251219 3500 251285 3501
rect 251219 3436 251220 3500
rect 251284 3436 251285 3500
rect 251219 3435 251285 3436
rect 252507 3500 252573 3501
rect 252507 3436 252508 3500
rect 252572 3436 252573 3500
rect 252507 3435 252573 3436
rect 253794 3454 254414 38898
rect 255270 3501 255330 375939
rect 257514 367174 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 259499 367708 259565 367709
rect 259499 367644 259500 367708
rect 259564 367644 259565 367708
rect 259499 367643 259565 367644
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257291 129028 257357 129029
rect 257291 128964 257292 129028
rect 257356 128964 257357 129028
rect 257291 128963 257357 128964
rect 255819 127124 255885 127125
rect 255819 127060 255820 127124
rect 255884 127060 255885 127124
rect 255819 127059 255885 127060
rect 255822 62797 255882 127059
rect 255819 62796 255885 62797
rect 255819 62732 255820 62796
rect 255884 62732 255885 62796
rect 255819 62731 255885 62732
rect 257294 40629 257354 128963
rect 257514 115174 258134 150618
rect 258763 131612 258829 131613
rect 258763 131548 258764 131612
rect 258828 131548 258829 131612
rect 258763 131547 258829 131548
rect 258579 130252 258645 130253
rect 258579 130188 258580 130252
rect 258644 130188 258645 130252
rect 258579 130187 258645 130188
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257291 40628 257357 40629
rect 257291 40564 257292 40628
rect 257356 40564 257357 40628
rect 257291 40563 257357 40564
rect 257514 7174 258134 42618
rect 258582 30973 258642 130187
rect 258766 73813 258826 131547
rect 258763 73812 258829 73813
rect 258763 73748 258764 73812
rect 258828 73748 258829 73812
rect 258763 73747 258829 73748
rect 258579 30972 258645 30973
rect 258579 30908 258580 30972
rect 258644 30908 258645 30972
rect 258579 30907 258645 30908
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 249011 3364 249077 3365
rect 249011 3300 249012 3364
rect 249076 3300 249077 3364
rect 249011 3299 249077 3300
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 255267 3500 255333 3501
rect 255267 3436 255268 3500
rect 255332 3436 255333 3500
rect 255267 3435 255333 3436
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 6618
rect 259502 3501 259562 367643
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 268331 307052 268397 307053
rect 268331 306988 268332 307052
rect 268396 306988 268397 307052
rect 268331 306987 268397 306988
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 262811 140180 262877 140181
rect 262811 140116 262812 140180
rect 262876 140116 262877 140180
rect 262811 140115 262877 140116
rect 262075 133244 262141 133245
rect 262075 133180 262076 133244
rect 262140 133180 262141 133244
rect 262075 133179 262141 133180
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 262078 24173 262138 133179
rect 262814 25533 262874 140115
rect 264099 132564 264165 132565
rect 264099 132500 264100 132564
rect 264164 132500 264165 132564
rect 264099 132499 264165 132500
rect 264102 72453 264162 132499
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 265755 98020 265821 98021
rect 265755 97956 265756 98020
rect 265820 97956 265821 98020
rect 265755 97955 265821 97956
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264099 72452 264165 72453
rect 264099 72388 264100 72452
rect 264164 72388 264165 72452
rect 264099 72387 264165 72388
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 262811 25532 262877 25533
rect 262811 25468 262812 25532
rect 262876 25468 262877 25532
rect 262811 25467 262877 25468
rect 262075 24172 262141 24173
rect 262075 24108 262076 24172
rect 262140 24108 262141 24172
rect 262075 24107 262141 24108
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 259499 3500 259565 3501
rect 259499 3436 259500 3500
rect 259564 3436 259565 3500
rect 259499 3435 259565 3436
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 265758 43485 265818 97955
rect 265755 43484 265821 43485
rect 265755 43420 265756 43484
rect 265820 43420 265821 43484
rect 265755 43419 265821 43420
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 268334 3365 268394 306987
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 278819 213212 278885 213213
rect 278819 213148 278820 213212
rect 278884 213148 278885 213212
rect 278819 213147 278885 213148
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 268515 175812 268581 175813
rect 268515 175748 268516 175812
rect 268580 175748 268581 175812
rect 268515 175747 268581 175748
rect 268518 174997 268578 175747
rect 268515 174996 268581 174997
rect 268515 174932 268516 174996
rect 268580 174932 268581 174996
rect 268515 174931 268581 174932
rect 278822 171150 278882 213147
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 178000 279854 208338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 288387 333300 288453 333301
rect 288387 333236 288388 333300
rect 288452 333236 288453 333300
rect 288387 333235 288453 333236
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 287099 293996 287165 293997
rect 287099 293932 287100 293996
rect 287164 293932 287165 293996
rect 287099 293931 287165 293932
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 285627 226948 285693 226949
rect 285627 226884 285628 226948
rect 285692 226884 285693 226948
rect 285627 226883 285693 226884
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 280291 192540 280357 192541
rect 280291 192476 280292 192540
rect 280356 192476 280357 192540
rect 280291 192475 280357 192476
rect 279371 177172 279437 177173
rect 279371 177108 279372 177172
rect 279436 177108 279437 177172
rect 279371 177107 279437 177108
rect 279374 175269 279434 177107
rect 279371 175268 279437 175269
rect 279371 175204 279372 175268
rect 279436 175204 279437 175268
rect 279371 175203 279437 175204
rect 278822 171090 279434 171150
rect 268515 167244 268581 167245
rect 268515 167180 268516 167244
rect 268580 167180 268581 167244
rect 268515 167179 268581 167180
rect 268518 166837 268578 167179
rect 268515 166836 268581 166837
rect 268515 166772 268516 166836
rect 268580 166772 268581 166836
rect 268515 166771 268581 166772
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 268515 163028 268581 163029
rect 268515 162964 268516 163028
rect 268580 162964 268581 163028
rect 268515 162963 268581 162964
rect 268518 159901 268578 162963
rect 268515 159900 268581 159901
rect 268515 159836 268516 159900
rect 268580 159836 268581 159900
rect 268515 159835 268581 159836
rect 279374 156773 279434 171090
rect 279371 156772 279437 156773
rect 279371 156708 279372 156772
rect 279436 156708 279437 156772
rect 279371 156707 279437 156708
rect 268515 147932 268581 147933
rect 268515 147868 268516 147932
rect 268580 147868 268581 147932
rect 268515 147867 268581 147868
rect 268518 146165 268578 147867
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 268515 146164 268581 146165
rect 268515 146100 268516 146164
rect 268580 146100 268581 146164
rect 268515 146099 268581 146100
rect 268515 140996 268581 140997
rect 268515 140932 268516 140996
rect 268580 140932 268581 140996
rect 268515 140931 268581 140932
rect 268518 140589 268578 140931
rect 268515 140588 268581 140589
rect 268515 140524 268516 140588
rect 268580 140524 268581 140588
rect 268515 140523 268581 140524
rect 280294 137053 280354 192475
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 281579 176220 281645 176221
rect 281579 176156 281580 176220
rect 281644 176156 281645 176220
rect 281579 176155 281645 176156
rect 281582 171733 281642 176155
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281579 171732 281645 171733
rect 281579 171668 281580 171732
rect 281644 171668 281645 171732
rect 281579 171667 281645 171668
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280291 137052 280357 137053
rect 280291 136988 280292 137052
rect 280356 136988 280357 137052
rect 280291 136987 280357 136988
rect 268515 134196 268581 134197
rect 268515 134132 268516 134196
rect 268580 134132 268581 134196
rect 268515 134131 268581 134132
rect 268518 133789 268578 134131
rect 268515 133788 268581 133789
rect 268515 133724 268516 133788
rect 268580 133724 268581 133788
rect 268515 133723 268581 133724
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 268515 128620 268581 128621
rect 268515 128556 268516 128620
rect 268580 128556 268581 128620
rect 268515 128555 268581 128556
rect 268518 128213 268578 128555
rect 268515 128212 268581 128213
rect 268515 128148 268516 128212
rect 268580 128148 268581 128212
rect 268515 128147 268581 128148
rect 268515 127260 268581 127261
rect 268515 127196 268516 127260
rect 268580 127196 268581 127260
rect 268515 127195 268581 127196
rect 268518 126853 268578 127195
rect 268515 126852 268581 126853
rect 268515 126788 268516 126852
rect 268580 126788 268581 126852
rect 268515 126787 268581 126788
rect 268515 123044 268581 123045
rect 268515 122980 268516 123044
rect 268580 122980 268581 123044
rect 268515 122979 268581 122980
rect 268518 122637 268578 122979
rect 268515 122636 268581 122637
rect 268515 122572 268516 122636
rect 268580 122572 268581 122636
rect 268515 122571 268581 122572
rect 268515 121684 268581 121685
rect 268515 121620 268516 121684
rect 268580 121620 268581 121684
rect 268515 121619 268581 121620
rect 268518 121277 268578 121619
rect 268515 121276 268581 121277
rect 268515 121212 268516 121276
rect 268580 121212 268581 121276
rect 268515 121211 268581 121212
rect 268515 117332 268581 117333
rect 268515 117268 268516 117332
rect 268580 117268 268581 117332
rect 268515 117267 268581 117268
rect 268518 116517 268578 117267
rect 268515 116516 268581 116517
rect 268515 116452 268516 116516
rect 268580 116452 268581 116516
rect 268515 116451 268581 116452
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 268515 107948 268581 107949
rect 268515 107884 268516 107948
rect 268580 107884 268581 107948
rect 268515 107883 268581 107884
rect 268518 107541 268578 107883
rect 268515 107540 268581 107541
rect 268515 107476 268516 107540
rect 268580 107476 268581 107540
rect 268515 107475 268581 107476
rect 282954 104614 283574 140058
rect 285630 106317 285690 226883
rect 285811 208996 285877 208997
rect 285811 208932 285812 208996
rect 285876 208932 285877 208996
rect 285811 208931 285877 208932
rect 285627 106316 285693 106317
rect 285627 106252 285628 106316
rect 285692 106252 285693 106316
rect 285627 106251 285693 106252
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 268515 102372 268581 102373
rect 268515 102308 268516 102372
rect 268580 102308 268581 102372
rect 268515 102307 268581 102308
rect 268518 100605 268578 102307
rect 268515 100604 268581 100605
rect 268515 100540 268516 100604
rect 268580 100540 268581 100604
rect 268515 100539 268581 100540
rect 281579 99380 281645 99381
rect 281579 99316 281580 99380
rect 281644 99316 281645 99380
rect 281579 99315 281645 99316
rect 268515 98020 268581 98021
rect 268515 97956 268516 98020
rect 268580 97956 268581 98020
rect 268515 97955 268581 97956
rect 279371 98020 279437 98021
rect 279371 97956 279372 98020
rect 279436 97956 279437 98020
rect 279371 97955 279437 97956
rect 268518 97205 268578 97955
rect 268515 97204 268581 97205
rect 268515 97140 268516 97204
rect 268580 97140 268581 97204
rect 268515 97139 268581 97140
rect 279374 95029 279434 97955
rect 279371 95028 279437 95029
rect 279371 94964 279372 95028
rect 279436 94964 279437 95028
rect 279371 94963 279437 94964
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 268331 3364 268397 3365
rect 268331 3300 268332 3364
rect 268396 3300 268397 3364
rect 268331 3299 268397 3300
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 281582 93533 281642 99315
rect 281579 93532 281645 93533
rect 281579 93468 281580 93532
rect 281644 93468 281645 93532
rect 281579 93467 281645 93468
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 285814 103189 285874 208931
rect 287102 106453 287162 293931
rect 287283 189684 287349 189685
rect 287283 189620 287284 189684
rect 287348 189620 287349 189684
rect 287283 189619 287349 189620
rect 287286 128757 287346 189619
rect 287283 128756 287349 128757
rect 287283 128692 287284 128756
rect 287348 128692 287349 128756
rect 287283 128691 287349 128692
rect 287099 106452 287165 106453
rect 287099 106388 287100 106452
rect 287164 106388 287165 106452
rect 287099 106387 287165 106388
rect 285811 103188 285877 103189
rect 285811 103124 285812 103188
rect 285876 103124 285877 103188
rect 285811 103123 285877 103124
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 288390 3501 288450 333235
rect 289794 327454 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 292619 336156 292685 336157
rect 292619 336092 292620 336156
rect 292684 336092 292685 336156
rect 292619 336091 292685 336092
rect 291147 334660 291213 334661
rect 291147 334596 291148 334660
rect 291212 334596 291213 334660
rect 291147 334595 291213 334596
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 288571 228308 288637 228309
rect 288571 228244 288572 228308
rect 288636 228244 288637 228308
rect 288571 228243 288637 228244
rect 288574 127125 288634 228243
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 290595 187100 290661 187101
rect 290595 187036 290596 187100
rect 290660 187036 290661 187100
rect 290595 187035 290661 187036
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288571 127124 288637 127125
rect 288571 127060 288572 127124
rect 288636 127060 288637 127124
rect 288571 127059 288637 127060
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 290598 109173 290658 187035
rect 290595 109172 290661 109173
rect 290595 109108 290596 109172
rect 290660 109108 290661 109172
rect 290595 109107 290661 109108
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288387 3500 288453 3501
rect 288387 3436 288388 3500
rect 288452 3436 288453 3500
rect 288387 3435 288453 3436
rect 289794 3454 290414 38898
rect 291150 3501 291210 334595
rect 291331 222868 291397 222869
rect 291331 222804 291332 222868
rect 291396 222804 291397 222868
rect 291331 222803 291397 222804
rect 291334 101013 291394 222803
rect 291331 101012 291397 101013
rect 291331 100948 291332 101012
rect 291396 100948 291397 101012
rect 291331 100947 291397 100948
rect 292622 3501 292682 336091
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 299611 369068 299677 369069
rect 299611 369004 299612 369068
rect 299676 369004 299677 369068
rect 299611 369003 299677 369004
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 295931 316708 295997 316709
rect 295931 316644 295932 316708
rect 295996 316644 295997 316708
rect 295931 316643 295997 316644
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 294275 178804 294341 178805
rect 294275 178740 294276 178804
rect 294340 178740 294341 178804
rect 294275 178739 294341 178740
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 294278 110533 294338 178739
rect 295379 178668 295445 178669
rect 295379 178604 295380 178668
rect 295444 178604 295445 178668
rect 295379 178603 295445 178604
rect 294275 110532 294341 110533
rect 294275 110468 294276 110532
rect 294340 110468 294341 110532
rect 294275 110467 294341 110468
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 291147 3500 291213 3501
rect 291147 3436 291148 3500
rect 291212 3436 291213 3500
rect 291147 3435 291213 3436
rect 292619 3500 292685 3501
rect 292619 3436 292620 3500
rect 292684 3436 292685 3500
rect 292619 3435 292685 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 6618
rect 295382 3501 295442 178603
rect 295934 3909 295994 316643
rect 297234 298894 297854 334338
rect 298691 329084 298757 329085
rect 298691 329020 298692 329084
rect 298756 329020 298757 329084
rect 298691 329019 298757 329020
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 295931 3908 295997 3909
rect 295931 3844 295932 3908
rect 295996 3844 295997 3908
rect 295931 3843 295997 3844
rect 295379 3500 295445 3501
rect 295379 3436 295380 3500
rect 295444 3436 295445 3500
rect 295379 3435 295445 3436
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 10338
rect 298694 3637 298754 329019
rect 298691 3636 298757 3637
rect 298691 3572 298692 3636
rect 298756 3572 298757 3636
rect 298691 3571 298757 3572
rect 299614 3501 299674 369003
rect 300954 338614 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 304947 370564 305013 370565
rect 304947 370500 304948 370564
rect 305012 370500 305013 370564
rect 304947 370499 305013 370500
rect 302739 363628 302805 363629
rect 302739 363564 302740 363628
rect 302804 363564 302805 363628
rect 302739 363563 302805 363564
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 3500 299677 3501
rect 299611 3436 299612 3500
rect 299676 3436 299677 3500
rect 299611 3435 299677 3436
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 302742 3909 302802 363563
rect 302739 3908 302805 3909
rect 302739 3844 302740 3908
rect 302804 3844 302805 3908
rect 302739 3843 302805 3844
rect 304950 3501 305010 370499
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 304947 3500 305013 3501
rect 304947 3436 304948 3500
rect 305012 3436 305013 3500
rect 304947 3435 305013 3436
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 76618 579218 76854 579454
rect 76618 578898 76854 579134
rect 87882 579218 88118 579454
rect 87882 578898 88118 579134
rect 99146 579218 99382 579454
rect 99146 578898 99382 579134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 82250 561218 82486 561454
rect 82250 560898 82486 561134
rect 93514 561218 93750 561454
rect 93514 560898 93750 561134
rect 76618 543218 76854 543454
rect 76618 542898 76854 543134
rect 87882 543218 88118 543454
rect 87882 542898 88118 543134
rect 99146 543218 99382 543454
rect 99146 542898 99382 543134
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 75618 471218 75854 471454
rect 75618 470898 75854 471134
rect 84882 471218 85118 471454
rect 84882 470898 85118 471134
rect 94146 471218 94382 471454
rect 94146 470898 94382 471134
rect 80250 453218 80486 453454
rect 80250 452898 80486 453134
rect 89514 453218 89750 453454
rect 89514 452898 89750 453134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76618 579454
rect 76854 579218 87882 579454
rect 88118 579218 99146 579454
rect 99382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76618 579134
rect 76854 578898 87882 579134
rect 88118 578898 99146 579134
rect 99382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 82250 561454
rect 82486 561218 93514 561454
rect 93750 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 82250 561134
rect 82486 560898 93514 561134
rect 93750 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76618 543454
rect 76854 543218 87882 543454
rect 88118 543218 99146 543454
rect 99382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76618 543134
rect 76854 542898 87882 543134
rect 88118 542898 99146 543134
rect 99382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 75618 471454
rect 75854 471218 84882 471454
rect 85118 471218 94146 471454
rect 94382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 75618 471134
rect 75854 470898 84882 471134
rect 85118 470898 94146 471134
rect 94382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 80250 453454
rect 80486 453218 89514 453454
rect 89750 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 80250 453134
rect 80486 452898 89514 453134
rect 89750 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 70000 0 1 440000
box -10 -52 30000 50000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 540000
box -10 -52 36000 42000
use wrapped_vga_clock  wrapped_vga_clock_1
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 46000 46000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 388000 74414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 492000 74414 538000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 584000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 388000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 388000 78134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 492000 78134 538000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 584000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 388000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 388000 81854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 492000 81854 538000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 584000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 388000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 388000 85574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 492000 85574 538000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 584000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 388000 99854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 492000 99854 538000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 584000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 388000 103574 538000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 584000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 388000 92414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 492000 92414 538000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 584000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 388000 96134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 492000 96134 538000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 584000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
