magic
tech sky130A
magscale 1 2
timestamp 1647706126
<< metal1 >>
rect 201494 703332 201500 703384
rect 201552 703372 201558 703384
rect 202782 703372 202788 703384
rect 201552 703344 202788 703372
rect 201552 703332 201558 703344
rect 202782 703332 202788 703344
rect 202840 703332 202846 703384
rect 77938 703264 77944 703316
rect 77996 703304 78002 703316
rect 267642 703304 267648 703316
rect 77996 703276 267648 703304
rect 77996 703264 78002 703276
rect 267642 703264 267648 703276
rect 267700 703264 267706 703316
rect 95142 703196 95148 703248
rect 95200 703236 95206 703248
rect 332502 703236 332508 703248
rect 95200 703208 332508 703236
rect 95200 703196 95206 703208
rect 332502 703196 332508 703208
rect 332560 703196 332566 703248
rect 109678 703128 109684 703180
rect 109736 703168 109742 703180
rect 348786 703168 348792 703180
rect 109736 703140 348792 703168
rect 109736 703128 109742 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 115198 703060 115204 703112
rect 115256 703100 115262 703112
rect 397454 703100 397460 703112
rect 115256 703072 397460 703100
rect 115256 703060 115262 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 76558 702992 76564 703044
rect 76616 703032 76622 703044
rect 358722 703032 358728 703044
rect 76616 703004 358728 703032
rect 76616 702992 76622 703004
rect 358722 702992 358728 703004
rect 358780 703032 358786 703044
rect 364978 703032 364984 703044
rect 358780 703004 364984 703032
rect 358780 702992 358786 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 104802 702924 104808 702976
rect 104860 702964 104866 702976
rect 413646 702964 413652 702976
rect 104860 702936 413652 702964
rect 104860 702924 104866 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 111702 702856 111708 702908
rect 111760 702896 111766 702908
rect 462314 702896 462320 702908
rect 111760 702868 462320 702896
rect 111760 702856 111766 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 75178 702788 75184 702840
rect 75236 702828 75242 702840
rect 429194 702828 429200 702840
rect 75236 702800 429200 702828
rect 75236 702788 75242 702800
rect 429194 702788 429200 702800
rect 429252 702828 429258 702840
rect 429838 702828 429844 702840
rect 429252 702800 429844 702828
rect 429252 702788 429258 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 117222 702720 117228 702772
rect 117280 702760 117286 702772
rect 478506 702760 478512 702772
rect 117280 702732 478512 702760
rect 117280 702720 117286 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 113082 702652 113088 702704
rect 113140 702692 113146 702704
rect 425698 702692 425704 702704
rect 113140 702664 425704 702692
rect 113140 702652 113146 702664
rect 425698 702652 425704 702664
rect 425756 702652 425762 702704
rect 492582 702652 492588 702704
rect 492640 702692 492646 702704
rect 494790 702692 494796 702704
rect 492640 702664 494796 702692
rect 492640 702652 492646 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 79318 702584 79324 702636
rect 79376 702624 79382 702636
rect 527174 702624 527180 702636
rect 79376 702596 527180 702624
rect 79376 702584 79382 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 108942 702516 108948 702568
rect 109000 702556 109006 702568
rect 521562 702556 521568 702568
rect 109000 702528 521568 702556
rect 109000 702516 109006 702528
rect 521562 702516 521568 702528
rect 521620 702516 521626 702568
rect 550542 702516 550548 702568
rect 550600 702556 550606 702568
rect 559650 702556 559656 702568
rect 550600 702528 559656 702556
rect 550600 702516 550606 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 68922 702448 68928 702500
rect 68980 702488 68986 702500
rect 543458 702488 543464 702500
rect 68980 702460 543464 702488
rect 68980 702448 68986 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 519538 700952 519544 701004
rect 519596 700992 519602 701004
rect 521562 700992 521568 701004
rect 519596 700964 521568 700992
rect 519596 700952 519602 700964
rect 521562 700952 521568 700964
rect 521620 700952 521626 701004
rect 137278 700408 137284 700460
rect 137336 700448 137342 700460
rect 137336 700420 142154 700448
rect 137336 700408 137342 700420
rect 69014 700340 69020 700392
rect 69072 700380 69078 700392
rect 137830 700380 137836 700392
rect 69072 700352 137836 700380
rect 69072 700340 69078 700352
rect 137830 700340 137836 700352
rect 137888 700340 137894 700392
rect 142126 700380 142154 700420
rect 154114 700380 154120 700392
rect 142126 700352 154120 700380
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 235166 700312 235172 700324
rect 62080 700284 235172 700312
rect 62080 700272 62086 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 238018 700272 238024 700324
rect 238076 700312 238082 700324
rect 283834 700312 283840 700324
rect 238076 700284 283840 700312
rect 238076 700272 238082 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 425698 700272 425704 700324
rect 425756 700312 425762 700324
rect 492582 700312 492588 700324
rect 425756 700284 492588 700312
rect 425756 700272 425762 700284
rect 492582 700272 492588 700284
rect 492640 700272 492646 700324
rect 521562 700272 521568 700324
rect 521620 700312 521626 700324
rect 550542 700312 550548 700324
rect 521620 700284 550548 700312
rect 521620 700272 521626 700284
rect 550542 700272 550548 700284
rect 550600 700272 550606 700324
rect 99282 698912 99288 698964
rect 99340 698952 99346 698964
rect 218974 698952 218980 698964
rect 99340 698924 218980 698952
rect 99340 698912 99346 698924
rect 218974 698912 218980 698924
rect 219032 698912 219038 698964
rect 24302 697620 24308 697672
rect 24360 697660 24366 697672
rect 106274 697660 106280 697672
rect 24360 697632 106280 697660
rect 24360 697620 24366 697632
rect 106274 697620 106280 697632
rect 106332 697620 106338 697672
rect 57882 697552 57888 697604
rect 57940 697592 57946 697604
rect 170306 697592 170312 697604
rect 57940 697564 170312 697592
rect 57940 697552 57946 697564
rect 170306 697552 170312 697564
rect 170364 697552 170370 697604
rect 334618 696940 334624 696992
rect 334676 696980 334682 696992
rect 580166 696980 580172 696992
rect 334676 696952 580172 696980
rect 334676 696940 334682 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 15838 683176 15844 683188
rect 3476 683148 15844 683176
rect 3476 683136 3482 683148
rect 15838 683136 15844 683148
rect 15896 683136 15902 683188
rect 320818 683136 320824 683188
rect 320876 683176 320882 683188
rect 580166 683176 580172 683188
rect 320876 683148 580172 683176
rect 320876 683136 320882 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 54478 670732 54484 670744
rect 3568 670704 54484 670732
rect 3568 670692 3574 670704
rect 54478 670692 54484 670704
rect 54536 670692 54542 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 87598 656928 87604 656940
rect 3476 656900 87604 656928
rect 3476 656888 3482 656900
rect 87598 656888 87604 656900
rect 87656 656888 87662 656940
rect 159358 643084 159364 643136
rect 159416 643124 159422 643136
rect 580166 643124 580172 643136
rect 159416 643096 580172 643124
rect 159416 643084 159422 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 276658 630640 276664 630692
rect 276716 630680 276722 630692
rect 579982 630680 579988 630692
rect 276716 630652 579988 630680
rect 276716 630640 276722 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 126238 616836 126244 616888
rect 126296 616876 126302 616888
rect 580166 616876 580172 616888
rect 126296 616848 580172 616876
rect 126296 616836 126302 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 35158 605860 35164 605872
rect 3568 605832 35164 605860
rect 3568 605820 3574 605832
rect 35158 605820 35164 605832
rect 35216 605820 35222 605872
rect 6914 598204 6920 598256
rect 6972 598244 6978 598256
rect 53098 598244 53104 598256
rect 6972 598216 53104 598244
rect 6972 598204 6978 598216
rect 53098 598204 53104 598216
rect 53156 598204 53162 598256
rect 53098 597524 53104 597576
rect 53156 597564 53162 597576
rect 85574 597564 85580 597576
rect 53156 597536 85580 597564
rect 53156 597524 53162 597536
rect 85574 597524 85580 597536
rect 85632 597524 85638 597576
rect 15838 596776 15844 596828
rect 15896 596816 15902 596828
rect 50982 596816 50988 596828
rect 15896 596788 50988 596816
rect 15896 596776 15902 596788
rect 50982 596776 50988 596788
rect 51040 596776 51046 596828
rect 50982 596164 50988 596216
rect 51040 596204 51046 596216
rect 71866 596204 71872 596216
rect 51040 596176 71872 596204
rect 51040 596164 51046 596176
rect 71866 596164 71872 596176
rect 71924 596164 71930 596216
rect 68830 594056 68836 594108
rect 68888 594096 68894 594108
rect 238018 594096 238024 594108
rect 68888 594068 238024 594096
rect 68888 594056 68894 594068
rect 238018 594056 238024 594068
rect 238076 594056 238082 594108
rect 81802 592628 81808 592680
rect 81860 592668 81866 592680
rect 580258 592668 580264 592680
rect 81860 592640 580264 592668
rect 81860 592628 81866 592640
rect 580258 592628 580264 592640
rect 580316 592628 580322 592680
rect 40034 592016 40040 592068
rect 40092 592056 40098 592068
rect 48222 592056 48228 592068
rect 40092 592028 48228 592056
rect 40092 592016 40098 592028
rect 48222 592016 48228 592028
rect 48280 592056 48286 592068
rect 74626 592056 74632 592068
rect 48280 592028 74632 592056
rect 48280 592016 48286 592028
rect 74626 592016 74632 592028
rect 74684 592016 74690 592068
rect 580258 592016 580264 592068
rect 580316 592056 580322 592068
rect 582374 592056 582380 592068
rect 580316 592028 582380 592056
rect 580316 592016 580322 592028
rect 582374 592016 582380 592028
rect 582432 592016 582438 592068
rect 385678 590656 385684 590708
rect 385736 590696 385742 590708
rect 579798 590696 579804 590708
rect 385736 590668 579804 590696
rect 385736 590656 385742 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3418 588548 3424 588600
rect 3476 588588 3482 588600
rect 57698 588588 57704 588600
rect 3476 588560 57704 588588
rect 3476 588548 3482 588560
rect 57698 588548 57704 588560
rect 57756 588548 57762 588600
rect 88334 588548 88340 588600
rect 88392 588588 88398 588600
rect 118878 588588 118884 588600
rect 88392 588560 118884 588588
rect 88392 588548 88398 588560
rect 118878 588548 118884 588560
rect 118936 588548 118942 588600
rect 57698 587868 57704 587920
rect 57756 587908 57762 587920
rect 95418 587908 95424 587920
rect 57756 587880 95424 587908
rect 57756 587868 57762 587880
rect 95418 587868 95424 587880
rect 95476 587868 95482 587920
rect 97902 586780 97908 586832
rect 97960 586820 97966 586832
rect 113358 586820 113364 586832
rect 97960 586792 113364 586820
rect 97960 586780 97966 586792
rect 113358 586780 113364 586792
rect 113416 586780 113422 586832
rect 52362 586712 52368 586764
rect 52420 586752 52426 586764
rect 85114 586752 85120 586764
rect 52420 586724 85120 586752
rect 52420 586712 52426 586724
rect 85114 586712 85120 586724
rect 85172 586712 85178 586764
rect 100570 586712 100576 586764
rect 100628 586752 100634 586764
rect 121638 586752 121644 586764
rect 100628 586724 121644 586752
rect 100628 586712 100634 586724
rect 121638 586712 121644 586724
rect 121696 586712 121702 586764
rect 49602 586644 49608 586696
rect 49660 586684 49666 586696
rect 81894 586684 81900 586696
rect 49660 586656 81900 586684
rect 49660 586644 49666 586656
rect 81894 586644 81900 586656
rect 81952 586644 81958 586696
rect 92842 586644 92848 586696
rect 92900 586684 92906 586696
rect 117314 586684 117320 586696
rect 92900 586656 117320 586684
rect 92900 586644 92906 586656
rect 117314 586644 117320 586656
rect 117372 586644 117378 586696
rect 48038 586576 48044 586628
rect 48096 586616 48102 586628
rect 84286 586616 84292 586628
rect 48096 586588 84292 586616
rect 48096 586576 48102 586588
rect 84286 586576 84292 586588
rect 84344 586576 84350 586628
rect 94866 586576 94872 586628
rect 94924 586616 94930 586628
rect 123110 586616 123116 586628
rect 94924 586588 123116 586616
rect 94924 586576 94930 586588
rect 123110 586576 123116 586588
rect 123168 586576 123174 586628
rect 42610 586508 42616 586560
rect 42668 586548 42674 586560
rect 80606 586548 80612 586560
rect 42668 586520 80612 586548
rect 42668 586508 42674 586520
rect 80606 586508 80612 586520
rect 80664 586508 80670 586560
rect 89622 586508 89628 586560
rect 89680 586548 89686 586560
rect 123018 586548 123024 586560
rect 89680 586520 123024 586548
rect 89680 586508 89686 586520
rect 123018 586508 123024 586520
rect 123076 586508 123082 586560
rect 68462 585760 68468 585812
rect 68520 585800 68526 585812
rect 137278 585800 137284 585812
rect 68520 585772 137284 585800
rect 68520 585760 68526 585772
rect 137278 585760 137284 585772
rect 137336 585760 137342 585812
rect 99282 585420 99288 585472
rect 99340 585460 99346 585472
rect 109034 585460 109040 585472
rect 99340 585432 109040 585460
rect 99340 585420 99346 585432
rect 109034 585420 109040 585432
rect 109092 585420 109098 585472
rect 87598 585352 87604 585404
rect 87656 585392 87662 585404
rect 110690 585392 110696 585404
rect 87656 585364 110696 585392
rect 87656 585352 87662 585364
rect 110690 585352 110696 585364
rect 110748 585352 110754 585404
rect 53650 585284 53656 585336
rect 53708 585324 53714 585336
rect 74902 585324 74908 585336
rect 53708 585296 74908 585324
rect 53708 585284 53714 585296
rect 74902 585284 74908 585296
rect 74960 585284 74966 585336
rect 94130 585284 94136 585336
rect 94188 585324 94194 585336
rect 94188 585296 99512 585324
rect 94188 585284 94194 585296
rect 46750 585216 46756 585268
rect 46808 585256 46814 585268
rect 83182 585256 83188 585268
rect 46808 585228 83188 585256
rect 46808 585216 46814 585228
rect 83182 585216 83188 585228
rect 83240 585216 83246 585268
rect 41230 585148 41236 585200
rect 41288 585188 41294 585200
rect 78030 585188 78036 585200
rect 41288 585160 78036 585188
rect 41288 585148 41294 585160
rect 78030 585148 78036 585160
rect 78088 585148 78094 585200
rect 98730 585148 98736 585200
rect 98788 585188 98794 585200
rect 99282 585188 99288 585200
rect 98788 585160 99288 585188
rect 98788 585148 98794 585160
rect 99282 585148 99288 585160
rect 99340 585148 99346 585200
rect 99484 585188 99512 585296
rect 118786 585188 118792 585200
rect 99484 585160 118792 585188
rect 118786 585148 118792 585160
rect 118844 585148 118850 585200
rect 103146 584400 103152 584452
rect 103204 584440 103210 584452
rect 104802 584440 104808 584452
rect 103204 584412 104808 584440
rect 103204 584400 103210 584412
rect 104802 584400 104808 584412
rect 104860 584440 104866 584452
rect 112070 584440 112076 584452
rect 104860 584412 112076 584440
rect 104860 584400 104866 584412
rect 112070 584400 112076 584412
rect 112128 584400 112134 584452
rect 55122 584060 55128 584112
rect 55180 584100 55186 584112
rect 73338 584100 73344 584112
rect 55180 584072 73344 584100
rect 55180 584060 55186 584072
rect 73338 584060 73344 584072
rect 73396 584060 73402 584112
rect 45462 583992 45468 584044
rect 45520 584032 45526 584044
rect 78674 584032 78680 584044
rect 45520 584004 78680 584032
rect 45520 583992 45526 584004
rect 78674 583992 78680 584004
rect 78732 583992 78738 584044
rect 88978 583992 88984 584044
rect 89036 584032 89042 584044
rect 111978 584032 111984 584044
rect 89036 584004 111984 584032
rect 89036 583992 89042 584004
rect 111978 583992 111984 584004
rect 112036 583992 112042 584044
rect 59170 583924 59176 583976
rect 59228 583964 59234 583976
rect 76558 583964 76564 583976
rect 59228 583936 76564 583964
rect 59228 583924 59234 583936
rect 76558 583924 76564 583936
rect 76616 583924 76622 583976
rect 77846 583924 77852 583976
rect 77904 583964 77910 583976
rect 79318 583964 79324 583976
rect 77904 583936 79324 583964
rect 77904 583924 77910 583936
rect 79318 583924 79324 583936
rect 79376 583924 79382 583976
rect 101306 583924 101312 583976
rect 101364 583964 101370 583976
rect 113266 583964 113272 583976
rect 101364 583936 113272 583964
rect 101364 583924 101370 583936
rect 113266 583924 113272 583936
rect 113324 583924 113330 583976
rect 70302 583856 70308 583908
rect 70360 583896 70366 583908
rect 82998 583896 83004 583908
rect 70360 583868 83004 583896
rect 70360 583856 70366 583868
rect 82998 583856 83004 583868
rect 83056 583856 83062 583908
rect 103882 583856 103888 583908
rect 103940 583896 103946 583908
rect 120166 583896 120172 583908
rect 103940 583868 120172 583896
rect 103940 583856 103946 583868
rect 120166 583856 120172 583868
rect 120224 583856 120230 583908
rect 47946 583788 47952 583840
rect 48004 583828 48010 583840
rect 77846 583828 77852 583840
rect 48004 583800 77852 583828
rect 48004 583788 48010 583800
rect 77846 583788 77852 583800
rect 77904 583788 77910 583840
rect 96522 583788 96528 583840
rect 96580 583828 96586 583840
rect 118694 583828 118700 583840
rect 96580 583800 118700 583828
rect 96580 583788 96586 583800
rect 118694 583788 118700 583800
rect 118752 583788 118758 583840
rect 65886 583720 65892 583772
rect 65944 583760 65950 583772
rect 70946 583760 70952 583772
rect 65944 583732 70952 583760
rect 65944 583720 65950 583732
rect 70946 583720 70952 583732
rect 71004 583720 71010 583772
rect 105538 583720 105544 583772
rect 105596 583760 105602 583772
rect 114554 583760 114560 583772
rect 105596 583732 114560 583760
rect 105596 583720 105602 583732
rect 114554 583720 114560 583732
rect 114612 583720 114618 583772
rect 56410 582972 56416 583024
rect 56468 583012 56474 583024
rect 71774 583012 71780 583024
rect 56468 582984 71780 583012
rect 56468 582972 56474 582984
rect 71774 582972 71780 582984
rect 71832 582972 71838 583024
rect 92290 582632 92296 582684
rect 92348 582672 92354 582684
rect 110506 582672 110512 582684
rect 92348 582644 110512 582672
rect 92348 582632 92354 582644
rect 110506 582632 110512 582644
rect 110564 582632 110570 582684
rect 70210 582564 70216 582616
rect 70268 582604 70274 582616
rect 84470 582604 84476 582616
rect 70268 582576 84476 582604
rect 70268 582564 70274 582576
rect 84470 582564 84476 582576
rect 84528 582564 84534 582616
rect 97442 582564 97448 582616
rect 97500 582604 97506 582616
rect 116026 582604 116032 582616
rect 97500 582576 116032 582604
rect 97500 582564 97506 582576
rect 116026 582564 116032 582576
rect 116084 582564 116090 582616
rect 50798 582496 50804 582548
rect 50856 582536 50862 582548
rect 76742 582536 76748 582548
rect 50856 582508 76748 582536
rect 50856 582496 50862 582508
rect 76742 582496 76748 582508
rect 76800 582496 76806 582548
rect 99282 582496 99288 582548
rect 99340 582536 99346 582548
rect 120074 582536 120080 582548
rect 99340 582508 120080 582536
rect 99340 582496 99346 582508
rect 120074 582496 120080 582508
rect 120132 582496 120138 582548
rect 3418 582428 3424 582480
rect 3476 582468 3482 582480
rect 107654 582468 107660 582480
rect 3476 582440 107660 582468
rect 3476 582428 3482 582440
rect 107654 582428 107660 582440
rect 107712 582428 107718 582480
rect 69106 582360 69112 582412
rect 69164 582400 69170 582412
rect 580166 582400 580172 582412
rect 69164 582372 580172 582400
rect 69164 582360 69170 582372
rect 580166 582360 580172 582372
rect 580224 582360 580230 582412
rect 65518 581680 65524 581732
rect 65576 581720 65582 581732
rect 75454 581720 75460 581732
rect 65576 581692 75460 581720
rect 65576 581680 65582 581692
rect 75454 581680 75460 581692
rect 75512 581680 75518 581732
rect 79318 581680 79324 581732
rect 79376 581680 79382 581732
rect 90266 581680 90272 581732
rect 90324 581720 90330 581732
rect 90324 581692 93854 581720
rect 90324 581680 90330 581692
rect 39758 581204 39764 581256
rect 39816 581244 39822 581256
rect 67634 581244 67640 581256
rect 39816 581216 67640 581244
rect 39816 581204 39822 581216
rect 67634 581204 67640 581216
rect 67692 581204 67698 581256
rect 59078 581136 59084 581188
rect 59136 581176 59142 581188
rect 79336 581176 79364 581680
rect 59136 581148 79364 581176
rect 59136 581136 59142 581148
rect 43806 581068 43812 581120
rect 43864 581108 43870 581120
rect 65518 581108 65524 581120
rect 43864 581080 65524 581108
rect 43864 581068 43870 581080
rect 65518 581068 65524 581080
rect 65576 581068 65582 581120
rect 36998 581000 37004 581052
rect 37056 581040 37062 581052
rect 70394 581040 70400 581052
rect 37056 581012 70400 581040
rect 37056 581000 37062 581012
rect 70394 581000 70400 581012
rect 70452 581000 70458 581052
rect 93826 581040 93854 581692
rect 104434 581680 104440 581732
rect 104492 581680 104498 581732
rect 104986 581680 104992 581732
rect 105044 581720 105050 581732
rect 105044 581692 113174 581720
rect 105044 581680 105050 581692
rect 104452 581108 104480 581680
rect 113146 581176 113174 581692
rect 114646 581176 114652 581188
rect 113146 581148 114652 581176
rect 114646 581136 114652 581148
rect 114704 581136 114710 581188
rect 126974 581108 126980 581120
rect 104452 581080 126980 581108
rect 126974 581068 126980 581080
rect 127032 581068 127038 581120
rect 121454 581040 121460 581052
rect 93826 581012 121460 581040
rect 121454 581000 121460 581012
rect 121512 581000 121518 581052
rect 108942 579708 108948 579760
rect 109000 579748 109006 579760
rect 128354 579748 128360 579760
rect 109000 579720 128360 579748
rect 109000 579708 109006 579720
rect 128354 579708 128360 579720
rect 128412 579708 128418 579760
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 15838 579680 15844 579692
rect 3384 579652 15844 579680
rect 3384 579640 3390 579652
rect 15838 579640 15844 579652
rect 15896 579640 15902 579692
rect 52178 579640 52184 579692
rect 52236 579680 52242 579692
rect 69014 579680 69020 579692
rect 52236 579652 69020 579680
rect 52236 579640 52242 579652
rect 69014 579640 69020 579652
rect 69072 579640 69078 579692
rect 57238 578212 57244 578264
rect 57296 578252 57302 578264
rect 67634 578252 67640 578264
rect 57296 578224 67640 578252
rect 57296 578212 57302 578224
rect 67634 578212 67640 578224
rect 67692 578212 67698 578264
rect 108942 578212 108948 578264
rect 109000 578252 109006 578264
rect 134150 578252 134156 578264
rect 109000 578224 134156 578252
rect 109000 578212 109006 578224
rect 134150 578212 134156 578224
rect 134208 578212 134214 578264
rect 356698 577464 356704 577516
rect 356756 577504 356762 577516
rect 429194 577504 429200 577516
rect 356756 577476 429200 577504
rect 356756 577464 356762 577476
rect 429194 577464 429200 577476
rect 429252 577464 429258 577516
rect 108942 576852 108948 576904
rect 109000 576892 109006 576904
rect 129826 576892 129832 576904
rect 109000 576864 129832 576892
rect 109000 576852 109006 576864
rect 129826 576852 129832 576864
rect 129884 576852 129890 576904
rect 108758 575560 108764 575612
rect 108816 575600 108822 575612
rect 131114 575600 131120 575612
rect 108816 575572 131120 575600
rect 108816 575560 108822 575572
rect 131114 575560 131120 575572
rect 131172 575560 131178 575612
rect 34422 575492 34428 575544
rect 34480 575532 34486 575544
rect 67634 575532 67640 575544
rect 34480 575504 67640 575532
rect 34480 575492 34486 575504
rect 67634 575492 67640 575504
rect 67692 575492 67698 575544
rect 108942 575492 108948 575544
rect 109000 575532 109006 575544
rect 122742 575532 122748 575544
rect 109000 575504 122748 575532
rect 109000 575492 109006 575504
rect 122742 575492 122748 575504
rect 122800 575532 122806 575544
rect 429838 575532 429844 575544
rect 122800 575504 429844 575532
rect 122800 575492 122806 575504
rect 429838 575492 429844 575504
rect 429896 575492 429902 575544
rect 59262 574064 59268 574116
rect 59320 574104 59326 574116
rect 67634 574104 67640 574116
rect 59320 574076 67640 574104
rect 59320 574064 59326 574076
rect 67634 574064 67640 574076
rect 67692 574064 67698 574116
rect 108942 574064 108948 574116
rect 109000 574104 109006 574116
rect 124214 574104 124220 574116
rect 109000 574076 124220 574104
rect 109000 574064 109006 574076
rect 124214 574064 124220 574076
rect 124272 574064 124278 574116
rect 65978 573316 65984 573368
rect 66036 573356 66042 573368
rect 68094 573356 68100 573368
rect 66036 573328 68100 573356
rect 66036 573316 66042 573328
rect 68094 573316 68100 573328
rect 68152 573316 68158 573368
rect 108666 573316 108672 573368
rect 108724 573356 108730 573368
rect 130378 573356 130384 573368
rect 108724 573328 130384 573356
rect 108724 573316 108730 573328
rect 130378 573316 130384 573328
rect 130436 573316 130442 573368
rect 61838 572704 61844 572756
rect 61896 572744 61902 572756
rect 67634 572744 67640 572756
rect 61896 572716 67640 572744
rect 61896 572704 61902 572716
rect 67634 572704 67640 572716
rect 67692 572704 67698 572756
rect 64690 571956 64696 572008
rect 64748 571996 64754 572008
rect 67818 571996 67824 572008
rect 64748 571968 67824 571996
rect 64748 571956 64754 571968
rect 67818 571956 67824 571968
rect 67876 571956 67882 572008
rect 105630 571956 105636 572008
rect 105688 571996 105694 572008
rect 110598 571996 110604 572008
rect 105688 571968 110604 571996
rect 105688 571956 105694 571968
rect 110598 571956 110604 571968
rect 110656 571956 110662 572008
rect 108942 571344 108948 571396
rect 109000 571384 109006 571396
rect 133874 571384 133880 571396
rect 109000 571356 133880 571384
rect 109000 571344 109006 571356
rect 133874 571344 133880 571356
rect 133932 571344 133938 571396
rect 108942 569984 108948 570036
rect 109000 570024 109006 570036
rect 120258 570024 120264 570036
rect 109000 569996 120264 570024
rect 109000 569984 109006 569996
rect 120258 569984 120264 569996
rect 120316 569984 120322 570036
rect 41322 569916 41328 569968
rect 41380 569956 41386 569968
rect 67634 569956 67640 569968
rect 41380 569928 67640 569956
rect 41380 569916 41386 569928
rect 67634 569916 67640 569928
rect 67692 569916 67698 569968
rect 108850 569916 108856 569968
rect 108908 569956 108914 569968
rect 142154 569956 142160 569968
rect 108908 569928 142160 569956
rect 108908 569916 108914 569928
rect 142154 569916 142160 569928
rect 142212 569916 142218 569968
rect 64598 568624 64604 568676
rect 64656 568664 64662 568676
rect 67726 568664 67732 568676
rect 64656 568636 67732 568664
rect 64656 568624 64662 568636
rect 67726 568624 67732 568636
rect 67784 568624 67790 568676
rect 61746 568556 61752 568608
rect 61804 568596 61810 568608
rect 67634 568596 67640 568608
rect 61804 568568 67640 568596
rect 61804 568556 61810 568568
rect 67634 568556 67640 568568
rect 67692 568556 67698 568608
rect 108942 568556 108948 568608
rect 109000 568596 109006 568608
rect 128998 568596 129004 568608
rect 109000 568568 129004 568596
rect 109000 568556 109006 568568
rect 128998 568556 129004 568568
rect 129056 568556 129062 568608
rect 106918 567808 106924 567860
rect 106976 567848 106982 567860
rect 117406 567848 117412 567860
rect 106976 567820 117412 567848
rect 106976 567808 106982 567820
rect 117406 567808 117412 567820
rect 117464 567808 117470 567860
rect 66070 567264 66076 567316
rect 66128 567304 66134 567316
rect 67726 567304 67732 567316
rect 66128 567276 67732 567304
rect 66128 567264 66134 567276
rect 67726 567264 67732 567276
rect 67784 567264 67790 567316
rect 108942 567264 108948 567316
rect 109000 567304 109006 567316
rect 117958 567304 117964 567316
rect 109000 567276 117964 567304
rect 109000 567264 109006 567276
rect 117958 567264 117964 567276
rect 118016 567264 118022 567316
rect 63218 567196 63224 567248
rect 63276 567236 63282 567248
rect 67634 567236 67640 567248
rect 63276 567208 67640 567236
rect 63276 567196 63282 567208
rect 67634 567196 67640 567208
rect 67692 567196 67698 567248
rect 108850 567196 108856 567248
rect 108908 567236 108914 567248
rect 125870 567236 125876 567248
rect 108908 567208 125876 567236
rect 108908 567196 108914 567208
rect 125870 567196 125876 567208
rect 125928 567196 125934 567248
rect 108942 565904 108948 565956
rect 109000 565944 109006 565956
rect 113174 565944 113180 565956
rect 109000 565916 113180 565944
rect 109000 565904 109006 565916
rect 113174 565904 113180 565916
rect 113232 565904 113238 565956
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 25498 565876 25504 565888
rect 3292 565848 25504 565876
rect 3292 565836 3298 565848
rect 25498 565836 25504 565848
rect 25556 565836 25562 565888
rect 64782 565836 64788 565888
rect 64840 565876 64846 565888
rect 67634 565876 67640 565888
rect 64840 565848 67640 565876
rect 64840 565836 64846 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 108390 565836 108396 565888
rect 108448 565876 108454 565888
rect 111886 565876 111892 565888
rect 108448 565848 111892 565876
rect 108448 565836 108454 565848
rect 111886 565836 111892 565848
rect 111944 565836 111950 565888
rect 429838 565088 429844 565140
rect 429896 565128 429902 565140
rect 497458 565128 497464 565140
rect 429896 565100 497464 565128
rect 429896 565088 429902 565100
rect 497458 565088 497464 565100
rect 497516 565128 497522 565140
rect 504358 565128 504364 565140
rect 497516 565100 504364 565128
rect 497516 565088 497522 565100
rect 504358 565088 504364 565100
rect 504416 565088 504422 565140
rect 41138 564476 41144 564528
rect 41196 564516 41202 564528
rect 67634 564516 67640 564528
rect 41196 564488 67640 564516
rect 41196 564476 41202 564488
rect 67634 564476 67640 564488
rect 67692 564476 67698 564528
rect 108942 564476 108948 564528
rect 109000 564516 109006 564528
rect 123202 564516 123208 564528
rect 109000 564488 123208 564516
rect 109000 564476 109006 564488
rect 123202 564476 123208 564488
rect 123260 564476 123266 564528
rect 108850 564408 108856 564460
rect 108908 564448 108914 564460
rect 133138 564448 133144 564460
rect 108908 564420 133144 564448
rect 108908 564408 108914 564420
rect 133138 564408 133144 564420
rect 133196 564448 133202 564460
rect 155218 564448 155224 564460
rect 133196 564420 155224 564448
rect 133196 564408 133202 564420
rect 155218 564408 155224 564420
rect 155276 564408 155282 564460
rect 108942 564340 108948 564392
rect 109000 564380 109006 564392
rect 117222 564380 117228 564392
rect 109000 564352 117228 564380
rect 109000 564340 109006 564352
rect 117222 564340 117228 564352
rect 117280 564340 117286 564392
rect 117222 563660 117228 563712
rect 117280 563700 117286 563712
rect 138014 563700 138020 563712
rect 117280 563672 138020 563700
rect 117280 563660 117286 563672
rect 138014 563660 138020 563672
rect 138072 563660 138078 563712
rect 504358 563660 504364 563712
rect 504416 563700 504422 563712
rect 580166 563700 580172 563712
rect 504416 563672 580172 563700
rect 504416 563660 504422 563672
rect 580166 563660 580172 563672
rect 580224 563660 580230 563712
rect 49418 563048 49424 563100
rect 49476 563088 49482 563100
rect 67634 563088 67640 563100
rect 49476 563060 67640 563088
rect 49476 563048 49482 563060
rect 67634 563048 67640 563060
rect 67692 563048 67698 563100
rect 61102 562300 61108 562352
rect 61160 562340 61166 562352
rect 62022 562340 62028 562352
rect 61160 562312 62028 562340
rect 61160 562300 61166 562312
rect 62022 562300 62028 562312
rect 62080 562340 62086 562352
rect 67634 562340 67640 562352
rect 62080 562312 67640 562340
rect 62080 562300 62086 562312
rect 67634 562300 67640 562312
rect 67692 562300 67698 562352
rect 60366 561688 60372 561740
rect 60424 561728 60430 561740
rect 67634 561728 67640 561740
rect 60424 561700 67640 561728
rect 60424 561688 60430 561700
rect 67634 561688 67640 561700
rect 67692 561688 67698 561740
rect 56502 561620 56508 561672
rect 56560 561660 56566 561672
rect 61102 561660 61108 561672
rect 56560 561632 61108 561660
rect 56560 561620 56566 561632
rect 61102 561620 61108 561632
rect 61160 561620 61166 561672
rect 60458 560328 60464 560380
rect 60516 560368 60522 560380
rect 67726 560368 67732 560380
rect 60516 560340 67732 560368
rect 60516 560328 60522 560340
rect 67726 560328 67732 560340
rect 67784 560328 67790 560380
rect 108942 560328 108948 560380
rect 109000 560368 109006 560380
rect 116118 560368 116124 560380
rect 109000 560340 116124 560368
rect 109000 560328 109006 560340
rect 116118 560328 116124 560340
rect 116176 560328 116182 560380
rect 57790 560260 57796 560312
rect 57848 560300 57854 560312
rect 67634 560300 67640 560312
rect 57848 560272 67640 560300
rect 57848 560260 57854 560272
rect 67634 560260 67640 560272
rect 67692 560260 67698 560312
rect 108206 560260 108212 560312
rect 108264 560300 108270 560312
rect 140774 560300 140780 560312
rect 108264 560272 140780 560300
rect 108264 560260 108270 560272
rect 140774 560260 140780 560272
rect 140832 560260 140838 560312
rect 136634 559512 136640 559564
rect 136692 559552 136698 559564
rect 201494 559552 201500 559564
rect 136692 559524 201500 559552
rect 136692 559512 136698 559524
rect 201494 559512 201500 559524
rect 201552 559512 201558 559564
rect 108942 558968 108948 559020
rect 109000 559008 109006 559020
rect 135438 559008 135444 559020
rect 109000 558980 135444 559008
rect 109000 558968 109006 558980
rect 135438 558968 135444 558980
rect 135496 558968 135502 559020
rect 42702 558900 42708 558952
rect 42760 558940 42766 558952
rect 67634 558940 67640 558952
rect 42760 558912 67640 558940
rect 42760 558900 42766 558912
rect 67634 558900 67640 558912
rect 67692 558900 67698 558952
rect 108850 558900 108856 558952
rect 108908 558940 108914 558952
rect 136634 558940 136640 558952
rect 108908 558912 136640 558940
rect 108908 558900 108914 558912
rect 136634 558900 136640 558912
rect 136692 558900 136698 558952
rect 66162 558288 66168 558340
rect 66220 558328 66226 558340
rect 68830 558328 68836 558340
rect 66220 558300 68836 558328
rect 66220 558288 66226 558300
rect 68830 558288 68836 558300
rect 68888 558288 68894 558340
rect 56318 557540 56324 557592
rect 56376 557580 56382 557592
rect 67634 557580 67640 557592
rect 56376 557552 67640 557580
rect 56376 557540 56382 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 108942 557540 108948 557592
rect 109000 557580 109006 557592
rect 115934 557580 115940 557592
rect 109000 557552 115940 557580
rect 109000 557540 109006 557552
rect 115934 557540 115940 557552
rect 115992 557540 115998 557592
rect 108942 556520 108948 556572
rect 109000 556560 109006 556572
rect 113910 556560 113916 556572
rect 109000 556532 113916 556560
rect 109000 556520 109006 556532
rect 113910 556520 113916 556532
rect 113968 556520 113974 556572
rect 43714 556248 43720 556300
rect 43772 556288 43778 556300
rect 67634 556288 67640 556300
rect 43772 556260 67640 556288
rect 43772 556248 43778 556260
rect 67634 556248 67640 556260
rect 67692 556248 67698 556300
rect 37090 556180 37096 556232
rect 37148 556220 37154 556232
rect 67818 556220 67824 556232
rect 37148 556192 67824 556220
rect 37148 556180 37154 556192
rect 67818 556180 67824 556192
rect 67876 556180 67882 556232
rect 55030 556112 55036 556164
rect 55088 556152 55094 556164
rect 57882 556152 57888 556164
rect 55088 556124 57888 556152
rect 55088 556112 55094 556124
rect 57882 556112 57888 556124
rect 57940 556152 57946 556164
rect 67726 556152 67732 556164
rect 57940 556124 67732 556152
rect 57940 556112 57946 556124
rect 67726 556112 67732 556124
rect 67784 556112 67790 556164
rect 108942 556112 108948 556164
rect 109000 556152 109006 556164
rect 110598 556152 110604 556164
rect 109000 556124 110604 556152
rect 109000 556112 109006 556124
rect 110598 556112 110604 556124
rect 110656 556112 110662 556164
rect 110598 555432 110604 555484
rect 110656 555472 110662 555484
rect 116578 555472 116584 555484
rect 110656 555444 116584 555472
rect 110656 555432 110662 555444
rect 116578 555432 116584 555444
rect 116636 555432 116642 555484
rect 37182 554752 37188 554804
rect 37240 554792 37246 554804
rect 67634 554792 67640 554804
rect 37240 554764 67640 554792
rect 37240 554752 37246 554764
rect 67634 554752 67640 554764
rect 67692 554752 67698 554804
rect 141510 554004 141516 554056
rect 141568 554044 141574 554056
rect 159358 554044 159364 554056
rect 141568 554016 159364 554044
rect 141568 554004 141574 554016
rect 159358 554004 159364 554016
rect 159416 554004 159422 554056
rect 108850 553460 108856 553512
rect 108908 553500 108914 553512
rect 118970 553500 118976 553512
rect 108908 553472 118976 553500
rect 108908 553460 108914 553472
rect 118970 553460 118976 553472
rect 119028 553460 119034 553512
rect 50890 553392 50896 553444
rect 50948 553432 50954 553444
rect 67634 553432 67640 553444
rect 50948 553404 67640 553432
rect 50948 553392 50954 553404
rect 67634 553392 67640 553404
rect 67692 553392 67698 553444
rect 108942 553392 108948 553444
rect 109000 553432 109006 553444
rect 141510 553432 141516 553444
rect 109000 553404 141516 553432
rect 109000 553392 109006 553404
rect 141510 553392 141516 553404
rect 141568 553432 141574 553444
rect 142062 553432 142068 553444
rect 141568 553404 142068 553432
rect 141568 553392 141574 553404
rect 142062 553392 142068 553404
rect 142120 553392 142126 553444
rect 53742 552032 53748 552084
rect 53800 552072 53806 552084
rect 67634 552072 67640 552084
rect 53800 552044 67640 552072
rect 53800 552032 53806 552044
rect 67634 552032 67640 552044
rect 67692 552032 67698 552084
rect 108942 552032 108948 552084
rect 109000 552072 109006 552084
rect 124582 552072 124588 552084
rect 109000 552044 124588 552072
rect 109000 552032 109006 552044
rect 124582 552032 124588 552044
rect 124640 552032 124646 552084
rect 107838 551488 107844 551540
rect 107896 551528 107902 551540
rect 110598 551528 110604 551540
rect 107896 551500 110604 551528
rect 107896 551488 107902 551500
rect 110598 551488 110604 551500
rect 110656 551488 110662 551540
rect 38562 550604 38568 550656
rect 38620 550644 38626 550656
rect 67634 550644 67640 550656
rect 38620 550616 67640 550644
rect 38620 550604 38626 550616
rect 67634 550604 67640 550616
rect 67692 550604 67698 550656
rect 108942 550604 108948 550656
rect 109000 550644 109006 550656
rect 138106 550644 138112 550656
rect 109000 550616 138112 550644
rect 109000 550604 109006 550616
rect 138106 550604 138112 550616
rect 138164 550604 138170 550656
rect 108942 549312 108948 549364
rect 109000 549352 109006 549364
rect 132494 549352 132500 549364
rect 109000 549324 132500 549352
rect 109000 549312 109006 549324
rect 132494 549312 132500 549324
rect 132552 549312 132558 549364
rect 35710 549244 35716 549296
rect 35768 549284 35774 549296
rect 67634 549284 67640 549296
rect 35768 549256 67640 549284
rect 35768 549244 35774 549256
rect 67634 549244 67640 549256
rect 67692 549244 67698 549296
rect 108850 549244 108856 549296
rect 108908 549284 108914 549296
rect 142246 549284 142252 549296
rect 108908 549256 142252 549284
rect 108908 549244 108914 549256
rect 142246 549244 142252 549256
rect 142304 549244 142310 549296
rect 52270 547952 52276 548004
rect 52328 547992 52334 548004
rect 67634 547992 67640 548004
rect 52328 547964 67640 547992
rect 52328 547952 52334 547964
rect 67634 547952 67640 547964
rect 67692 547952 67698 548004
rect 39850 547884 39856 547936
rect 39908 547924 39914 547936
rect 67726 547924 67732 547936
rect 39908 547896 67732 547924
rect 39908 547884 39914 547896
rect 67726 547884 67732 547896
rect 67784 547884 67790 547936
rect 61930 546524 61936 546576
rect 61988 546564 61994 546576
rect 67726 546564 67732 546576
rect 61988 546536 67732 546564
rect 61988 546524 61994 546536
rect 67726 546524 67732 546536
rect 67784 546524 67790 546576
rect 60642 546456 60648 546508
rect 60700 546496 60706 546508
rect 67634 546496 67640 546508
rect 60700 546468 67640 546496
rect 60700 546456 60706 546468
rect 67634 546456 67640 546468
rect 67692 546456 67698 546508
rect 108942 546456 108948 546508
rect 109000 546496 109006 546508
rect 135254 546496 135260 546508
rect 109000 546468 135260 546496
rect 109000 546456 109006 546468
rect 135254 546456 135260 546468
rect 135312 546456 135318 546508
rect 108942 545708 108948 545760
rect 109000 545748 109006 545760
rect 113082 545748 113088 545760
rect 109000 545720 113088 545748
rect 109000 545708 109006 545720
rect 113082 545708 113088 545720
rect 113140 545748 113146 545760
rect 125778 545748 125784 545760
rect 113140 545720 125784 545748
rect 113140 545708 113146 545720
rect 125778 545708 125784 545720
rect 125836 545708 125842 545760
rect 110414 545164 110420 545216
rect 110472 545204 110478 545216
rect 111702 545204 111708 545216
rect 110472 545176 111708 545204
rect 110472 545164 110478 545176
rect 111702 545164 111708 545176
rect 111760 545204 111766 545216
rect 133966 545204 133972 545216
rect 111760 545176 133972 545204
rect 111760 545164 111766 545176
rect 133966 545164 133972 545176
rect 134024 545164 134030 545216
rect 35802 545096 35808 545148
rect 35860 545136 35866 545148
rect 68554 545136 68560 545148
rect 35860 545108 68560 545136
rect 35860 545096 35866 545108
rect 68554 545096 68560 545108
rect 68612 545096 68618 545148
rect 108942 545096 108948 545148
rect 109000 545136 109006 545148
rect 139486 545136 139492 545148
rect 109000 545108 139492 545136
rect 109000 545096 109006 545108
rect 139486 545096 139492 545108
rect 139544 545096 139550 545148
rect 108850 545028 108856 545080
rect 108908 545068 108914 545080
rect 110414 545068 110420 545080
rect 108908 545040 110420 545068
rect 108908 545028 108914 545040
rect 110414 545028 110420 545040
rect 110472 545028 110478 545080
rect 25498 544348 25504 544400
rect 25556 544388 25562 544400
rect 68002 544388 68008 544400
rect 25556 544360 68008 544388
rect 25556 544348 25562 544360
rect 68002 544348 68008 544360
rect 68060 544348 68066 544400
rect 63402 542444 63408 542496
rect 63460 542484 63466 542496
rect 67634 542484 67640 542496
rect 63460 542456 67640 542484
rect 63460 542444 63466 542456
rect 67634 542444 67640 542456
rect 67692 542444 67698 542496
rect 46842 542376 46848 542428
rect 46900 542416 46906 542428
rect 67726 542416 67732 542428
rect 46900 542388 67732 542416
rect 46900 542376 46906 542388
rect 67726 542376 67732 542388
rect 67784 542376 67790 542428
rect 108942 542376 108948 542428
rect 109000 542416 109006 542428
rect 136726 542416 136732 542428
rect 109000 542388 136732 542416
rect 109000 542376 109006 542388
rect 136726 542376 136732 542388
rect 136784 542376 136790 542428
rect 129734 541628 129740 541680
rect 129792 541668 129798 541680
rect 299474 541668 299480 541680
rect 129792 541640 299480 541668
rect 129792 541628 129798 541640
rect 299474 541628 299480 541640
rect 299532 541628 299538 541680
rect 109770 541016 109776 541068
rect 109828 541056 109834 541068
rect 129734 541056 129740 541068
rect 109828 541028 129740 541056
rect 109828 541016 109834 541028
rect 129734 541016 129740 541028
rect 129792 541016 129798 541068
rect 63310 540948 63316 541000
rect 63368 540988 63374 541000
rect 67634 540988 67640 541000
rect 63368 540960 67640 540988
rect 63368 540948 63374 540960
rect 67634 540948 67640 540960
rect 67692 540948 67698 541000
rect 108942 540948 108948 541000
rect 109000 540988 109006 541000
rect 142338 540988 142344 541000
rect 109000 540960 142344 540988
rect 109000 540948 109006 540960
rect 142338 540948 142344 540960
rect 142396 540948 142402 541000
rect 107470 540880 107476 540932
rect 107528 540920 107534 540932
rect 109678 540920 109684 540932
rect 107528 540892 109684 540920
rect 107528 540880 107534 540892
rect 109678 540880 109684 540892
rect 109736 540880 109742 540932
rect 62022 539588 62028 539640
rect 62080 539628 62086 539640
rect 67634 539628 67640 539640
rect 62080 539600 67640 539628
rect 62080 539588 62086 539600
rect 67634 539588 67640 539600
rect 67692 539588 67698 539640
rect 4798 539520 4804 539572
rect 4856 539560 4862 539572
rect 99006 539560 99012 539572
rect 4856 539532 99012 539560
rect 4856 539520 4862 539532
rect 99006 539520 99012 539532
rect 99064 539520 99070 539572
rect 95142 539112 95148 539164
rect 95200 539152 95206 539164
rect 118786 539152 118792 539164
rect 95200 539124 118792 539152
rect 95200 539112 95206 539124
rect 118786 539112 118792 539124
rect 118844 539112 118850 539164
rect 97902 539044 97908 539096
rect 97960 539084 97966 539096
rect 113358 539084 113364 539096
rect 97960 539056 113364 539084
rect 97960 539044 97966 539056
rect 113358 539044 113364 539056
rect 113416 539044 113422 539096
rect 59078 538976 59084 539028
rect 59136 539016 59142 539028
rect 73154 539016 73160 539028
rect 59136 538988 73160 539016
rect 59136 538976 59142 538988
rect 73154 538976 73160 538988
rect 73212 538976 73218 539028
rect 88058 538976 88064 539028
rect 88116 539016 88122 539028
rect 118786 539016 118792 539028
rect 88116 538988 118792 539016
rect 88116 538976 88122 538988
rect 118786 538976 118792 538988
rect 118844 539016 118850 539028
rect 126238 539016 126244 539028
rect 118844 538988 126244 539016
rect 118844 538976 118850 538988
rect 126238 538976 126244 538988
rect 126296 538976 126302 539028
rect 57698 538908 57704 538960
rect 57756 538948 57762 538960
rect 90358 538948 90364 538960
rect 57756 538920 90364 538948
rect 57756 538908 57762 538920
rect 90358 538908 90364 538920
rect 90416 538908 90422 538960
rect 98638 538908 98644 538960
rect 98696 538948 98702 538960
rect 120166 538948 120172 538960
rect 98696 538920 120172 538948
rect 98696 538908 98702 538920
rect 120166 538908 120172 538920
rect 120224 538908 120230 538960
rect 54478 538840 54484 538892
rect 54536 538880 54542 538892
rect 57882 538880 57888 538892
rect 54536 538852 57888 538880
rect 54536 538840 54542 538852
rect 57882 538840 57888 538852
rect 57940 538880 57946 538892
rect 91278 538880 91284 538892
rect 57940 538852 91284 538880
rect 57940 538840 57946 538852
rect 91278 538840 91284 538852
rect 91336 538840 91342 538892
rect 99006 538840 99012 538892
rect 99064 538880 99070 538892
rect 124490 538880 124496 538892
rect 99064 538852 124496 538880
rect 99064 538840 99070 538852
rect 124490 538840 124496 538852
rect 124548 538840 124554 538892
rect 15838 538160 15844 538212
rect 15896 538200 15902 538212
rect 98362 538200 98368 538212
rect 15896 538172 98368 538200
rect 15896 538160 15902 538172
rect 98362 538160 98368 538172
rect 98420 538160 98426 538212
rect 103514 538160 103520 538212
rect 103572 538200 103578 538212
rect 109770 538200 109776 538212
rect 103572 538172 109776 538200
rect 103572 538160 103578 538172
rect 109770 538160 109776 538172
rect 109828 538160 109834 538212
rect 155218 538160 155224 538212
rect 155276 538200 155282 538212
rect 580166 538200 580172 538212
rect 155276 538172 580172 538200
rect 155276 538160 155282 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 102226 537752 102232 537804
rect 102284 537792 102290 537804
rect 110782 537792 110788 537804
rect 102284 537764 110788 537792
rect 102284 537752 102290 537764
rect 110782 537752 110788 537764
rect 110840 537752 110846 537804
rect 70302 537684 70308 537736
rect 70360 537724 70366 537736
rect 81526 537724 81532 537736
rect 70360 537696 81532 537724
rect 70360 537684 70366 537696
rect 81526 537684 81532 537696
rect 81584 537684 81590 537736
rect 102870 537684 102876 537736
rect 102928 537724 102934 537736
rect 127618 537724 127624 537736
rect 102928 537696 127624 537724
rect 102928 537684 102934 537696
rect 127618 537684 127624 537696
rect 127676 537684 127682 537736
rect 45370 537616 45376 537668
rect 45428 537656 45434 537668
rect 56410 537656 56416 537668
rect 45428 537628 56416 537656
rect 45428 537616 45434 537628
rect 56410 537616 56416 537628
rect 56468 537616 56474 537668
rect 57698 537616 57704 537668
rect 57756 537656 57762 537668
rect 81618 537656 81624 537668
rect 57756 537628 81624 537656
rect 57756 537616 57762 537628
rect 81618 537616 81624 537628
rect 81676 537616 81682 537668
rect 83458 537616 83464 537668
rect 83516 537656 83522 537668
rect 90634 537656 90640 537668
rect 83516 537628 90640 537656
rect 83516 537616 83522 537628
rect 90634 537616 90640 537628
rect 90692 537616 90698 537668
rect 98362 537616 98368 537668
rect 98420 537656 98426 537668
rect 122926 537656 122932 537668
rect 98420 537628 122932 537656
rect 98420 537616 98426 537628
rect 122926 537616 122932 537628
rect 122984 537616 122990 537668
rect 44082 537548 44088 537600
rect 44140 537588 44146 537600
rect 73246 537588 73252 537600
rect 44140 537560 73252 537588
rect 44140 537548 44146 537560
rect 73246 537548 73252 537560
rect 73304 537548 73310 537600
rect 79686 537548 79692 537600
rect 79744 537588 79750 537600
rect 87046 537588 87052 537600
rect 79744 537560 87052 537588
rect 79744 537548 79750 537560
rect 87046 537548 87052 537560
rect 87104 537548 87110 537600
rect 95786 537548 95792 537600
rect 95844 537588 95850 537600
rect 121546 537588 121552 537600
rect 95844 537560 121552 537588
rect 95844 537548 95850 537560
rect 121546 537548 121552 537560
rect 121604 537548 121610 537600
rect 52086 537480 52092 537532
rect 52144 537520 52150 537532
rect 82906 537520 82912 537532
rect 52144 537492 82912 537520
rect 52144 537480 52150 537492
rect 82906 537480 82912 537492
rect 82964 537480 82970 537532
rect 84194 537480 84200 537532
rect 84252 537520 84258 537532
rect 98546 537520 98552 537532
rect 84252 537492 98552 537520
rect 84252 537480 84258 537492
rect 98546 537480 98552 537492
rect 98604 537480 98610 537532
rect 100294 537480 100300 537532
rect 100352 537520 100358 537532
rect 132586 537520 132592 537532
rect 100352 537492 132592 537520
rect 100352 537480 100358 537492
rect 132586 537480 132592 537492
rect 132644 537480 132650 537532
rect 94498 537412 94504 537464
rect 94556 537452 94562 537464
rect 100754 537452 100760 537464
rect 94556 537424 100760 537452
rect 94556 537412 94562 537424
rect 100754 537412 100760 537424
rect 100812 537412 100818 537464
rect 70210 536800 70216 536852
rect 70268 536840 70274 536852
rect 75086 536840 75092 536852
rect 70268 536812 75092 536840
rect 70268 536800 70274 536812
rect 75086 536800 75092 536812
rect 75144 536800 75150 536852
rect 84102 536800 84108 536852
rect 84160 536840 84166 536852
rect 84838 536840 84844 536852
rect 84160 536812 84844 536840
rect 84160 536800 84166 536812
rect 84838 536800 84844 536812
rect 84896 536800 84902 536852
rect 102042 536800 102048 536852
rect 102100 536840 102106 536852
rect 104158 536840 104164 536852
rect 102100 536812 104164 536840
rect 102100 536800 102106 536812
rect 104158 536800 104164 536812
rect 104216 536800 104222 536852
rect 35158 536732 35164 536784
rect 35216 536772 35222 536784
rect 106274 536772 106280 536784
rect 35216 536744 106280 536772
rect 35216 536732 35222 536744
rect 106274 536732 106280 536744
rect 106332 536732 106338 536784
rect 100754 536664 100760 536716
rect 100812 536704 100818 536716
rect 118878 536704 118884 536716
rect 100812 536676 118884 536704
rect 100812 536664 100818 536676
rect 118878 536664 118884 536676
rect 118936 536664 118942 536716
rect 97810 536120 97816 536172
rect 97868 536160 97874 536172
rect 110506 536160 110512 536172
rect 97868 536132 110512 536160
rect 97868 536120 97874 536132
rect 110506 536120 110512 536132
rect 110564 536120 110570 536172
rect 118878 536120 118884 536172
rect 118936 536160 118942 536172
rect 128538 536160 128544 536172
rect 118936 536132 128544 536160
rect 118936 536120 118942 536132
rect 128538 536120 128544 536132
rect 128596 536120 128602 536172
rect 106274 536052 106280 536104
rect 106332 536092 106338 536104
rect 131206 536092 131212 536104
rect 106332 536064 131212 536092
rect 106332 536052 106338 536064
rect 131206 536052 131212 536064
rect 131264 536052 131270 536104
rect 71038 535372 71044 535424
rect 71096 535412 71102 535424
rect 77110 535412 77116 535424
rect 71096 535384 77116 535412
rect 71096 535372 71102 535384
rect 77110 535372 77116 535384
rect 77168 535372 77174 535424
rect 48130 534828 48136 534880
rect 48188 534868 48194 534880
rect 75178 534868 75184 534880
rect 48188 534840 75184 534868
rect 48188 534828 48194 534840
rect 75178 534828 75184 534840
rect 75236 534828 75242 534880
rect 99282 534828 99288 534880
rect 99340 534868 99346 534880
rect 114646 534868 114652 534880
rect 99340 534840 114652 534868
rect 99340 534828 99346 534840
rect 114646 534828 114652 534840
rect 114704 534828 114710 534880
rect 115198 534828 115204 534880
rect 115256 534868 115262 534880
rect 128354 534868 128360 534880
rect 115256 534840 128360 534868
rect 115256 534828 115262 534840
rect 128354 534828 128360 534840
rect 128412 534828 128418 534880
rect 53558 534760 53564 534812
rect 53616 534800 53622 534812
rect 83550 534800 83556 534812
rect 53616 534772 83556 534800
rect 53616 534760 53622 534772
rect 83550 534760 83556 534772
rect 83608 534760 83614 534812
rect 93854 534760 93860 534812
rect 93912 534800 93918 534812
rect 120166 534800 120172 534812
rect 93912 534772 120172 534800
rect 93912 534760 93918 534772
rect 120166 534760 120172 534772
rect 120224 534760 120230 534812
rect 46566 534692 46572 534744
rect 46624 534732 46630 534744
rect 78398 534732 78404 534744
rect 46624 534704 78404 534732
rect 46624 534692 46630 534704
rect 78398 534692 78404 534704
rect 78456 534692 78462 534744
rect 89990 534692 89996 534744
rect 90048 534732 90054 534744
rect 118878 534732 118884 534744
rect 90048 534704 118884 534732
rect 90048 534692 90054 534704
rect 118878 534692 118884 534704
rect 118936 534692 118942 534744
rect 46750 533332 46756 533384
rect 46808 533372 46814 533384
rect 76558 533372 76564 533384
rect 46808 533344 76564 533372
rect 46808 533332 46814 533344
rect 76558 533332 76564 533344
rect 76616 533332 76622 533384
rect 49510 532108 49516 532160
rect 49568 532148 49574 532160
rect 76466 532148 76472 532160
rect 49568 532120 76472 532148
rect 49568 532108 49574 532120
rect 76466 532108 76472 532120
rect 76524 532108 76530 532160
rect 97074 532108 97080 532160
rect 97132 532148 97138 532160
rect 121730 532148 121736 532160
rect 97132 532120 121736 532148
rect 97132 532108 97138 532120
rect 121730 532108 121736 532120
rect 121788 532108 121794 532160
rect 52362 532040 52368 532092
rect 52420 532080 52426 532092
rect 79318 532080 79324 532092
rect 52420 532052 79324 532080
rect 52420 532040 52426 532052
rect 79318 532040 79324 532052
rect 79376 532040 79382 532092
rect 87414 532040 87420 532092
rect 87472 532080 87478 532092
rect 109218 532080 109224 532092
rect 87472 532052 109224 532080
rect 87472 532040 87478 532052
rect 109218 532040 109224 532052
rect 109276 532040 109282 532092
rect 54938 531972 54944 532024
rect 54996 532012 55002 532024
rect 86126 532012 86132 532024
rect 54996 531984 86132 532012
rect 54996 531972 55002 531984
rect 86126 531972 86132 531984
rect 86184 531972 86190 532024
rect 95050 531972 95056 532024
rect 95108 532012 95114 532024
rect 121638 532012 121644 532024
rect 95108 531984 121644 532012
rect 95108 531972 95114 531984
rect 121638 531972 121644 531984
rect 121696 531972 121702 532024
rect 56410 529320 56416 529372
rect 56468 529360 56474 529372
rect 72602 529360 72608 529372
rect 56468 529332 72608 529360
rect 56468 529320 56474 529332
rect 72602 529320 72608 529332
rect 72660 529320 72666 529372
rect 46658 529252 46664 529304
rect 46716 529292 46722 529304
rect 70486 529292 70492 529304
rect 46716 529264 70492 529292
rect 46716 529252 46722 529264
rect 70486 529252 70492 529264
rect 70544 529252 70550 529304
rect 40954 529184 40960 529236
rect 41012 529224 41018 529236
rect 74534 529224 74540 529236
rect 41012 529196 74540 529224
rect 41012 529184 41018 529196
rect 74534 529184 74540 529196
rect 74592 529184 74598 529236
rect 110414 529184 110420 529236
rect 110472 529224 110478 529236
rect 110598 529224 110604 529236
rect 110472 529196 110604 529224
rect 110472 529184 110478 529196
rect 110598 529184 110604 529196
rect 110656 529224 110662 529236
rect 128354 529224 128360 529236
rect 110656 529196 128360 529224
rect 110656 529184 110662 529196
rect 128354 529184 128360 529196
rect 128412 529184 128418 529236
rect 110414 528612 110420 528624
rect 106246 528584 110420 528612
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 106246 528544 106274 528584
rect 110414 528572 110420 528584
rect 110472 528572 110478 528624
rect 3200 528516 106274 528544
rect 3200 528504 3206 528516
rect 39666 526396 39672 526448
rect 39724 526436 39730 526448
rect 71958 526436 71964 526448
rect 39724 526408 71964 526436
rect 39724 526396 39730 526408
rect 71958 526396 71964 526408
rect 72016 526396 72022 526448
rect 34238 525784 34244 525836
rect 34296 525824 34302 525836
rect 34296 525796 64874 525824
rect 34296 525784 34302 525796
rect 64846 525756 64874 525796
rect 69014 525756 69020 525768
rect 64846 525728 69020 525756
rect 69014 525716 69020 525728
rect 69072 525756 69078 525768
rect 579798 525756 579804 525768
rect 69072 525728 579804 525756
rect 69072 525716 69078 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 431218 510620 431224 510672
rect 431276 510660 431282 510672
rect 580166 510660 580172 510672
rect 431276 510632 580172 510660
rect 431276 510620 431282 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 88242 500284 88248 500336
rect 88300 500324 88306 500336
rect 117406 500324 117412 500336
rect 88300 500296 117412 500324
rect 88300 500284 88306 500296
rect 117406 500284 117412 500296
rect 117464 500324 117470 500336
rect 125594 500324 125600 500336
rect 117464 500296 125600 500324
rect 117464 500284 117470 500296
rect 125594 500284 125600 500296
rect 125652 500284 125658 500336
rect 95234 500216 95240 500268
rect 95292 500256 95298 500268
rect 136818 500256 136824 500268
rect 95292 500228 136824 500256
rect 95292 500216 95298 500228
rect 136818 500216 136824 500228
rect 136876 500256 136882 500268
rect 137094 500256 137100 500268
rect 136876 500228 137100 500256
rect 136876 500216 136882 500228
rect 137094 500216 137100 500228
rect 137152 500216 137158 500268
rect 89346 498788 89352 498840
rect 89404 498828 89410 498840
rect 111794 498828 111800 498840
rect 89404 498800 111800 498828
rect 89404 498788 89410 498800
rect 111794 498788 111800 498800
rect 111852 498788 111858 498840
rect 85482 497564 85488 497616
rect 85540 497604 85546 497616
rect 109310 497604 109316 497616
rect 85540 497576 109316 497604
rect 85540 497564 85546 497576
rect 109310 497564 109316 497576
rect 109368 497564 109374 497616
rect 84102 497496 84108 497548
rect 84160 497536 84166 497548
rect 110414 497536 110420 497548
rect 84160 497508 110420 497536
rect 84160 497496 84166 497508
rect 110414 497496 110420 497508
rect 110472 497496 110478 497548
rect 38470 497428 38476 497480
rect 38528 497468 38534 497480
rect 70394 497468 70400 497480
rect 38528 497440 70400 497468
rect 38528 497428 38534 497440
rect 70394 497428 70400 497440
rect 70452 497428 70458 497480
rect 81618 497428 81624 497480
rect 81676 497468 81682 497480
rect 88242 497468 88248 497480
rect 81676 497440 88248 497468
rect 81676 497428 81682 497440
rect 88242 497428 88248 497440
rect 88300 497428 88306 497480
rect 96430 497428 96436 497480
rect 96488 497468 96494 497480
rect 131298 497468 131304 497480
rect 96488 497440 131304 497468
rect 96488 497428 96494 497440
rect 131298 497428 131304 497440
rect 131356 497428 131362 497480
rect 88058 496272 88064 496324
rect 88116 496312 88122 496324
rect 123110 496312 123116 496324
rect 88116 496284 123116 496312
rect 88116 496272 88122 496284
rect 123110 496272 123116 496284
rect 123168 496312 123174 496324
rect 123168 496284 132494 496312
rect 123168 496272 123174 496284
rect 89622 496204 89628 496256
rect 89680 496244 89686 496256
rect 125686 496244 125692 496256
rect 89680 496216 125692 496244
rect 89680 496204 89686 496216
rect 125686 496204 125692 496216
rect 125744 496244 125750 496256
rect 127066 496244 127072 496256
rect 125744 496216 127072 496244
rect 125744 496204 125750 496216
rect 127066 496204 127072 496216
rect 127124 496204 127130 496256
rect 76466 496136 76472 496188
rect 76524 496176 76530 496188
rect 81526 496176 81532 496188
rect 76524 496148 81532 496176
rect 76524 496136 76530 496148
rect 81526 496136 81532 496148
rect 81584 496176 81590 496188
rect 123294 496176 123300 496188
rect 81584 496148 123300 496176
rect 81584 496136 81590 496148
rect 123294 496136 123300 496148
rect 123352 496136 123358 496188
rect 4798 496068 4804 496120
rect 4856 496108 4862 496120
rect 91094 496108 91100 496120
rect 4856 496080 91100 496108
rect 4856 496068 4862 496080
rect 91094 496068 91100 496080
rect 91152 496068 91158 496120
rect 132466 496108 132494 496284
rect 135346 496108 135352 496120
rect 132466 496080 135352 496108
rect 135346 496068 135352 496080
rect 135404 496068 135410 496120
rect 91094 495456 91100 495508
rect 91152 495496 91158 495508
rect 116026 495496 116032 495508
rect 91152 495468 116032 495496
rect 91152 495456 91158 495468
rect 116026 495456 116032 495468
rect 116084 495496 116090 495508
rect 116394 495496 116400 495508
rect 116084 495468 116400 495496
rect 116084 495456 116090 495468
rect 116394 495456 116400 495468
rect 116452 495456 116458 495508
rect 93210 494980 93216 495032
rect 93268 495020 93274 495032
rect 112162 495020 112168 495032
rect 93268 494992 112168 495020
rect 93268 494980 93274 494992
rect 112162 494980 112168 494992
rect 112220 494980 112226 495032
rect 58986 494844 58992 494896
rect 59044 494884 59050 494896
rect 80974 494884 80980 494896
rect 59044 494856 80980 494884
rect 59044 494844 59050 494856
rect 80974 494844 80980 494856
rect 81032 494844 81038 494896
rect 82262 494844 82268 494896
rect 82320 494884 82326 494896
rect 111978 494884 111984 494896
rect 82320 494856 111984 494884
rect 82320 494844 82326 494856
rect 111978 494844 111984 494856
rect 112036 494884 112042 494896
rect 119062 494884 119068 494896
rect 112036 494856 119068 494884
rect 112036 494844 112042 494856
rect 119062 494844 119068 494856
rect 119120 494844 119126 494896
rect 43898 494776 43904 494828
rect 43956 494816 43962 494828
rect 49602 494816 49608 494828
rect 43956 494788 49608 494816
rect 43956 494776 43962 494788
rect 49602 494776 49608 494788
rect 49660 494816 49666 494828
rect 75454 494816 75460 494828
rect 49660 494788 75460 494816
rect 49660 494776 49666 494788
rect 75454 494776 75460 494788
rect 75512 494776 75518 494828
rect 82906 494776 82912 494828
rect 82964 494816 82970 494828
rect 123018 494816 123024 494828
rect 82964 494788 123024 494816
rect 82964 494776 82970 494788
rect 123018 494776 123024 494788
rect 123076 494816 123082 494828
rect 127250 494816 127256 494828
rect 123076 494788 127256 494816
rect 123076 494776 123082 494788
rect 127250 494776 127256 494788
rect 127308 494776 127314 494828
rect 3510 494708 3516 494760
rect 3568 494748 3574 494760
rect 82814 494748 82820 494760
rect 3568 494720 82820 494748
rect 3568 494708 3574 494720
rect 82814 494708 82820 494720
rect 82872 494708 82878 494760
rect 90634 494708 90640 494760
rect 90692 494748 90698 494760
rect 118694 494748 118700 494760
rect 90692 494720 118700 494748
rect 90692 494708 90698 494720
rect 118694 494708 118700 494720
rect 118752 494748 118758 494760
rect 134058 494748 134064 494760
rect 118752 494720 134064 494748
rect 118752 494708 118758 494720
rect 134058 494708 134064 494720
rect 134116 494708 134122 494760
rect 47854 494504 47860 494556
rect 47912 494544 47918 494556
rect 48038 494544 48044 494556
rect 47912 494516 48044 494544
rect 47912 494504 47918 494516
rect 48038 494504 48044 494516
rect 48096 494504 48102 494556
rect 47854 494028 47860 494080
rect 47912 494068 47918 494080
rect 77386 494068 77392 494080
rect 47912 494040 77392 494068
rect 47912 494028 47918 494040
rect 77386 494028 77392 494040
rect 77444 494028 77450 494080
rect 82814 493960 82820 494012
rect 82872 494000 82878 494012
rect 83550 494000 83556 494012
rect 82872 493972 83556 494000
rect 82872 493960 82878 493972
rect 83550 493960 83556 493972
rect 83608 494000 83614 494012
rect 121454 494000 121460 494012
rect 83608 493972 121460 494000
rect 83608 493960 83614 493972
rect 121454 493960 121460 493972
rect 121512 493960 121518 494012
rect 120074 493892 120080 493944
rect 120132 493932 120138 493944
rect 121822 493932 121828 493944
rect 120132 493904 121828 493932
rect 120132 493892 120138 493904
rect 121822 493892 121828 493904
rect 121880 493892 121886 493944
rect 88702 493824 88708 493876
rect 88760 493864 88766 493876
rect 89530 493864 89536 493876
rect 88760 493836 89536 493864
rect 88760 493824 88766 493836
rect 89530 493824 89536 493836
rect 89588 493824 89594 493876
rect 110506 493552 110512 493604
rect 110564 493592 110570 493604
rect 110690 493592 110696 493604
rect 110564 493564 110696 493592
rect 110564 493552 110570 493564
rect 110690 493552 110696 493564
rect 110748 493592 110754 493604
rect 124398 493592 124404 493604
rect 110748 493564 124404 493592
rect 110748 493552 110754 493564
rect 124398 493552 124404 493564
rect 124456 493552 124462 493604
rect 97718 493484 97724 493536
rect 97776 493524 97782 493536
rect 114738 493524 114744 493536
rect 97776 493496 114744 493524
rect 97776 493484 97782 493496
rect 114738 493484 114744 493496
rect 114796 493484 114802 493536
rect 95142 493416 95148 493468
rect 95200 493456 95206 493468
rect 113266 493456 113272 493468
rect 95200 493428 113272 493456
rect 95200 493416 95206 493428
rect 113266 493416 113272 493428
rect 113324 493456 113330 493468
rect 113324 493428 116440 493456
rect 113324 493416 113330 493428
rect 93210 493348 93216 493400
rect 93268 493388 93274 493400
rect 93268 493360 113174 493388
rect 93268 493348 93274 493360
rect 54754 493280 54760 493332
rect 54812 493320 54818 493332
rect 59170 493320 59176 493332
rect 54812 493292 59176 493320
rect 54812 493280 54818 493292
rect 59170 493280 59176 493292
rect 59228 493320 59234 493332
rect 70026 493320 70032 493332
rect 59228 493292 70032 493320
rect 59228 493280 59234 493292
rect 70026 493280 70032 493292
rect 70084 493280 70090 493332
rect 80974 493280 80980 493332
rect 81032 493320 81038 493332
rect 110506 493320 110512 493332
rect 81032 493292 110512 493320
rect 81032 493280 81038 493292
rect 110506 493280 110512 493292
rect 110564 493280 110570 493332
rect 113146 493252 113174 493360
rect 116412 493320 116440 493428
rect 121454 493348 121460 493400
rect 121512 493388 121518 493400
rect 128446 493388 128452 493400
rect 121512 493360 128452 493388
rect 121512 493348 121518 493360
rect 128446 493348 128452 493360
rect 128504 493348 128510 493400
rect 137278 493320 137284 493332
rect 116412 493292 137284 493320
rect 137278 493280 137284 493292
rect 137336 493280 137342 493332
rect 120074 493252 120080 493264
rect 113146 493224 120080 493252
rect 120074 493212 120080 493224
rect 120132 493212 120138 493264
rect 85482 493144 85488 493196
rect 85540 493184 85546 493196
rect 89622 493184 89628 493196
rect 85540 493156 89628 493184
rect 85540 493144 85546 493156
rect 89622 493144 89628 493156
rect 89680 493144 89686 493196
rect 47946 492668 47952 492720
rect 48004 492708 48010 492720
rect 71130 492708 71136 492720
rect 48004 492680 71136 492708
rect 48004 492668 48010 492680
rect 71130 492668 71136 492680
rect 71188 492668 71194 492720
rect 88702 492668 88708 492720
rect 88760 492708 88766 492720
rect 102134 492708 102140 492720
rect 88760 492680 102140 492708
rect 88760 492668 88766 492680
rect 102134 492668 102140 492680
rect 102192 492668 102198 492720
rect 75178 492600 75184 492652
rect 75236 492640 75242 492652
rect 78398 492640 78404 492652
rect 75236 492612 78404 492640
rect 75236 492600 75242 492612
rect 78398 492600 78404 492612
rect 78456 492600 78462 492652
rect 39942 492056 39948 492108
rect 40000 492096 40006 492108
rect 45462 492096 45468 492108
rect 40000 492068 45468 492096
rect 40000 492056 40006 492068
rect 45462 492056 45468 492068
rect 45520 492096 45526 492108
rect 72234 492096 72240 492108
rect 45520 492068 72240 492096
rect 45520 492056 45526 492068
rect 72234 492056 72240 492068
rect 72292 492056 72298 492108
rect 49602 491988 49608 492040
rect 49660 492028 49666 492040
rect 53098 492028 53104 492040
rect 49660 492000 53104 492028
rect 49660 491988 49666 492000
rect 53098 491988 53104 492000
rect 53156 492028 53162 492040
rect 80054 492028 80060 492040
rect 53156 492000 80060 492028
rect 53156 491988 53162 492000
rect 80054 491988 80060 492000
rect 80112 491988 80118 492040
rect 91922 491988 91928 492040
rect 91980 492028 91986 492040
rect 97902 492028 97908 492040
rect 91980 492000 97908 492028
rect 91980 491988 91986 492000
rect 97902 491988 97908 492000
rect 97960 492028 97966 492040
rect 101398 492028 101404 492040
rect 97960 492000 101404 492028
rect 97960 491988 97966 492000
rect 101398 491988 101404 492000
rect 101456 491988 101462 492040
rect 56226 491920 56232 491972
rect 56284 491960 56290 491972
rect 83458 491960 83464 491972
rect 56284 491932 83464 491960
rect 56284 491920 56290 491932
rect 83458 491920 83464 491932
rect 83516 491920 83522 491972
rect 86126 491920 86132 491972
rect 86184 491960 86190 491972
rect 96982 491960 96988 491972
rect 86184 491932 96988 491960
rect 86184 491920 86190 491932
rect 96982 491920 96988 491932
rect 97040 491920 97046 491972
rect 98362 491920 98368 491972
rect 98420 491960 98426 491972
rect 126974 491960 126980 491972
rect 98420 491932 126980 491960
rect 98420 491920 98426 491932
rect 126974 491920 126980 491932
rect 127032 491960 127038 491972
rect 139394 491960 139400 491972
rect 127032 491932 139400 491960
rect 127032 491920 127038 491932
rect 139394 491920 139400 491932
rect 139452 491920 139458 491972
rect 78398 491648 78404 491700
rect 78456 491688 78462 491700
rect 103606 491688 103612 491700
rect 78456 491660 103612 491688
rect 78456 491648 78462 491660
rect 103606 491648 103612 491660
rect 103664 491648 103670 491700
rect 76650 491580 76656 491632
rect 76708 491620 76714 491632
rect 113266 491620 113272 491632
rect 76708 491592 113272 491620
rect 76708 491580 76714 491592
rect 113266 491580 113272 491592
rect 113324 491580 113330 491632
rect 99650 491512 99656 491564
rect 99708 491552 99714 491564
rect 114554 491552 114560 491564
rect 99708 491524 114560 491552
rect 99708 491512 99714 491524
rect 114554 491512 114560 491524
rect 114612 491552 114618 491564
rect 114612 491524 115888 491552
rect 114612 491512 114618 491524
rect 90358 491444 90364 491496
rect 90416 491484 90422 491496
rect 110598 491484 110604 491496
rect 90416 491456 110604 491484
rect 90416 491444 90422 491456
rect 110598 491444 110604 491456
rect 110656 491444 110662 491496
rect 58618 491376 58624 491428
rect 58676 491416 58682 491428
rect 70394 491416 70400 491428
rect 58676 491388 70400 491416
rect 58676 491376 58682 491388
rect 70394 491376 70400 491388
rect 70452 491376 70458 491428
rect 86770 491376 86776 491428
rect 86828 491416 86834 491428
rect 92474 491416 92480 491428
rect 86828 491388 92480 491416
rect 86828 491376 86834 491388
rect 92474 491376 92480 491388
rect 92532 491376 92538 491428
rect 41230 491308 41236 491360
rect 41288 491348 41294 491360
rect 71774 491348 71780 491360
rect 41288 491320 71780 491348
rect 41288 491308 41294 491320
rect 71774 491308 71780 491320
rect 71832 491308 71838 491360
rect 50798 491240 50804 491292
rect 50856 491280 50862 491292
rect 58618 491280 58624 491292
rect 50856 491252 58624 491280
rect 50856 491240 50862 491252
rect 58618 491240 58624 491252
rect 58676 491240 58682 491292
rect 107562 491240 107568 491292
rect 107620 491280 107626 491292
rect 109034 491280 109040 491292
rect 107620 491252 109040 491280
rect 107620 491240 107626 491252
rect 109034 491240 109040 491252
rect 109092 491240 109098 491292
rect 115860 491212 115888 491524
rect 116394 491240 116400 491292
rect 116452 491280 116458 491292
rect 120074 491280 120080 491292
rect 116452 491252 120080 491280
rect 116452 491240 116458 491252
rect 120074 491240 120080 491252
rect 120132 491240 120138 491292
rect 120350 491212 120356 491224
rect 115860 491184 120356 491212
rect 120350 491172 120356 491184
rect 120408 491172 120414 491224
rect 87414 490696 87420 490748
rect 87472 490736 87478 490748
rect 95050 490736 95056 490748
rect 87472 490708 95056 490736
rect 87472 490696 87478 490708
rect 95050 490696 95056 490708
rect 95108 490736 95114 490748
rect 100018 490736 100024 490748
rect 95108 490708 100024 490736
rect 95108 490696 95114 490708
rect 100018 490696 100024 490708
rect 100076 490696 100082 490748
rect 92842 490628 92848 490680
rect 92900 490668 92906 490680
rect 107562 490668 107568 490680
rect 92900 490640 107568 490668
rect 92900 490628 92906 490640
rect 107562 490628 107568 490640
rect 107620 490628 107626 490680
rect 50798 490560 50804 490612
rect 50856 490600 50862 490612
rect 79042 490600 79048 490612
rect 50856 490572 79048 490600
rect 50856 490560 50862 490572
rect 79042 490560 79048 490572
rect 79100 490560 79106 490612
rect 92014 490560 92020 490612
rect 92072 490600 92078 490612
rect 109402 490600 109408 490612
rect 92072 490572 109408 490600
rect 92072 490560 92078 490572
rect 109402 490560 109408 490572
rect 109460 490560 109466 490612
rect 42610 489948 42616 490000
rect 42668 489988 42674 490000
rect 74350 489988 74356 490000
rect 42668 489960 74356 489988
rect 42668 489948 42674 489960
rect 74350 489948 74356 489960
rect 74408 489948 74414 490000
rect 45278 489880 45284 489932
rect 45336 489920 45342 489932
rect 73430 489920 73436 489932
rect 45336 489892 73436 489920
rect 45336 489880 45342 489892
rect 73430 489880 73436 489892
rect 73488 489880 73494 489932
rect 43806 489812 43812 489864
rect 43864 489852 43870 489864
rect 69014 489852 69020 489864
rect 43864 489824 69020 489852
rect 43864 489812 43870 489824
rect 69014 489812 69020 489824
rect 69072 489812 69078 489864
rect 97994 489812 98000 489864
rect 98052 489852 98058 489864
rect 98638 489852 98644 489864
rect 98052 489824 98644 489852
rect 98052 489812 98058 489824
rect 98638 489812 98644 489824
rect 98696 489852 98702 489864
rect 99190 489852 99196 489864
rect 98696 489824 99196 489852
rect 98696 489812 98702 489824
rect 99190 489812 99196 489824
rect 99248 489812 99254 489864
rect 101214 489812 101220 489864
rect 101272 489852 101278 489864
rect 117314 489852 117320 489864
rect 101272 489824 117320 489852
rect 101272 489812 101278 489824
rect 117314 489812 117320 489824
rect 117372 489812 117378 489864
rect 102226 489268 102232 489320
rect 102284 489308 102290 489320
rect 115198 489308 115204 489320
rect 102284 489280 115204 489308
rect 102284 489268 102290 489280
rect 115198 489268 115204 489280
rect 115256 489268 115262 489320
rect 99190 489200 99196 489252
rect 99248 489240 99254 489252
rect 113818 489240 113824 489252
rect 99248 489212 113824 489240
rect 99248 489200 99254 489212
rect 113818 489200 113824 489212
rect 113876 489200 113882 489252
rect 106182 489132 106188 489184
rect 106240 489172 106246 489184
rect 134150 489172 134156 489184
rect 106240 489144 134156 489172
rect 106240 489132 106246 489144
rect 134150 489132 134156 489144
rect 134208 489172 134214 489184
rect 151814 489172 151820 489184
rect 134208 489144 151820 489172
rect 134208 489132 134214 489144
rect 151814 489132 151820 489144
rect 151872 489132 151878 489184
rect 53650 488452 53656 488504
rect 53708 488492 53714 488504
rect 67634 488492 67640 488504
rect 53708 488464 67640 488492
rect 53708 488452 53714 488464
rect 67634 488452 67640 488464
rect 67692 488452 67698 488504
rect 102318 488452 102324 488504
rect 102376 488492 102382 488504
rect 109126 488492 109132 488504
rect 102376 488464 109132 488492
rect 102376 488452 102382 488464
rect 109126 488452 109132 488464
rect 109184 488452 109190 488504
rect 102226 488044 102232 488096
rect 102284 488084 102290 488096
rect 106182 488084 106188 488096
rect 102284 488056 106188 488084
rect 102284 488044 102290 488056
rect 106182 488044 106188 488056
rect 106240 488044 106246 488096
rect 48222 487772 48228 487824
rect 48280 487812 48286 487824
rect 67634 487812 67640 487824
rect 48280 487784 67640 487812
rect 48280 487772 48286 487784
rect 67634 487772 67640 487784
rect 67692 487772 67698 487824
rect 109126 487772 109132 487824
rect 109184 487812 109190 487824
rect 116026 487812 116032 487824
rect 109184 487784 116032 487812
rect 109184 487772 109190 487784
rect 116026 487772 116032 487784
rect 116084 487772 116090 487824
rect 129918 487200 129924 487212
rect 103486 487172 129924 487200
rect 55122 487092 55128 487144
rect 55180 487132 55186 487144
rect 68002 487132 68008 487144
rect 55180 487104 68008 487132
rect 55180 487092 55186 487104
rect 68002 487092 68008 487104
rect 68060 487092 68066 487144
rect 102226 487092 102232 487144
rect 102284 487132 102290 487144
rect 103486 487132 103514 487172
rect 129918 487160 129924 487172
rect 129976 487160 129982 487212
rect 102284 487104 103514 487132
rect 102284 487092 102290 487104
rect 99466 485800 99472 485852
rect 99524 485840 99530 485852
rect 141050 485840 141056 485852
rect 99524 485812 141056 485840
rect 99524 485800 99530 485812
rect 141050 485800 141056 485812
rect 141108 485800 141114 485852
rect 103422 485052 103428 485104
rect 103480 485092 103486 485104
rect 111978 485092 111984 485104
rect 103480 485064 111984 485092
rect 103480 485052 103486 485064
rect 111978 485052 111984 485064
rect 112036 485052 112042 485104
rect 67634 484412 67640 484424
rect 53116 484384 67640 484412
rect 53116 484356 53144 484384
rect 67634 484372 67640 484384
rect 67692 484372 67698 484424
rect 286318 484372 286324 484424
rect 286376 484412 286382 484424
rect 580166 484412 580172 484424
rect 286376 484384 580172 484412
rect 286376 484372 286382 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 50982 484304 50988 484356
rect 51040 484344 51046 484356
rect 53098 484344 53104 484356
rect 51040 484316 53104 484344
rect 51040 484304 51046 484316
rect 53098 484304 53104 484316
rect 53156 484304 53162 484356
rect 36998 483624 37004 483676
rect 37056 483664 37062 483676
rect 65886 483664 65892 483676
rect 37056 483636 65892 483664
rect 37056 483624 37062 483636
rect 65886 483624 65892 483636
rect 65944 483664 65950 483676
rect 67634 483664 67640 483676
rect 65944 483636 67640 483664
rect 65944 483624 65950 483636
rect 67634 483624 67640 483636
rect 67692 483624 67698 483676
rect 103422 483624 103428 483676
rect 103480 483664 103486 483676
rect 122834 483664 122840 483676
rect 103480 483636 122840 483664
rect 103480 483624 103486 483636
rect 122834 483624 122840 483636
rect 122892 483664 122898 483676
rect 123386 483664 123392 483676
rect 122892 483636 123392 483664
rect 122892 483624 122898 483636
rect 123386 483624 123392 483636
rect 123444 483624 123450 483676
rect 39758 482944 39764 482996
rect 39816 482984 39822 482996
rect 68094 482984 68100 482996
rect 39816 482956 68100 482984
rect 39816 482944 39822 482956
rect 68094 482944 68100 482956
rect 68152 482944 68158 482996
rect 115198 482944 115204 482996
rect 115256 482984 115262 482996
rect 117406 482984 117412 482996
rect 115256 482956 117412 482984
rect 115256 482944 115262 482956
rect 117406 482944 117412 482956
rect 117464 482944 117470 482996
rect 67358 482400 67364 482452
rect 67416 482440 67422 482452
rect 69842 482440 69848 482452
rect 67416 482412 69848 482440
rect 67416 482400 67422 482412
rect 69842 482400 69848 482412
rect 69900 482400 69906 482452
rect 36906 482264 36912 482316
rect 36964 482304 36970 482316
rect 66898 482304 66904 482316
rect 36964 482276 66904 482304
rect 36964 482264 36970 482276
rect 66898 482264 66904 482276
rect 66956 482304 66962 482316
rect 67450 482304 67456 482316
rect 66956 482276 67456 482304
rect 66956 482264 66962 482276
rect 67450 482264 67456 482276
rect 67508 482264 67514 482316
rect 103422 482264 103428 482316
rect 103480 482304 103486 482316
rect 114554 482304 114560 482316
rect 103480 482276 114560 482304
rect 103480 482264 103486 482276
rect 114554 482264 114560 482276
rect 114612 482264 114618 482316
rect 106274 481788 106280 481840
rect 106332 481828 106338 481840
rect 107010 481828 107016 481840
rect 106332 481800 107016 481828
rect 106332 481788 106338 481800
rect 107010 481788 107016 481800
rect 107068 481828 107074 481840
rect 107068 481800 113174 481828
rect 107068 481788 107074 481800
rect 103330 481720 103336 481772
rect 103388 481760 103394 481772
rect 110322 481760 110328 481772
rect 103388 481732 110328 481760
rect 103388 481720 103394 481732
rect 110322 481720 110328 481732
rect 110380 481720 110386 481772
rect 113146 481692 113174 481800
rect 129826 481720 129832 481772
rect 129884 481760 129890 481772
rect 130378 481760 130384 481772
rect 129884 481732 130384 481760
rect 129884 481720 129890 481732
rect 130378 481720 130384 481732
rect 130436 481760 130442 481772
rect 143718 481760 143724 481772
rect 130436 481732 143724 481760
rect 130436 481720 130442 481732
rect 143718 481720 143724 481732
rect 143776 481720 143782 481772
rect 146294 481692 146300 481704
rect 113146 481664 146300 481692
rect 146294 481652 146300 481664
rect 146352 481652 146358 481704
rect 52178 481584 52184 481636
rect 52236 481624 52242 481636
rect 69106 481624 69112 481636
rect 52236 481596 69112 481624
rect 52236 481584 52242 481596
rect 69106 481584 69112 481596
rect 69164 481584 69170 481636
rect 103422 481584 103428 481636
rect 103480 481624 103486 481636
rect 129826 481624 129832 481636
rect 103480 481596 129832 481624
rect 103480 481584 103486 481596
rect 129826 481584 129832 481596
rect 129884 481584 129890 481636
rect 103330 481516 103336 481568
rect 103388 481556 103394 481568
rect 106274 481556 106280 481568
rect 103388 481528 106280 481556
rect 103388 481516 103394 481528
rect 106274 481516 106280 481528
rect 106332 481516 106338 481568
rect 110322 481516 110328 481568
rect 110380 481556 110386 481568
rect 124214 481556 124220 481568
rect 110380 481528 124220 481556
rect 110380 481516 110386 481528
rect 124214 481516 124220 481528
rect 124272 481516 124278 481568
rect 54846 480224 54852 480276
rect 54904 480264 54910 480276
rect 57238 480264 57244 480276
rect 54904 480236 57244 480264
rect 54904 480224 54910 480236
rect 57238 480224 57244 480236
rect 57296 480264 57302 480276
rect 57296 480236 57974 480264
rect 57296 480224 57302 480236
rect 57946 480196 57974 480236
rect 67634 480196 67640 480208
rect 57946 480168 67640 480196
rect 67634 480156 67640 480168
rect 67692 480156 67698 480208
rect 103330 479544 103336 479596
rect 103388 479584 103394 479596
rect 107654 479584 107660 479596
rect 103388 479556 107660 479584
rect 103388 479544 103394 479556
rect 107654 479544 107660 479556
rect 107712 479584 107718 479596
rect 115198 479584 115204 479596
rect 107712 479556 115204 479584
rect 107712 479544 107718 479556
rect 115198 479544 115204 479556
rect 115256 479544 115262 479596
rect 103422 479476 103428 479528
rect 103480 479516 103486 479528
rect 133874 479516 133880 479528
rect 103480 479488 133880 479516
rect 103480 479476 103486 479488
rect 133874 479476 133880 479488
rect 133932 479476 133938 479528
rect 64414 478864 64420 478916
rect 64472 478904 64478 478916
rect 65794 478904 65800 478916
rect 64472 478876 65800 478904
rect 64472 478864 64478 478876
rect 65794 478864 65800 478876
rect 65852 478864 65858 478916
rect 105630 478864 105636 478916
rect 105688 478904 105694 478916
rect 109218 478904 109224 478916
rect 105688 478876 109224 478904
rect 105688 478864 105694 478876
rect 109218 478864 109224 478876
rect 109276 478864 109282 478916
rect 128998 478864 129004 478916
rect 129056 478904 129062 478916
rect 129826 478904 129832 478916
rect 129056 478876 129832 478904
rect 129056 478864 129062 478876
rect 129826 478864 129832 478876
rect 129884 478864 129890 478916
rect 60550 478796 60556 478848
rect 60608 478836 60614 478848
rect 67266 478836 67272 478848
rect 60608 478808 67272 478836
rect 60608 478796 60614 478808
rect 67266 478796 67272 478808
rect 67324 478796 67330 478848
rect 103422 477504 103428 477556
rect 103480 477544 103486 477556
rect 103480 477516 109034 477544
rect 103480 477504 103486 477516
rect 109006 477488 109034 477516
rect 108942 477436 108948 477488
rect 109000 477476 109034 477488
rect 142154 477476 142160 477488
rect 109000 477448 142160 477476
rect 109000 477436 109006 477448
rect 142154 477436 142160 477448
rect 142212 477436 142218 477488
rect 103330 476824 103336 476876
rect 103388 476864 103394 476876
rect 125870 476864 125876 476876
rect 103388 476836 125876 476864
rect 103388 476824 103394 476836
rect 125870 476824 125876 476836
rect 125928 476824 125934 476876
rect 105170 476756 105176 476808
rect 105228 476796 105234 476808
rect 129826 476796 129832 476808
rect 105228 476768 129832 476796
rect 105228 476756 105234 476768
rect 129826 476756 129832 476768
rect 129884 476756 129890 476808
rect 34330 476076 34336 476128
rect 34388 476116 34394 476128
rect 67634 476116 67640 476128
rect 34388 476088 67640 476116
rect 34388 476076 34394 476088
rect 67634 476076 67640 476088
rect 67692 476076 67698 476128
rect 117958 476076 117964 476128
rect 118016 476116 118022 476128
rect 124306 476116 124312 476128
rect 118016 476088 124312 476116
rect 118016 476076 118022 476088
rect 124306 476076 124312 476088
rect 124364 476076 124370 476128
rect 103238 476008 103244 476060
rect 103296 476048 103302 476060
rect 120258 476048 120264 476060
rect 103296 476020 120264 476048
rect 103296 476008 103302 476020
rect 120258 476008 120264 476020
rect 120316 476008 120322 476060
rect 102226 475940 102232 475992
rect 102284 475980 102290 475992
rect 117958 475980 117964 475992
rect 102284 475952 117964 475980
rect 102284 475940 102290 475952
rect 117958 475940 117964 475952
rect 118016 475940 118022 475992
rect 102318 475872 102324 475924
rect 102376 475912 102382 475924
rect 111886 475912 111892 475924
rect 102376 475884 111892 475912
rect 102376 475872 102382 475884
rect 111886 475872 111892 475884
rect 111944 475912 111950 475924
rect 112622 475912 112628 475924
rect 111944 475884 112628 475912
rect 111944 475872 111950 475884
rect 112622 475872 112628 475884
rect 112680 475872 112686 475924
rect 59078 475396 59084 475448
rect 59136 475436 59142 475448
rect 67634 475436 67640 475448
rect 59136 475408 67640 475436
rect 59136 475396 59142 475408
rect 67634 475396 67640 475408
rect 67692 475396 67698 475448
rect 35618 475328 35624 475380
rect 35676 475368 35682 475380
rect 65978 475368 65984 475380
rect 35676 475340 65984 475368
rect 35676 475328 35682 475340
rect 65978 475328 65984 475340
rect 66036 475368 66042 475380
rect 67726 475368 67732 475380
rect 66036 475340 67732 475368
rect 66036 475328 66042 475340
rect 67726 475328 67732 475340
rect 67784 475328 67790 475380
rect 112622 475328 112628 475380
rect 112680 475368 112686 475380
rect 122834 475368 122840 475380
rect 112680 475340 122840 475368
rect 112680 475328 112686 475340
rect 122834 475328 122840 475340
rect 122892 475328 122898 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 11698 474756 11704 474768
rect 3476 474728 11704 474756
rect 3476 474716 3482 474728
rect 11698 474716 11704 474728
rect 11756 474716 11762 474768
rect 102226 474648 102232 474700
rect 102284 474688 102290 474700
rect 113174 474688 113180 474700
rect 102284 474660 113180 474688
rect 102284 474648 102290 474660
rect 113174 474648 113180 474660
rect 113232 474688 113238 474700
rect 115474 474688 115480 474700
rect 113232 474660 115480 474688
rect 113232 474648 113238 474660
rect 115474 474648 115480 474660
rect 115532 474648 115538 474700
rect 61838 474308 61844 474360
rect 61896 474348 61902 474360
rect 65978 474348 65984 474360
rect 61896 474320 65984 474348
rect 61896 474308 61902 474320
rect 65978 474308 65984 474320
rect 66036 474348 66042 474360
rect 67634 474348 67640 474360
rect 66036 474320 67640 474348
rect 66036 474308 66042 474320
rect 67634 474308 67640 474320
rect 67692 474308 67698 474360
rect 42610 473356 42616 473408
rect 42668 473396 42674 473408
rect 53834 473396 53840 473408
rect 42668 473368 53840 473396
rect 42668 473356 42674 473368
rect 53834 473356 53840 473368
rect 53892 473356 53898 473408
rect 64690 473288 64696 473340
rect 64748 473328 64754 473340
rect 67634 473328 67640 473340
rect 64748 473300 67640 473328
rect 64748 473288 64754 473300
rect 67634 473288 67640 473300
rect 67692 473288 67698 473340
rect 102226 473288 102232 473340
rect 102284 473328 102290 473340
rect 133138 473328 133144 473340
rect 102284 473300 133144 473328
rect 102284 473288 102290 473300
rect 133138 473288 133144 473300
rect 133196 473328 133202 473340
rect 133782 473328 133788 473340
rect 133196 473300 133788 473328
rect 133196 473288 133202 473300
rect 133782 473288 133788 473300
rect 133840 473288 133846 473340
rect 52178 472608 52184 472660
rect 52236 472648 52242 472660
rect 64690 472648 64696 472660
rect 52236 472620 64696 472648
rect 52236 472608 52242 472620
rect 64690 472608 64696 472620
rect 64748 472608 64754 472660
rect 102226 472608 102232 472660
rect 102284 472648 102290 472660
rect 123202 472648 123208 472660
rect 102284 472620 123208 472648
rect 102284 472608 102290 472620
rect 123202 472608 123208 472620
rect 123260 472648 123266 472660
rect 124122 472648 124128 472660
rect 123260 472620 124128 472648
rect 123260 472608 123266 472620
rect 124122 472608 124128 472620
rect 124180 472608 124186 472660
rect 133782 472608 133788 472660
rect 133840 472648 133846 472660
rect 142154 472648 142160 472660
rect 133840 472620 142160 472648
rect 133840 472608 133846 472620
rect 142154 472608 142160 472620
rect 142212 472608 142218 472660
rect 102318 471996 102324 472048
rect 102376 472036 102382 472048
rect 103422 472036 103428 472048
rect 102376 472008 103428 472036
rect 102376 471996 102382 472008
rect 103422 471996 103428 472008
rect 103480 472036 103486 472048
rect 146386 472036 146392 472048
rect 103480 472008 146392 472036
rect 103480 471996 103486 472008
rect 146386 471996 146392 472008
rect 146444 471996 146450 472048
rect 124122 471248 124128 471300
rect 124180 471288 124186 471300
rect 145006 471288 145012 471300
rect 124180 471260 145012 471288
rect 124180 471248 124186 471260
rect 145006 471248 145012 471260
rect 145064 471248 145070 471300
rect 61378 470608 61384 470620
rect 60706 470580 61384 470608
rect 41322 470500 41328 470552
rect 41380 470540 41386 470552
rect 60706 470540 60734 470580
rect 61378 470568 61384 470580
rect 61436 470608 61442 470620
rect 67634 470608 67640 470620
rect 61436 470580 67640 470608
rect 61436 470568 61442 470580
rect 67634 470568 67640 470580
rect 67692 470568 67698 470620
rect 102226 470568 102232 470620
rect 102284 470608 102290 470620
rect 102284 470580 106274 470608
rect 102284 470568 102290 470580
rect 41380 470512 60734 470540
rect 41380 470500 41386 470512
rect 64598 470500 64604 470552
rect 64656 470540 64662 470552
rect 65978 470540 65984 470552
rect 64656 470512 65984 470540
rect 64656 470500 64662 470512
rect 65978 470500 65984 470512
rect 66036 470540 66042 470552
rect 67726 470540 67732 470552
rect 66036 470512 67732 470540
rect 66036 470500 66042 470512
rect 67726 470500 67732 470512
rect 67784 470500 67790 470552
rect 106246 470540 106274 470580
rect 145006 470568 145012 470620
rect 145064 470608 145070 470620
rect 579982 470608 579988 470620
rect 145064 470580 579988 470608
rect 145064 470568 145070 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 138014 470540 138020 470552
rect 106246 470512 138020 470540
rect 138014 470500 138020 470512
rect 138072 470500 138078 470552
rect 102226 469888 102232 469940
rect 102284 469928 102290 469940
rect 105538 469928 105544 469940
rect 102284 469900 105544 469928
rect 102284 469888 102290 469900
rect 105538 469888 105544 469900
rect 105596 469928 105602 469940
rect 140958 469928 140964 469940
rect 105596 469900 140964 469928
rect 105596 469888 105602 469900
rect 140958 469888 140964 469900
rect 141016 469888 141022 469940
rect 103606 469820 103612 469872
rect 103664 469860 103670 469872
rect 140774 469860 140780 469872
rect 103664 469832 140780 469860
rect 103664 469820 103670 469832
rect 140774 469820 140780 469832
rect 140832 469860 140838 469872
rect 147858 469860 147864 469872
rect 140832 469832 147864 469860
rect 140832 469820 140838 469832
rect 147858 469820 147864 469832
rect 147916 469820 147922 469872
rect 61746 469548 61752 469600
rect 61804 469588 61810 469600
rect 67634 469588 67640 469600
rect 61804 469560 67640 469588
rect 61804 469548 61810 469560
rect 67634 469548 67640 469560
rect 67692 469548 67698 469600
rect 102226 469208 102232 469260
rect 102284 469248 102290 469260
rect 102284 469220 106274 469248
rect 102284 469208 102290 469220
rect 106246 469192 106274 469220
rect 138014 469208 138020 469260
rect 138072 469248 138078 469260
rect 138198 469248 138204 469260
rect 138072 469220 138204 469248
rect 138072 469208 138078 469220
rect 138198 469208 138204 469220
rect 138256 469208 138262 469260
rect 106182 469180 106188 469192
rect 106141 469152 106188 469180
rect 106182 469140 106188 469152
rect 106240 469180 106274 469192
rect 116118 469180 116124 469192
rect 106240 469152 116124 469180
rect 106240 469140 106246 469152
rect 116118 469140 116124 469152
rect 116176 469140 116182 469192
rect 103606 468460 103612 468512
rect 103664 468500 103670 468512
rect 135438 468500 135444 468512
rect 103664 468472 135444 468500
rect 103664 468460 103670 468472
rect 135438 468460 135444 468472
rect 135496 468500 135502 468512
rect 149146 468500 149152 468512
rect 135496 468472 149152 468500
rect 135496 468460 135502 468472
rect 149146 468460 149152 468472
rect 149204 468460 149210 468512
rect 56318 468324 56324 468376
rect 56376 468364 56382 468376
rect 64138 468364 64144 468376
rect 56376 468336 64144 468364
rect 56376 468324 56382 468336
rect 64138 468324 64144 468336
rect 64196 468324 64202 468376
rect 59262 467848 59268 467900
rect 59320 467888 59326 467900
rect 63218 467888 63224 467900
rect 59320 467860 63224 467888
rect 59320 467848 59326 467860
rect 63218 467848 63224 467860
rect 63276 467888 63282 467900
rect 67634 467888 67640 467900
rect 63276 467860 67640 467888
rect 63276 467848 63282 467860
rect 67634 467848 67640 467860
rect 67692 467848 67698 467900
rect 64782 467780 64788 467832
rect 64840 467820 64846 467832
rect 67450 467820 67456 467832
rect 64840 467792 67456 467820
rect 64840 467780 64846 467792
rect 67450 467780 67456 467792
rect 67508 467780 67514 467832
rect 104158 467100 104164 467152
rect 104216 467140 104222 467152
rect 114830 467140 114836 467152
rect 104216 467112 114836 467140
rect 104216 467100 104222 467112
rect 114830 467100 114836 467112
rect 114888 467100 114894 467152
rect 102226 466488 102232 466540
rect 102284 466528 102290 466540
rect 133782 466528 133788 466540
rect 102284 466500 133788 466528
rect 102284 466488 102290 466500
rect 133782 466488 133788 466500
rect 133840 466488 133846 466540
rect 144914 466460 144920 466472
rect 108316 466432 144920 466460
rect 108316 466404 108344 466432
rect 144914 466420 144920 466432
rect 144972 466420 144978 466472
rect 102318 466352 102324 466404
rect 102376 466392 102382 466404
rect 108298 466392 108304 466404
rect 102376 466364 108304 466392
rect 102376 466352 102382 466364
rect 108298 466352 108304 466364
rect 108356 466352 108362 466404
rect 133782 466352 133788 466404
rect 133840 466392 133846 466404
rect 136634 466392 136640 466404
rect 133840 466364 136640 466392
rect 133840 466352 133846 466364
rect 136634 466352 136640 466364
rect 136692 466352 136698 466404
rect 41046 465672 41052 465724
rect 41104 465712 41110 465724
rect 67634 465712 67640 465724
rect 41104 465684 67640 465712
rect 41104 465672 41110 465684
rect 67634 465672 67640 465684
rect 67692 465672 67698 465724
rect 102226 465672 102232 465724
rect 102284 465712 102290 465724
rect 115934 465712 115940 465724
rect 102284 465684 115940 465712
rect 102284 465672 102290 465684
rect 115934 465672 115940 465684
rect 115992 465712 115998 465724
rect 116854 465712 116860 465724
rect 115992 465684 116860 465712
rect 115992 465672 115998 465684
rect 116854 465672 116860 465684
rect 116912 465672 116918 465724
rect 66070 465332 66076 465384
rect 66128 465372 66134 465384
rect 67542 465372 67548 465384
rect 66128 465344 67548 465372
rect 66128 465332 66134 465344
rect 67542 465332 67548 465344
rect 67600 465372 67606 465384
rect 67910 465372 67916 465384
rect 67600 465344 67916 465372
rect 67600 465332 67606 465344
rect 67910 465332 67916 465344
rect 67968 465332 67974 465384
rect 113910 465100 113916 465112
rect 113146 465072 113916 465100
rect 102226 464992 102232 465044
rect 102284 465032 102290 465044
rect 113146 465032 113174 465072
rect 113910 465060 113916 465072
rect 113968 465100 113974 465112
rect 150618 465100 150624 465112
rect 113968 465072 150624 465100
rect 113968 465060 113974 465072
rect 150618 465060 150624 465072
rect 150676 465060 150682 465112
rect 102284 465004 113174 465032
rect 102284 464992 102290 465004
rect 116854 464992 116860 465044
rect 116912 465032 116918 465044
rect 121638 465032 121644 465044
rect 116912 465004 121644 465032
rect 116912 464992 116918 465004
rect 121638 464992 121644 465004
rect 121696 464992 121702 465044
rect 49418 464312 49424 464364
rect 49476 464352 49482 464364
rect 67634 464352 67640 464364
rect 49476 464324 67640 464352
rect 49476 464312 49482 464324
rect 67634 464312 67640 464324
rect 67692 464312 67698 464364
rect 108298 464312 108304 464364
rect 108356 464352 108362 464364
rect 110782 464352 110788 464364
rect 108356 464324 110788 464352
rect 108356 464312 108362 464324
rect 110782 464312 110788 464324
rect 110840 464312 110846 464364
rect 128630 463740 128636 463752
rect 117240 463712 128636 463740
rect 49418 463632 49424 463684
rect 49476 463672 49482 463684
rect 50338 463672 50344 463684
rect 49476 463644 50344 463672
rect 49476 463632 49482 463644
rect 50338 463632 50344 463644
rect 50396 463632 50402 463684
rect 102226 463632 102232 463684
rect 102284 463672 102290 463684
rect 116578 463672 116584 463684
rect 102284 463644 116584 463672
rect 102284 463632 102290 463644
rect 116578 463632 116584 463644
rect 116636 463672 116642 463684
rect 117240 463672 117268 463712
rect 128630 463700 128636 463712
rect 128688 463700 128694 463752
rect 116636 463644 117268 463672
rect 116636 463632 116642 463644
rect 56502 462952 56508 463004
rect 56560 462992 56566 463004
rect 67634 462992 67640 463004
rect 56560 462964 67640 462992
rect 56560 462952 56566 462964
rect 67634 462952 67640 462964
rect 67692 462952 67698 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 102226 462272 102232 462324
rect 102284 462312 102290 462324
rect 140774 462312 140780 462324
rect 102284 462284 140780 462312
rect 102284 462272 102290 462284
rect 140774 462272 140780 462284
rect 140832 462272 140838 462324
rect 60458 461592 60464 461644
rect 60516 461632 60522 461644
rect 67634 461632 67640 461644
rect 60516 461604 67640 461632
rect 60516 461592 60522 461604
rect 67634 461592 67640 461604
rect 67692 461592 67698 461644
rect 102318 460980 102324 461032
rect 102376 461020 102382 461032
rect 115934 461020 115940 461032
rect 102376 460992 115940 461020
rect 102376 460980 102382 460992
rect 115934 460980 115940 460992
rect 115992 460980 115998 461032
rect 147766 460952 147772 460964
rect 108960 460924 147772 460952
rect 102226 460844 102232 460896
rect 102284 460884 102290 460896
rect 108390 460884 108396 460896
rect 102284 460856 108396 460884
rect 102284 460844 102290 460856
rect 108390 460844 108396 460856
rect 108448 460884 108454 460896
rect 108960 460884 108988 460924
rect 147766 460912 147772 460924
rect 147824 460912 147830 460964
rect 108448 460856 108988 460884
rect 108448 460844 108454 460856
rect 115934 460844 115940 460896
rect 115992 460884 115998 460896
rect 118970 460884 118976 460896
rect 115992 460856 118976 460884
rect 115992 460844 115998 460856
rect 118970 460844 118976 460856
rect 119028 460844 119034 460896
rect 108390 460232 108396 460284
rect 108448 460272 108454 460284
rect 124582 460272 124588 460284
rect 108448 460244 124588 460272
rect 108448 460232 108454 460244
rect 124582 460232 124588 460244
rect 124640 460232 124646 460284
rect 42702 460164 42708 460216
rect 42760 460204 42766 460216
rect 52454 460204 52460 460216
rect 42760 460176 52460 460204
rect 42760 460164 42766 460176
rect 52454 460164 52460 460176
rect 52512 460164 52518 460216
rect 57790 460164 57796 460216
rect 57848 460204 57854 460216
rect 67634 460204 67640 460216
rect 57848 460176 67640 460204
rect 57848 460164 57854 460176
rect 67634 460164 67640 460176
rect 67692 460164 67698 460216
rect 102318 460164 102324 460216
rect 102376 460204 102382 460216
rect 138106 460204 138112 460216
rect 102376 460176 138112 460204
rect 102376 460164 102382 460176
rect 138106 460164 138112 460176
rect 138164 460204 138170 460216
rect 151906 460204 151912 460216
rect 138164 460176 151912 460204
rect 138164 460164 138170 460176
rect 151906 460164 151912 460176
rect 151964 460164 151970 460216
rect 52454 459552 52460 459604
rect 52512 459592 52518 459604
rect 53650 459592 53656 459604
rect 52512 459564 53656 459592
rect 52512 459552 52518 459564
rect 53650 459552 53656 459564
rect 53708 459592 53714 459604
rect 67634 459592 67640 459604
rect 53708 459564 67640 459592
rect 53708 459552 53714 459564
rect 67634 459552 67640 459564
rect 67692 459552 67698 459604
rect 102410 459552 102416 459604
rect 102468 459592 102474 459604
rect 108390 459592 108396 459604
rect 102468 459564 108396 459592
rect 102468 459552 102474 459564
rect 108390 459552 108396 459564
rect 108448 459592 108454 459604
rect 108850 459592 108856 459604
rect 108448 459564 108856 459592
rect 108448 459552 108454 459564
rect 108850 459552 108856 459564
rect 108908 459552 108914 459604
rect 125134 459552 125140 459604
rect 125192 459592 125198 459604
rect 128354 459592 128360 459604
rect 125192 459564 128360 459592
rect 125192 459552 125198 459564
rect 128354 459552 128360 459564
rect 128412 459552 128418 459604
rect 66162 459484 66168 459536
rect 66220 459524 66226 459536
rect 67726 459524 67732 459536
rect 66220 459496 67732 459524
rect 66220 459484 66226 459496
rect 67726 459484 67732 459496
rect 67784 459484 67790 459536
rect 43990 458872 43996 458924
rect 44048 458912 44054 458924
rect 57790 458912 57796 458924
rect 44048 458884 57796 458912
rect 44048 458872 44054 458884
rect 57790 458872 57796 458884
rect 57848 458872 57854 458924
rect 64138 458872 64144 458924
rect 64196 458912 64202 458924
rect 64782 458912 64788 458924
rect 64196 458884 64788 458912
rect 64196 458872 64202 458884
rect 64782 458872 64788 458884
rect 64840 458912 64846 458924
rect 67634 458912 67640 458924
rect 64840 458884 67640 458912
rect 64840 458872 64846 458884
rect 67634 458872 67640 458884
rect 67692 458872 67698 458924
rect 102226 458872 102232 458924
rect 102284 458912 102290 458924
rect 124214 458912 124220 458924
rect 102284 458884 124220 458912
rect 102284 458872 102290 458884
rect 124214 458872 124220 458884
rect 124272 458912 124278 458924
rect 125134 458912 125140 458924
rect 124272 458884 125140 458912
rect 124272 458872 124278 458884
rect 125134 458872 125140 458884
rect 125192 458872 125198 458924
rect 45462 458804 45468 458856
rect 45520 458844 45526 458856
rect 66162 458844 66168 458856
rect 45520 458816 66168 458844
rect 45520 458804 45526 458816
rect 66162 458804 66168 458816
rect 66220 458804 66226 458856
rect 103606 458804 103612 458856
rect 103664 458844 103670 458856
rect 142246 458844 142252 458856
rect 103664 458816 142252 458844
rect 103664 458804 103670 458816
rect 142246 458804 142252 458816
rect 142304 458844 142310 458856
rect 151998 458844 152004 458856
rect 142304 458816 152004 458844
rect 142304 458804 142310 458816
rect 151998 458804 152004 458816
rect 152056 458804 152062 458856
rect 108482 458192 108488 458244
rect 108540 458232 108546 458244
rect 138106 458232 138112 458244
rect 108540 458204 138112 458232
rect 108540 458192 108546 458204
rect 138106 458192 138112 458204
rect 138164 458192 138170 458244
rect 39758 458124 39764 458176
rect 39816 458164 39822 458176
rect 43714 458164 43720 458176
rect 39816 458136 43720 458164
rect 39816 458124 39822 458136
rect 43714 458124 43720 458136
rect 43772 458164 43778 458176
rect 67726 458164 67732 458176
rect 43772 458136 67732 458164
rect 43772 458124 43778 458136
rect 67726 458124 67732 458136
rect 67784 458124 67790 458176
rect 36998 457444 37004 457496
rect 37056 457484 37062 457496
rect 67634 457484 67640 457496
rect 37056 457456 67640 457484
rect 37056 457444 37062 457456
rect 67634 457444 67640 457456
rect 67692 457444 67698 457496
rect 143626 456804 143632 456816
rect 107580 456776 143632 456804
rect 102226 456696 102232 456748
rect 102284 456736 102290 456748
rect 106918 456736 106924 456748
rect 102284 456708 106924 456736
rect 102284 456696 102290 456708
rect 106918 456696 106924 456708
rect 106976 456736 106982 456748
rect 107580 456736 107608 456776
rect 143626 456764 143632 456776
rect 143684 456764 143690 456816
rect 446398 456764 446404 456816
rect 446456 456804 446462 456816
rect 580166 456804 580172 456816
rect 446456 456776 580172 456804
rect 446456 456764 446462 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 106976 456708 107608 456736
rect 106976 456696 106982 456708
rect 100202 456152 100208 456204
rect 100260 456192 100266 456204
rect 109310 456192 109316 456204
rect 100260 456164 109316 456192
rect 100260 456152 100266 456164
rect 109310 456152 109316 456164
rect 109368 456152 109374 456204
rect 102318 456084 102324 456136
rect 102376 456124 102382 456136
rect 132494 456124 132500 456136
rect 102376 456096 132500 456124
rect 102376 456084 102382 456096
rect 132494 456084 132500 456096
rect 132552 456084 132558 456136
rect 106090 456016 106096 456068
rect 106148 456056 106154 456068
rect 135254 456056 135260 456068
rect 106148 456028 135260 456056
rect 106148 456016 106154 456028
rect 135254 456016 135260 456028
rect 135312 456056 135318 456068
rect 142246 456056 142252 456068
rect 135312 456028 142252 456056
rect 135312 456016 135318 456028
rect 142246 456016 142252 456028
rect 142304 456016 142310 456068
rect 67634 455444 67640 455456
rect 64800 455416 67640 455444
rect 37182 455336 37188 455388
rect 37240 455376 37246 455388
rect 64138 455376 64144 455388
rect 37240 455348 64144 455376
rect 37240 455336 37246 455348
rect 64138 455336 64144 455348
rect 64196 455376 64202 455388
rect 64800 455376 64828 455416
rect 67634 455404 67640 455416
rect 67692 455404 67698 455456
rect 64196 455348 64828 455376
rect 64196 455336 64202 455348
rect 102318 455336 102324 455388
rect 102376 455376 102382 455388
rect 108482 455376 108488 455388
rect 102376 455348 108488 455376
rect 102376 455336 102382 455348
rect 108482 455336 108488 455348
rect 108540 455336 108546 455388
rect 55030 455268 55036 455320
rect 55088 455308 55094 455320
rect 57330 455308 57336 455320
rect 55088 455280 57336 455308
rect 55088 455268 55094 455280
rect 57330 455268 57336 455280
rect 57388 455268 57394 455320
rect 102226 455268 102232 455320
rect 102284 455308 102290 455320
rect 106090 455308 106096 455320
rect 102284 455280 106096 455308
rect 102284 455268 102290 455280
rect 106090 455268 106096 455280
rect 106148 455268 106154 455320
rect 107378 454656 107384 454708
rect 107436 454696 107442 454708
rect 139486 454696 139492 454708
rect 107436 454668 139492 454696
rect 107436 454656 107442 454668
rect 139486 454656 139492 454668
rect 139544 454696 139550 454708
rect 150526 454696 150532 454708
rect 139544 454668 150532 454696
rect 139544 454656 139550 454668
rect 150526 454656 150532 454668
rect 150584 454656 150590 454708
rect 57330 454044 57336 454096
rect 57388 454084 57394 454096
rect 67634 454084 67640 454096
rect 57388 454056 67640 454084
rect 57388 454044 57394 454056
rect 67634 454044 67640 454056
rect 67692 454044 67698 454096
rect 102226 453976 102232 454028
rect 102284 454016 102290 454028
rect 125778 454016 125784 454028
rect 102284 453988 125784 454016
rect 102284 453976 102290 453988
rect 125778 453976 125784 453988
rect 125836 453976 125842 454028
rect 102318 453908 102324 453960
rect 102376 453948 102382 453960
rect 107378 453948 107384 453960
rect 102376 453920 107384 453948
rect 102376 453908 102382 453920
rect 107378 453908 107384 453920
rect 107436 453908 107442 453960
rect 53742 452684 53748 452736
rect 53800 452724 53806 452736
rect 57790 452724 57796 452736
rect 53800 452696 57796 452724
rect 53800 452684 53806 452696
rect 57790 452684 57796 452696
rect 57848 452724 57854 452736
rect 67634 452724 67640 452736
rect 57848 452696 67640 452724
rect 57848 452684 57854 452696
rect 67634 452684 67640 452696
rect 67692 452684 67698 452736
rect 67726 452656 67732 452668
rect 51736 452628 67732 452656
rect 51736 452600 51764 452628
rect 67726 452616 67732 452628
rect 67784 452616 67790 452668
rect 50890 452548 50896 452600
rect 50948 452588 50954 452600
rect 51718 452588 51724 452600
rect 50948 452560 51724 452588
rect 50948 452548 50954 452560
rect 51718 452548 51724 452560
rect 51776 452548 51782 452600
rect 102226 452548 102232 452600
rect 102284 452588 102290 452600
rect 133966 452588 133972 452600
rect 102284 452560 133972 452588
rect 102284 452548 102290 452560
rect 133966 452548 133972 452560
rect 134024 452588 134030 452600
rect 135162 452588 135168 452600
rect 134024 452560 135168 452588
rect 134024 452548 134030 452560
rect 135162 452548 135168 452560
rect 135220 452548 135226 452600
rect 136726 452480 136732 452532
rect 136784 452520 136790 452532
rect 137370 452520 137376 452532
rect 136784 452492 137376 452520
rect 136784 452480 136790 452492
rect 137370 452480 137376 452492
rect 137428 452480 137434 452532
rect 135162 451868 135168 451920
rect 135220 451908 135226 451920
rect 147674 451908 147680 451920
rect 135220 451880 147680 451908
rect 135220 451868 135226 451880
rect 147674 451868 147680 451880
rect 147732 451868 147738 451920
rect 62482 451460 62488 451512
rect 62540 451500 62546 451512
rect 67634 451500 67640 451512
rect 62540 451472 67640 451500
rect 62540 451460 62546 451472
rect 67634 451460 67640 451472
rect 67692 451460 67698 451512
rect 102778 451256 102784 451308
rect 102836 451296 102842 451308
rect 137370 451296 137376 451308
rect 102836 451268 137376 451296
rect 102836 451256 102842 451268
rect 137370 451256 137376 451268
rect 137428 451256 137434 451308
rect 35710 451188 35716 451240
rect 35768 451228 35774 451240
rect 67634 451228 67640 451240
rect 35768 451200 67640 451228
rect 35768 451188 35774 451200
rect 67634 451188 67640 451200
rect 67692 451188 67698 451240
rect 38562 451120 38568 451172
rect 38620 451160 38626 451172
rect 62482 451160 62488 451172
rect 38620 451132 62488 451160
rect 38620 451120 38626 451132
rect 62482 451120 62488 451132
rect 62540 451120 62546 451172
rect 102226 450236 102232 450288
rect 102284 450276 102290 450288
rect 104986 450276 104992 450288
rect 102284 450248 104992 450276
rect 102284 450236 102290 450248
rect 104986 450236 104992 450248
rect 105044 450276 105050 450288
rect 105906 450276 105912 450288
rect 105044 450248 105912 450276
rect 105044 450236 105050 450248
rect 105906 450236 105912 450248
rect 105964 450236 105970 450288
rect 33042 449896 33048 449948
rect 33100 449936 33106 449948
rect 35710 449936 35716 449948
rect 33100 449908 35716 449936
rect 33100 449896 33106 449908
rect 35710 449896 35716 449908
rect 35768 449896 35774 449948
rect 102226 448672 102232 448724
rect 102284 448712 102290 448724
rect 106826 448712 106832 448724
rect 102284 448684 106832 448712
rect 102284 448672 102290 448684
rect 106826 448672 106832 448684
rect 106884 448672 106890 448724
rect 107378 448604 107384 448656
rect 107436 448644 107442 448656
rect 119338 448644 119344 448656
rect 107436 448616 119344 448644
rect 107436 448604 107442 448616
rect 119338 448604 119344 448616
rect 119396 448604 119402 448656
rect 60458 448536 60464 448588
rect 60516 448576 60522 448588
rect 61746 448576 61752 448588
rect 60516 448548 61752 448576
rect 60516 448536 60522 448548
rect 61746 448536 61752 448548
rect 61804 448536 61810 448588
rect 131114 448576 131120 448588
rect 106200 448548 131120 448576
rect 39850 448468 39856 448520
rect 39908 448508 39914 448520
rect 67818 448508 67824 448520
rect 39908 448480 67824 448508
rect 39908 448468 39914 448480
rect 67818 448468 67824 448480
rect 67876 448468 67882 448520
rect 102226 448468 102232 448520
rect 102284 448508 102290 448520
rect 106200 448508 106228 448548
rect 131114 448536 131120 448548
rect 131172 448536 131178 448588
rect 102284 448480 106228 448508
rect 102284 448468 102290 448480
rect 139486 448468 139492 448520
rect 139544 448508 139550 448520
rect 140682 448508 140688 448520
rect 139544 448480 140688 448508
rect 139544 448468 139550 448480
rect 140682 448468 140688 448480
rect 140740 448508 140746 448520
rect 142338 448508 142344 448520
rect 140740 448480 142344 448508
rect 140740 448468 140746 448480
rect 142338 448468 142344 448480
rect 142396 448468 142402 448520
rect 61930 448400 61936 448452
rect 61988 448440 61994 448452
rect 62114 448440 62120 448452
rect 61988 448412 62120 448440
rect 61988 448400 61994 448412
rect 62114 448400 62120 448412
rect 62172 448400 62178 448452
rect 102318 448400 102324 448452
rect 102376 448440 102382 448452
rect 107378 448440 107384 448452
rect 102376 448412 107384 448440
rect 102376 448400 102382 448412
rect 107378 448400 107384 448412
rect 107436 448400 107442 448452
rect 106826 447788 106832 447840
rect 106884 447828 106890 447840
rect 139486 447828 139492 447840
rect 106884 447800 139492 447828
rect 106884 447788 106890 447800
rect 139486 447788 139492 447800
rect 139544 447788 139550 447840
rect 62114 447176 62120 447228
rect 62172 447216 62178 447228
rect 67634 447216 67640 447228
rect 62172 447188 67640 447216
rect 62172 447176 62178 447188
rect 67634 447176 67640 447188
rect 67692 447176 67698 447228
rect 104710 447108 104716 447160
rect 104768 447148 104774 447160
rect 110598 447148 110604 447160
rect 104768 447120 110604 447148
rect 104768 447108 104774 447120
rect 110598 447108 110604 447120
rect 110656 447108 110662 447160
rect 60734 445816 60740 445868
rect 60792 445856 60798 445868
rect 61930 445856 61936 445868
rect 60792 445828 61936 445856
rect 60792 445816 60798 445828
rect 61930 445816 61936 445828
rect 61988 445856 61994 445868
rect 67726 445856 67732 445868
rect 61988 445828 67732 445856
rect 61988 445816 61994 445828
rect 67726 445816 67732 445828
rect 67784 445816 67790 445868
rect 102042 445816 102048 445868
rect 102100 445856 102106 445868
rect 102410 445856 102416 445868
rect 102100 445828 102416 445856
rect 102100 445816 102106 445828
rect 102410 445816 102416 445828
rect 102468 445856 102474 445868
rect 135254 445856 135260 445868
rect 102468 445828 135260 445856
rect 102468 445816 102474 445828
rect 135254 445816 135260 445828
rect 135312 445816 135318 445868
rect 65518 445788 65524 445800
rect 65076 445760 65524 445788
rect 35802 445680 35808 445732
rect 35860 445720 35866 445732
rect 65076 445720 65104 445760
rect 65518 445748 65524 445760
rect 65576 445788 65582 445800
rect 67634 445788 67640 445800
rect 65576 445760 67640 445788
rect 65576 445748 65582 445760
rect 67634 445748 67640 445760
rect 67692 445748 67698 445800
rect 102318 445748 102324 445800
rect 102376 445788 102382 445800
rect 143534 445788 143540 445800
rect 102376 445760 143540 445788
rect 102376 445748 102382 445760
rect 143534 445748 143540 445760
rect 143592 445748 143598 445800
rect 35860 445692 65104 445720
rect 35860 445680 35866 445692
rect 102226 445680 102232 445732
rect 102284 445720 102290 445732
rect 104894 445720 104900 445732
rect 102284 445692 104900 445720
rect 102284 445680 102290 445692
rect 104894 445680 104900 445692
rect 104952 445720 104958 445732
rect 105538 445720 105544 445732
rect 104952 445692 105544 445720
rect 104952 445680 104958 445692
rect 105538 445680 105544 445692
rect 105596 445680 105602 445732
rect 127618 444456 127624 444508
rect 127676 444496 127682 444508
rect 140866 444496 140872 444508
rect 127676 444468 140872 444496
rect 127676 444456 127682 444468
rect 140866 444456 140872 444468
rect 140924 444456 140930 444508
rect 104802 444388 104808 444440
rect 104860 444428 104866 444440
rect 129734 444428 129740 444440
rect 104860 444400 129740 444428
rect 104860 444388 104866 444400
rect 129734 444388 129740 444400
rect 129792 444388 129798 444440
rect 102226 443980 102232 444032
rect 102284 444020 102290 444032
rect 104802 444020 104808 444032
rect 102284 443992 104808 444020
rect 102284 443980 102290 443992
rect 104802 443980 104808 443992
rect 104860 443980 104866 444032
rect 46842 443640 46848 443692
rect 46900 443680 46906 443692
rect 67634 443680 67640 443692
rect 46900 443652 67640 443680
rect 46900 443640 46906 443652
rect 67634 443640 67640 443652
rect 67692 443640 67698 443692
rect 62758 442416 62764 442468
rect 62816 442456 62822 442468
rect 63402 442456 63408 442468
rect 62816 442428 63408 442456
rect 62816 442416 62822 442428
rect 63402 442416 63408 442428
rect 63460 442456 63466 442468
rect 67634 442456 67640 442468
rect 63460 442428 67640 442456
rect 63460 442416 63466 442428
rect 67634 442416 67640 442428
rect 67692 442416 67698 442468
rect 34238 442212 34244 442264
rect 34296 442252 34302 442264
rect 67634 442252 67640 442264
rect 34296 442224 67640 442252
rect 34296 442212 34302 442224
rect 67634 442212 67640 442224
rect 67692 442212 67698 442264
rect 102226 442212 102232 442264
rect 102284 442252 102290 442264
rect 108298 442252 108304 442264
rect 102284 442224 108304 442252
rect 102284 442212 102290 442224
rect 108298 442212 108304 442224
rect 108356 442212 108362 442264
rect 62022 441532 62028 441584
rect 62080 441572 62086 441584
rect 64506 441572 64512 441584
rect 62080 441544 64512 441572
rect 62080 441532 62086 441544
rect 64506 441532 64512 441544
rect 64564 441532 64570 441584
rect 102226 441532 102232 441584
rect 102284 441572 102290 441584
rect 132586 441572 132592 441584
rect 102284 441544 132592 441572
rect 102284 441532 102290 441544
rect 132586 441532 132592 441544
rect 132644 441532 132650 441584
rect 61746 441464 61752 441516
rect 61804 441504 61810 441516
rect 63310 441504 63316 441516
rect 61804 441476 63316 441504
rect 61804 441464 61810 441476
rect 63310 441464 63316 441476
rect 63368 441504 63374 441516
rect 67634 441504 67640 441516
rect 63368 441476 67640 441504
rect 63368 441464 63374 441476
rect 67634 441464 67640 441476
rect 67692 441464 67698 441516
rect 64506 440920 64512 440972
rect 64564 440960 64570 440972
rect 67634 440960 67640 440972
rect 64564 440932 67640 440960
rect 64564 440920 64570 440932
rect 67634 440920 67640 440932
rect 67692 440920 67698 440972
rect 112162 440960 112168 440972
rect 99346 440932 112168 440960
rect 38470 440852 38476 440904
rect 38528 440892 38534 440904
rect 38528 440864 60734 440892
rect 38528 440852 38534 440864
rect 60706 440688 60734 440864
rect 71038 440688 71044 440700
rect 60706 440660 71044 440688
rect 71038 440648 71044 440660
rect 71096 440648 71102 440700
rect 94130 440648 94136 440700
rect 94188 440688 94194 440700
rect 99346 440688 99374 440932
rect 112162 440920 112168 440932
rect 112220 440920 112226 440972
rect 94188 440660 99374 440688
rect 94188 440648 94194 440660
rect 91738 440580 91744 440632
rect 91796 440620 91802 440632
rect 111794 440620 111800 440632
rect 91796 440592 111800 440620
rect 91796 440580 91802 440592
rect 111794 440580 111800 440592
rect 111852 440580 111858 440632
rect 132586 440308 132592 440360
rect 132644 440348 132650 440360
rect 133966 440348 133972 440360
rect 132644 440320 133972 440348
rect 132644 440308 132650 440320
rect 133966 440308 133972 440320
rect 134024 440308 134030 440360
rect 37090 440240 37096 440292
rect 37148 440280 37154 440292
rect 38470 440280 38476 440292
rect 37148 440252 38476 440280
rect 37148 440240 37154 440252
rect 38470 440240 38476 440252
rect 38528 440240 38534 440292
rect 100662 440240 100668 440292
rect 100720 440280 100726 440292
rect 136726 440280 136732 440292
rect 100720 440252 136732 440280
rect 100720 440240 100726 440252
rect 136726 440240 136732 440252
rect 136784 440240 136790 440292
rect 66990 439560 66996 439612
rect 67048 439600 67054 439612
rect 76558 439600 76564 439612
rect 67048 439572 76564 439600
rect 67048 439560 67054 439572
rect 76558 439560 76564 439572
rect 76616 439560 76622 439612
rect 53742 439492 53748 439544
rect 53800 439532 53806 439544
rect 57698 439532 57704 439544
rect 53800 439504 57704 439532
rect 53800 439492 53806 439504
rect 57698 439492 57704 439504
rect 57756 439532 57762 439544
rect 73154 439532 73160 439544
rect 57756 439504 73160 439532
rect 57756 439492 57762 439504
rect 73154 439492 73160 439504
rect 73212 439492 73218 439544
rect 91646 439152 91652 439204
rect 91704 439192 91710 439204
rect 91922 439192 91928 439204
rect 91704 439164 91928 439192
rect 91704 439152 91710 439164
rect 91922 439152 91928 439164
rect 91980 439152 91986 439204
rect 67358 439084 67364 439136
rect 67416 439124 67422 439136
rect 73338 439124 73344 439136
rect 67416 439096 73344 439124
rect 67416 439084 67422 439096
rect 73338 439084 73344 439096
rect 73396 439084 73402 439136
rect 110414 439124 110420 439136
rect 89686 439096 110420 439124
rect 43714 439016 43720 439068
rect 43772 439056 43778 439068
rect 45370 439056 45376 439068
rect 43772 439028 45376 439056
rect 43772 439016 43778 439028
rect 45370 439016 45376 439028
rect 45428 439056 45434 439068
rect 73890 439056 73896 439068
rect 45428 439028 73896 439056
rect 45428 439016 45434 439028
rect 73890 439016 73896 439028
rect 73948 439016 73954 439068
rect 84838 439016 84844 439068
rect 84896 439056 84902 439068
rect 89686 439056 89714 439096
rect 110414 439084 110420 439096
rect 110472 439084 110478 439136
rect 95234 439056 95240 439068
rect 84896 439028 89714 439056
rect 91848 439028 95240 439056
rect 84896 439016 84902 439028
rect 57882 438948 57888 439000
rect 57940 438988 57946 439000
rect 91646 438988 91652 439000
rect 57940 438960 91652 438988
rect 57940 438948 57946 438960
rect 91646 438948 91652 438960
rect 91704 438948 91710 439000
rect 11698 438880 11704 438932
rect 11756 438920 11762 438932
rect 91848 438920 91876 439028
rect 95234 439016 95240 439028
rect 95292 439056 95298 439068
rect 96430 439056 96436 439068
rect 95292 439028 96436 439056
rect 95292 439016 95298 439028
rect 96430 439016 96436 439028
rect 96488 439016 96494 439068
rect 103606 439016 103612 439068
rect 103664 439056 103670 439068
rect 106918 439056 106924 439068
rect 103664 439028 106924 439056
rect 103664 439016 103670 439028
rect 106918 439016 106924 439028
rect 106976 439016 106982 439068
rect 94038 438948 94044 439000
rect 94096 438988 94102 439000
rect 95142 438988 95148 439000
rect 94096 438960 95148 438988
rect 94096 438948 94102 438960
rect 95142 438948 95148 438960
rect 95200 438988 95206 439000
rect 128538 438988 128544 439000
rect 95200 438960 128544 438988
rect 95200 438948 95206 438960
rect 128538 438948 128544 438960
rect 128596 438948 128602 439000
rect 11756 438892 91876 438920
rect 11756 438880 11762 438892
rect 91922 438880 91928 438932
rect 91980 438920 91986 438932
rect 95878 438920 95884 438932
rect 91980 438892 95884 438920
rect 91980 438880 91986 438892
rect 95878 438880 95884 438892
rect 95936 438880 95942 438932
rect 96430 438880 96436 438932
rect 96488 438920 96494 438932
rect 121546 438920 121552 438932
rect 96488 438892 121552 438920
rect 96488 438880 96494 438892
rect 121546 438880 121552 438892
rect 121604 438880 121610 438932
rect 50982 438812 50988 438864
rect 51040 438852 51046 438864
rect 53558 438852 53564 438864
rect 51040 438824 53564 438852
rect 51040 438812 51046 438824
rect 53558 438812 53564 438824
rect 53616 438852 53622 438864
rect 83550 438852 83556 438864
rect 53616 438824 83556 438852
rect 53616 438812 53622 438824
rect 83550 438812 83556 438824
rect 83608 438812 83614 438864
rect 88978 438812 88984 438864
rect 89036 438852 89042 438864
rect 118786 438852 118792 438864
rect 89036 438824 118792 438852
rect 89036 438812 89042 438824
rect 118786 438812 118792 438824
rect 118844 438812 118850 438864
rect 73154 438744 73160 438796
rect 73212 438784 73218 438796
rect 82262 438784 82268 438796
rect 73212 438756 82268 438784
rect 73212 438744 73218 438756
rect 82262 438744 82268 438756
rect 82320 438744 82326 438796
rect 89990 438744 89996 438796
rect 90048 438784 90054 438796
rect 91002 438784 91008 438796
rect 90048 438756 91008 438784
rect 90048 438744 90054 438756
rect 91002 438744 91008 438756
rect 91060 438784 91066 438796
rect 118878 438784 118884 438796
rect 91060 438756 118884 438784
rect 91060 438744 91066 438756
rect 118878 438744 118884 438756
rect 118936 438744 118942 438796
rect 48130 438676 48136 438728
rect 48188 438716 48194 438728
rect 75822 438716 75828 438728
rect 48188 438688 75828 438716
rect 48188 438676 48194 438688
rect 75822 438676 75828 438688
rect 75880 438676 75886 438728
rect 99006 438676 99012 438728
rect 99064 438716 99070 438728
rect 99282 438716 99288 438728
rect 99064 438688 99288 438716
rect 99064 438676 99070 438688
rect 99282 438676 99288 438688
rect 99340 438716 99346 438728
rect 122926 438716 122932 438728
rect 99340 438688 122932 438716
rect 99340 438676 99346 438688
rect 122926 438676 122932 438688
rect 122984 438676 122990 438728
rect 80698 438608 80704 438660
rect 80756 438648 80762 438660
rect 104158 438648 104164 438660
rect 80756 438620 104164 438648
rect 80756 438608 80762 438620
rect 104158 438608 104164 438620
rect 104216 438608 104222 438660
rect 98362 438540 98368 438592
rect 98420 438580 98426 438592
rect 99190 438580 99196 438592
rect 98420 438552 99196 438580
rect 98420 438540 98426 438552
rect 99190 438540 99196 438552
rect 99248 438580 99254 438592
rect 114738 438580 114744 438592
rect 99248 438552 114744 438580
rect 99248 438540 99254 438552
rect 114738 438540 114744 438552
rect 114796 438540 114802 438592
rect 65886 438268 65892 438320
rect 65944 438308 65950 438320
rect 75178 438308 75184 438320
rect 65944 438280 75184 438308
rect 65944 438268 65950 438280
rect 75178 438268 75184 438280
rect 75236 438268 75242 438320
rect 56410 438200 56416 438252
rect 56468 438240 56474 438252
rect 73246 438240 73252 438252
rect 56468 438212 73252 438240
rect 56468 438200 56474 438212
rect 73246 438200 73252 438212
rect 73304 438200 73310 438252
rect 4798 438132 4804 438184
rect 4856 438172 4862 438184
rect 50982 438172 50988 438184
rect 4856 438144 50988 438172
rect 4856 438132 4862 438144
rect 50982 438132 50988 438144
rect 51040 438132 51046 438184
rect 57238 438132 57244 438184
rect 57296 438172 57302 438184
rect 91278 438172 91284 438184
rect 57296 438144 91284 438172
rect 57296 438132 57302 438144
rect 91278 438132 91284 438144
rect 91336 438132 91342 438184
rect 99650 438132 99656 438184
rect 99708 438172 99714 438184
rect 102042 438172 102048 438184
rect 99708 438144 102048 438172
rect 99708 438132 99714 438144
rect 102042 438132 102048 438144
rect 102100 438172 102106 438184
rect 124490 438172 124496 438184
rect 102100 438144 124496 438172
rect 102100 438132 102106 438144
rect 124490 438132 124496 438144
rect 124548 438132 124554 438184
rect 83550 437928 83556 437980
rect 83608 437968 83614 437980
rect 84838 437968 84844 437980
rect 83608 437940 84844 437968
rect 83608 437928 83614 437940
rect 84838 437928 84844 437940
rect 84896 437928 84902 437980
rect 89346 437724 89352 437776
rect 89404 437764 89410 437776
rect 91738 437764 91744 437776
rect 89404 437736 91744 437764
rect 89404 437724 89410 437736
rect 91738 437724 91744 437736
rect 91796 437724 91802 437776
rect 56226 437452 56232 437504
rect 56284 437492 56290 437504
rect 57238 437492 57244 437504
rect 56284 437464 57244 437492
rect 56284 437452 56290 437464
rect 57238 437452 57244 437464
rect 57296 437452 57302 437504
rect 54938 437384 54944 437436
rect 54996 437424 55002 437436
rect 85574 437424 85580 437436
rect 54996 437396 85580 437424
rect 54996 437384 55002 437396
rect 85574 437384 85580 437396
rect 85632 437424 85638 437436
rect 86770 437424 86776 437436
rect 85632 437396 86776 437424
rect 85632 437384 85638 437396
rect 86770 437384 86776 437396
rect 86828 437384 86834 437436
rect 100202 437424 100208 437436
rect 93826 437396 100208 437424
rect 46566 437316 46572 437368
rect 46624 437356 46630 437368
rect 78398 437356 78404 437368
rect 46624 437328 78404 437356
rect 46624 437316 46630 437328
rect 78398 437316 78404 437328
rect 78456 437316 78462 437368
rect 86218 437316 86224 437368
rect 86276 437356 86282 437368
rect 93826 437356 93854 437396
rect 100202 437384 100208 437396
rect 100260 437384 100266 437436
rect 86276 437328 93854 437356
rect 86276 437316 86282 437328
rect 94866 437316 94872 437368
rect 94924 437356 94930 437368
rect 120166 437356 120172 437368
rect 94924 437328 120172 437356
rect 94924 437316 94930 437328
rect 120166 437316 120172 437328
rect 120224 437316 120230 437368
rect 52086 437248 52092 437300
rect 52144 437288 52150 437300
rect 82906 437288 82912 437300
rect 52144 437260 82912 437288
rect 52144 437248 52150 437260
rect 82906 437248 82912 437260
rect 82964 437248 82970 437300
rect 97074 437248 97080 437300
rect 97132 437288 97138 437300
rect 97132 437260 113174 437288
rect 97132 437248 97138 437260
rect 44082 437180 44088 437232
rect 44140 437220 44146 437232
rect 55858 437220 55864 437232
rect 44140 437192 55864 437220
rect 44140 437180 44146 437192
rect 55858 437180 55864 437192
rect 55916 437220 55922 437232
rect 56410 437220 56416 437232
rect 55916 437192 56416 437220
rect 55916 437180 55922 437192
rect 56410 437180 56416 437192
rect 56468 437180 56474 437232
rect 58986 437180 58992 437232
rect 59044 437220 59050 437232
rect 81618 437220 81624 437232
rect 59044 437192 81624 437220
rect 59044 437180 59050 437192
rect 81618 437180 81624 437192
rect 81676 437180 81682 437232
rect 87690 437180 87696 437232
rect 87748 437220 87754 437232
rect 105630 437220 105636 437232
rect 87748 437192 105636 437220
rect 87748 437180 87754 437192
rect 105630 437180 105636 437192
rect 105688 437180 105694 437232
rect 113146 437220 113174 437260
rect 131298 437220 131304 437232
rect 113146 437192 131304 437220
rect 131298 437180 131304 437192
rect 131356 437180 131362 437232
rect 69198 436908 69204 436960
rect 69256 436948 69262 436960
rect 72418 436948 72424 436960
rect 69256 436920 72424 436948
rect 69256 436908 69262 436920
rect 72418 436908 72424 436920
rect 72476 436908 72482 436960
rect 39666 436704 39672 436756
rect 39724 436744 39730 436756
rect 46750 436744 46756 436756
rect 39724 436716 46756 436744
rect 39724 436704 39730 436716
rect 46750 436704 46756 436716
rect 46808 436744 46814 436756
rect 71682 436744 71688 436756
rect 46808 436716 71688 436744
rect 46808 436704 46814 436716
rect 71682 436704 71688 436716
rect 71740 436704 71746 436756
rect 78398 436432 78404 436484
rect 78456 436472 78462 436484
rect 83458 436472 83464 436484
rect 78456 436444 83464 436472
rect 78456 436432 78462 436444
rect 83458 436432 83464 436444
rect 83516 436432 83522 436484
rect 97074 436364 97080 436416
rect 97132 436404 97138 436416
rect 97902 436404 97908 436416
rect 97132 436376 97908 436404
rect 97132 436364 97138 436376
rect 97902 436364 97908 436376
rect 97960 436364 97966 436416
rect 50798 436024 50804 436076
rect 50856 436064 50862 436076
rect 78766 436064 78772 436076
rect 50856 436036 78772 436064
rect 50856 436024 50862 436036
rect 78766 436024 78772 436036
rect 78824 436024 78830 436076
rect 92566 436024 92572 436076
rect 92624 436064 92630 436076
rect 93670 436064 93676 436076
rect 92624 436036 93676 436064
rect 92624 436024 92630 436036
rect 93670 436024 93676 436036
rect 93728 436064 93734 436076
rect 109402 436064 109408 436076
rect 93728 436036 109408 436064
rect 93728 436024 93734 436036
rect 109402 436024 109408 436036
rect 109460 436024 109466 436076
rect 40954 434664 40960 434716
rect 41012 434704 41018 434716
rect 74534 434704 74540 434716
rect 41012 434676 74540 434704
rect 41012 434664 41018 434676
rect 74534 434664 74540 434676
rect 74592 434664 74598 434716
rect 56318 434596 56324 434648
rect 56376 434636 56382 434648
rect 71866 434636 71872 434648
rect 56376 434608 71872 434636
rect 56376 434596 56382 434608
rect 71866 434596 71872 434608
rect 71924 434636 71930 434648
rect 72602 434636 72608 434648
rect 71924 434608 72608 434636
rect 71924 434596 71930 434608
rect 72602 434596 72608 434608
rect 72660 434596 72666 434648
rect 59078 433984 59084 434036
rect 59136 434024 59142 434036
rect 69658 434024 69664 434036
rect 59136 433996 69664 434024
rect 59136 433984 59142 433996
rect 69658 433984 69664 433996
rect 69716 433984 69722 434036
rect 49510 433236 49516 433288
rect 49568 433276 49574 433288
rect 76466 433276 76472 433288
rect 49568 433248 76472 433276
rect 49568 433236 49574 433248
rect 76466 433236 76472 433248
rect 76524 433236 76530 433288
rect 42702 432556 42708 432608
rect 42760 432596 42766 432608
rect 49510 432596 49516 432608
rect 42760 432568 49516 432596
rect 42760 432556 42766 432568
rect 49510 432556 49516 432568
rect 49568 432556 49574 432608
rect 69014 432556 69020 432608
rect 69072 432596 69078 432608
rect 80790 432596 80796 432608
rect 69072 432568 80796 432596
rect 69072 432556 69078 432568
rect 80790 432556 80796 432568
rect 80848 432556 80854 432608
rect 100754 431264 100760 431316
rect 100812 431304 100818 431316
rect 104986 431304 104992 431316
rect 100812 431276 104992 431304
rect 100812 431264 100818 431276
rect 104986 431264 104992 431276
rect 105044 431264 105050 431316
rect 83458 431196 83464 431248
rect 83516 431236 83522 431248
rect 580166 431236 580172 431248
rect 83516 431208 580172 431236
rect 83516 431196 83522 431208
rect 580166 431196 580172 431208
rect 580224 431196 580230 431248
rect 69106 431060 69112 431112
rect 69164 431100 69170 431112
rect 71958 431100 71964 431112
rect 69164 431072 71964 431100
rect 69164 431060 69170 431072
rect 71958 431060 71964 431072
rect 72016 431060 72022 431112
rect 104986 430584 104992 430636
rect 105044 430624 105050 430636
rect 111150 430624 111156 430636
rect 105044 430596 111156 430624
rect 105044 430584 105050 430596
rect 111150 430584 111156 430596
rect 111208 430584 111214 430636
rect 3418 429836 3424 429888
rect 3476 429876 3482 429888
rect 100754 429876 100760 429888
rect 3476 429848 100760 429876
rect 3476 429836 3482 429848
rect 100754 429836 100760 429848
rect 100812 429836 100818 429888
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 113174 422328 113180 422340
rect 3568 422300 113180 422328
rect 3568 422288 3574 422300
rect 113174 422288 113180 422300
rect 113232 422288 113238 422340
rect 113174 421540 113180 421592
rect 113232 421580 113238 421592
rect 119430 421580 119436 421592
rect 113232 421552 119436 421580
rect 113232 421540 113238 421552
rect 119430 421540 119436 421552
rect 119488 421580 119494 421592
rect 120350 421580 120356 421592
rect 119488 421552 120356 421580
rect 119488 421540 119494 421552
rect 120350 421540 120356 421552
rect 120408 421540 120414 421592
rect 370498 418140 370504 418192
rect 370556 418180 370562 418192
rect 580166 418180 580172 418192
rect 370556 418152 580172 418180
rect 370556 418140 370562 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 99374 406784 99380 406836
rect 99432 406824 99438 406836
rect 100110 406824 100116 406836
rect 99432 406796 100116 406824
rect 99432 406784 99438 406796
rect 100110 406784 100116 406796
rect 100168 406784 100174 406836
rect 75914 406240 75920 406292
rect 75972 406280 75978 406292
rect 76558 406280 76564 406292
rect 75972 406252 76564 406280
rect 75972 406240 75978 406252
rect 76558 406240 76564 406252
rect 76616 406240 76622 406292
rect 76558 405764 76564 405816
rect 76616 405804 76622 405816
rect 173158 405804 173164 405816
rect 76616 405776 173164 405804
rect 76616 405764 76622 405776
rect 173158 405764 173164 405776
rect 173216 405764 173222 405816
rect 99374 405696 99380 405748
rect 99432 405736 99438 405748
rect 342254 405736 342260 405748
rect 99432 405708 342260 405736
rect 99432 405696 99438 405708
rect 342254 405696 342260 405708
rect 342312 405696 342318 405748
rect 95878 405016 95884 405068
rect 95936 405056 95942 405068
rect 128538 405056 128544 405068
rect 95936 405028 128544 405056
rect 95936 405016 95942 405028
rect 128538 405016 128544 405028
rect 128596 405016 128602 405068
rect 97902 404948 97908 405000
rect 97960 404988 97966 405000
rect 132586 404988 132592 405000
rect 97960 404960 132592 404988
rect 97960 404948 97966 404960
rect 132586 404948 132592 404960
rect 132644 404948 132650 405000
rect 544378 404336 544384 404388
rect 544436 404376 544442 404388
rect 580166 404376 580172 404388
rect 544436 404348 580172 404376
rect 544436 404336 544442 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 89806 403588 89812 403640
rect 89864 403628 89870 403640
rect 113266 403628 113272 403640
rect 89864 403600 113272 403628
rect 89864 403588 89870 403600
rect 113266 403588 113272 403600
rect 113324 403628 113330 403640
rect 353294 403628 353300 403640
rect 113324 403600 353300 403628
rect 113324 403588 113330 403600
rect 353294 403588 353300 403600
rect 353352 403588 353358 403640
rect 74534 402976 74540 403028
rect 74592 403016 74598 403028
rect 75178 403016 75184 403028
rect 74592 402988 75184 403016
rect 74592 402976 74598 402988
rect 75178 402976 75184 402988
rect 75236 403016 75242 403028
rect 153838 403016 153844 403028
rect 75236 402988 153844 403016
rect 75236 402976 75242 402988
rect 153838 402976 153844 402988
rect 153896 402976 153902 403028
rect 106182 402296 106188 402348
rect 106240 402336 106246 402348
rect 117590 402336 117596 402348
rect 106240 402308 117596 402336
rect 106240 402296 106246 402308
rect 117590 402296 117596 402308
rect 117648 402296 117654 402348
rect 45278 402228 45284 402280
rect 45336 402268 45342 402280
rect 85482 402268 85488 402280
rect 45336 402240 85488 402268
rect 45336 402228 45342 402240
rect 85482 402228 85488 402240
rect 85540 402228 85546 402280
rect 94038 402228 94044 402280
rect 94096 402268 94102 402280
rect 120258 402268 120264 402280
rect 94096 402240 120264 402268
rect 94096 402228 94102 402240
rect 120258 402228 120264 402240
rect 120316 402228 120322 402280
rect 80790 401616 80796 401668
rect 80848 401656 80854 401668
rect 327074 401656 327080 401668
rect 80848 401628 327080 401656
rect 80848 401616 80854 401628
rect 327074 401616 327080 401628
rect 327132 401616 327138 401668
rect 99190 401004 99196 401056
rect 99248 401044 99254 401056
rect 131298 401044 131304 401056
rect 99248 401016 131304 401044
rect 99248 401004 99254 401016
rect 131298 401004 131304 401016
rect 131356 401004 131362 401056
rect 92658 400936 92664 400988
rect 92716 400976 92722 400988
rect 111702 400976 111708 400988
rect 92716 400948 111708 400976
rect 92716 400936 92722 400948
rect 111702 400936 111708 400948
rect 111760 400976 111766 400988
rect 166258 400976 166264 400988
rect 111760 400948 166264 400976
rect 111760 400936 111766 400948
rect 166258 400936 166264 400948
rect 166316 400936 166322 400988
rect 97994 400868 98000 400920
rect 98052 400908 98058 400920
rect 117498 400908 117504 400920
rect 98052 400880 117504 400908
rect 98052 400868 98058 400880
rect 117498 400868 117504 400880
rect 117556 400908 117562 400920
rect 351914 400908 351920 400920
rect 117556 400880 351920 400908
rect 117556 400868 117562 400880
rect 351914 400868 351920 400880
rect 351972 400868 351978 400920
rect 69198 400188 69204 400240
rect 69256 400228 69262 400240
rect 226978 400228 226984 400240
rect 69256 400200 226984 400228
rect 69256 400188 69262 400200
rect 226978 400188 226984 400200
rect 227036 400188 227042 400240
rect 56410 399576 56416 399628
rect 56468 399616 56474 399628
rect 84838 399616 84844 399628
rect 56468 399588 84844 399616
rect 56468 399576 56474 399588
rect 84838 399576 84844 399588
rect 84896 399576 84902 399628
rect 54938 399508 54944 399560
rect 54996 399548 55002 399560
rect 85574 399548 85580 399560
rect 54996 399520 85580 399548
rect 54996 399508 55002 399520
rect 85574 399508 85580 399520
rect 85632 399508 85638 399560
rect 43898 399440 43904 399492
rect 43956 399480 43962 399492
rect 87506 399480 87512 399492
rect 43956 399452 87512 399480
rect 43956 399440 43962 399452
rect 87506 399440 87512 399452
rect 87564 399480 87570 399492
rect 88242 399480 88248 399492
rect 87564 399452 88248 399480
rect 87564 399440 87570 399452
rect 88242 399440 88248 399452
rect 88300 399440 88306 399492
rect 95142 399440 95148 399492
rect 95200 399480 95206 399492
rect 127342 399480 127348 399492
rect 95200 399452 127348 399480
rect 95200 399440 95206 399452
rect 127342 399440 127348 399452
rect 127400 399440 127406 399492
rect 88242 398896 88248 398948
rect 88300 398936 88306 398948
rect 159358 398936 159364 398948
rect 88300 398908 159364 398936
rect 88300 398896 88306 398908
rect 159358 398896 159364 398908
rect 159416 398896 159422 398948
rect 72418 398828 72424 398880
rect 72476 398868 72482 398880
rect 149238 398868 149244 398880
rect 72476 398840 149244 398868
rect 72476 398828 72482 398840
rect 149238 398828 149244 398840
rect 149296 398868 149302 398880
rect 204898 398868 204904 398880
rect 149296 398840 204904 398868
rect 149296 398828 149302 398840
rect 204898 398828 204904 398840
rect 204956 398828 204962 398880
rect 117222 398216 117228 398268
rect 117280 398256 117286 398268
rect 125870 398256 125876 398268
rect 117280 398228 125876 398256
rect 117280 398216 117286 398228
rect 125870 398216 125876 398228
rect 125928 398216 125934 398268
rect 98546 398148 98552 398200
rect 98604 398188 98610 398200
rect 127066 398188 127072 398200
rect 98604 398160 127072 398188
rect 98604 398148 98610 398160
rect 127066 398148 127072 398160
rect 127124 398188 127130 398200
rect 157978 398188 157984 398200
rect 127124 398160 157984 398188
rect 127124 398148 127130 398160
rect 157978 398148 157984 398160
rect 158036 398148 158042 398200
rect 53650 398080 53656 398132
rect 53708 398120 53714 398132
rect 69290 398120 69296 398132
rect 53708 398092 69296 398120
rect 53708 398080 53714 398092
rect 69290 398080 69296 398092
rect 69348 398080 69354 398132
rect 88334 398080 88340 398132
rect 88392 398120 88398 398132
rect 123294 398120 123300 398132
rect 88392 398092 123300 398120
rect 88392 398080 88398 398092
rect 123294 398080 123300 398092
rect 123352 398120 123358 398132
rect 162118 398120 162124 398132
rect 123352 398092 162124 398120
rect 123352 398080 123358 398092
rect 162118 398080 162124 398092
rect 162176 398080 162182 398132
rect 116578 397576 116584 397588
rect 55186 397548 116584 397576
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 50982 397508 50988 397520
rect 3476 397480 50988 397508
rect 3476 397468 3482 397480
rect 50982 397468 50988 397480
rect 51040 397508 51046 397520
rect 55186 397508 55214 397548
rect 116578 397536 116584 397548
rect 116636 397576 116642 397588
rect 117222 397576 117228 397588
rect 116636 397548 117228 397576
rect 116636 397536 116642 397548
rect 117222 397536 117228 397548
rect 117280 397536 117286 397588
rect 51040 397480 55214 397508
rect 51040 397468 51046 397480
rect 69290 397468 69296 397520
rect 69348 397508 69354 397520
rect 268378 397508 268384 397520
rect 69348 397480 268384 397508
rect 69348 397468 69354 397480
rect 268378 397468 268384 397480
rect 268436 397468 268442 397520
rect 108850 396856 108856 396908
rect 108908 396896 108914 396908
rect 117498 396896 117504 396908
rect 108908 396868 117504 396896
rect 108908 396856 108914 396868
rect 117498 396856 117504 396868
rect 117556 396856 117562 396908
rect 43806 396788 43812 396840
rect 43864 396828 43870 396840
rect 71866 396828 71872 396840
rect 43864 396800 71872 396828
rect 43864 396788 43870 396800
rect 71866 396788 71872 396800
rect 71924 396788 71930 396840
rect 99282 396788 99288 396840
rect 99340 396828 99346 396840
rect 131206 396828 131212 396840
rect 99340 396800 131212 396828
rect 99340 396788 99346 396800
rect 131206 396788 131212 396800
rect 131264 396788 131270 396840
rect 53466 396720 53472 396772
rect 53524 396760 53530 396772
rect 83550 396760 83556 396772
rect 53524 396732 83556 396760
rect 53524 396720 53530 396732
rect 83550 396720 83556 396732
rect 83608 396720 83614 396772
rect 93762 396720 93768 396772
rect 93820 396760 93826 396772
rect 127158 396760 127164 396772
rect 93820 396732 127164 396760
rect 93820 396720 93826 396732
rect 127158 396720 127164 396732
rect 127216 396720 127222 396772
rect 102134 396584 102140 396636
rect 102192 396624 102198 396636
rect 102778 396624 102784 396636
rect 102192 396596 102784 396624
rect 102192 396584 102198 396596
rect 102778 396584 102784 396596
rect 102836 396584 102842 396636
rect 41138 396040 41144 396092
rect 41196 396080 41202 396092
rect 102134 396080 102140 396092
rect 41196 396052 102140 396080
rect 41196 396040 41202 396052
rect 102134 396040 102140 396052
rect 102192 396040 102198 396092
rect 69106 395972 69112 396024
rect 69164 396012 69170 396024
rect 69658 396012 69664 396024
rect 69164 395984 69664 396012
rect 69164 395972 69170 395984
rect 69658 395972 69664 395984
rect 69716 395972 69722 396024
rect 106918 395972 106924 396024
rect 106976 396012 106982 396024
rect 134702 396012 134708 396024
rect 106976 395984 134708 396012
rect 106976 395972 106982 395984
rect 134702 395972 134708 395984
rect 134760 395972 134766 396024
rect 276014 395972 276020 396024
rect 276072 396012 276078 396024
rect 276658 396012 276664 396024
rect 276072 395984 276664 396012
rect 276072 395972 276078 395984
rect 276658 395972 276664 395984
rect 276716 395972 276722 396024
rect 127250 395468 127256 395480
rect 122806 395440 127256 395468
rect 45278 395360 45284 395412
rect 45336 395400 45342 395412
rect 78674 395400 78680 395412
rect 45336 395372 78680 395400
rect 45336 395360 45342 395372
rect 78674 395360 78680 395372
rect 78732 395360 78738 395412
rect 95970 395360 95976 395412
rect 96028 395400 96034 395412
rect 122806 395400 122834 395440
rect 127250 395428 127256 395440
rect 127308 395468 127314 395480
rect 142338 395468 142344 395480
rect 127308 395440 142344 395468
rect 127308 395428 127314 395440
rect 142338 395428 142344 395440
rect 142396 395428 142402 395480
rect 150434 395400 150440 395412
rect 96028 395372 122834 395400
rect 132466 395372 150440 395400
rect 96028 395360 96034 395372
rect 48038 395292 48044 395344
rect 48096 395332 48102 395344
rect 82814 395332 82820 395344
rect 48096 395304 82820 395332
rect 48096 395292 48102 395304
rect 82814 395292 82820 395304
rect 82872 395292 82878 395344
rect 96706 395292 96712 395344
rect 96764 395332 96770 395344
rect 128446 395332 128452 395344
rect 96764 395304 128452 395332
rect 96764 395292 96770 395304
rect 128446 395292 128452 395304
rect 128504 395332 128510 395344
rect 132466 395332 132494 395372
rect 150434 395360 150440 395372
rect 150492 395360 150498 395412
rect 128504 395304 132494 395332
rect 128504 395292 128510 395304
rect 134702 395292 134708 395344
rect 134760 395332 134766 395344
rect 276014 395332 276020 395344
rect 134760 395304 276020 395332
rect 134760 395292 134766 395304
rect 276014 395292 276020 395304
rect 276072 395292 276078 395344
rect 292482 395292 292488 395344
rect 292540 395332 292546 395344
rect 385678 395332 385684 395344
rect 292540 395304 385684 395332
rect 292540 395292 292546 395304
rect 385678 395292 385684 395304
rect 385736 395292 385742 395344
rect 82814 394748 82820 394800
rect 82872 394788 82878 394800
rect 82998 394788 83004 394800
rect 82872 394760 83004 394788
rect 82872 394748 82878 394760
rect 82998 394748 83004 394760
rect 83056 394788 83062 394800
rect 126330 394788 126336 394800
rect 83056 394760 126336 394788
rect 83056 394748 83062 394760
rect 126330 394748 126336 394760
rect 126388 394748 126394 394800
rect 69106 394680 69112 394732
rect 69164 394720 69170 394732
rect 231854 394720 231860 394732
rect 69164 394692 231860 394720
rect 69164 394680 69170 394692
rect 231854 394680 231860 394692
rect 231912 394680 231918 394732
rect 68738 394612 68744 394664
rect 68796 394652 68802 394664
rect 68922 394652 68928 394664
rect 68796 394624 68928 394652
rect 68796 394612 68802 394624
rect 68922 394612 68928 394624
rect 68980 394612 68986 394664
rect 53098 394068 53104 394120
rect 53156 394108 53162 394120
rect 75362 394108 75368 394120
rect 53156 394080 75368 394108
rect 53156 394068 53162 394080
rect 75362 394068 75368 394080
rect 75420 394068 75426 394120
rect 52362 394000 52368 394052
rect 52420 394040 52426 394052
rect 82906 394040 82912 394052
rect 52420 394012 82912 394040
rect 52420 394000 52426 394012
rect 82906 394000 82912 394012
rect 82964 394000 82970 394052
rect 101398 394000 101404 394052
rect 101456 394040 101462 394052
rect 106274 394040 106280 394052
rect 101456 394012 106280 394040
rect 101456 394000 101462 394012
rect 106274 394000 106280 394012
rect 106332 394000 106338 394052
rect 108298 394000 108304 394052
rect 108356 394040 108362 394052
rect 135438 394040 135444 394052
rect 108356 394012 135444 394040
rect 108356 394000 108362 394012
rect 135438 394000 135444 394012
rect 135496 394000 135502 394052
rect 49510 393932 49516 393984
rect 49568 393972 49574 393984
rect 80698 393972 80704 393984
rect 49568 393944 80704 393972
rect 49568 393932 49574 393944
rect 80698 393932 80704 393944
rect 80756 393932 80762 393984
rect 95234 393932 95240 393984
rect 95292 393972 95298 393984
rect 128998 393972 129004 393984
rect 95292 393944 129004 393972
rect 95292 393932 95298 393944
rect 128998 393932 129004 393944
rect 129056 393932 129062 393984
rect 82814 393456 82820 393508
rect 82872 393496 82878 393508
rect 83090 393496 83096 393508
rect 82872 393468 83096 393496
rect 82872 393456 82878 393468
rect 83090 393456 83096 393468
rect 83148 393496 83154 393508
rect 138014 393496 138020 393508
rect 83148 393468 138020 393496
rect 83148 393456 83154 393468
rect 138014 393456 138020 393468
rect 138072 393456 138078 393508
rect 75362 393388 75368 393440
rect 75420 393428 75426 393440
rect 134150 393428 134156 393440
rect 75420 393400 134156 393428
rect 75420 393388 75426 393400
rect 134150 393388 134156 393400
rect 134208 393388 134214 393440
rect 135438 393388 135444 393440
rect 135496 393428 135502 393440
rect 316678 393428 316684 393440
rect 135496 393400 316684 393428
rect 135496 393388 135502 393400
rect 316678 393388 316684 393400
rect 316736 393388 316742 393440
rect 68922 393320 68928 393372
rect 68980 393360 68986 393372
rect 278038 393360 278044 393372
rect 68980 393332 278044 393360
rect 68980 393320 68986 393332
rect 278038 393320 278044 393332
rect 278096 393320 278102 393372
rect 41230 393252 41236 393304
rect 41288 393292 41294 393304
rect 82814 393292 82820 393304
rect 41288 393264 82820 393292
rect 41288 393252 41294 393264
rect 82814 393252 82820 393264
rect 82872 393252 82878 393304
rect 110874 392776 110880 392828
rect 110932 392816 110938 392828
rect 125686 392816 125692 392828
rect 110932 392788 125692 392816
rect 110932 392776 110938 392788
rect 125686 392776 125692 392788
rect 125744 392776 125750 392828
rect 114278 392708 114284 392760
rect 114336 392748 114342 392760
rect 139394 392748 139400 392760
rect 114336 392720 139400 392748
rect 114336 392708 114342 392720
rect 139394 392708 139400 392720
rect 139452 392748 139458 392760
rect 146938 392748 146944 392760
rect 139452 392720 146944 392748
rect 139452 392708 139458 392720
rect 146938 392708 146944 392720
rect 146996 392708 147002 392760
rect 57698 392640 57704 392692
rect 57756 392680 57762 392692
rect 87598 392680 87604 392692
rect 57756 392652 87604 392680
rect 57756 392640 57762 392652
rect 87598 392640 87604 392652
rect 87656 392640 87662 392692
rect 104526 392640 104532 392692
rect 104584 392680 104590 392692
rect 134058 392680 134064 392692
rect 104584 392652 134064 392680
rect 104584 392640 104590 392652
rect 134058 392640 134064 392652
rect 134116 392640 134122 392692
rect 36906 392572 36912 392624
rect 36964 392612 36970 392624
rect 70394 392612 70400 392624
rect 36964 392584 70400 392612
rect 36964 392572 36970 392584
rect 70394 392572 70400 392584
rect 70452 392572 70458 392624
rect 94130 392572 94136 392624
rect 94188 392612 94194 392624
rect 124398 392612 124404 392624
rect 94188 392584 124404 392612
rect 94188 392572 94194 392584
rect 124398 392572 124404 392584
rect 124456 392612 124462 392624
rect 152090 392612 152096 392624
rect 124456 392584 152096 392612
rect 124456 392572 124462 392584
rect 152090 392572 152096 392584
rect 152148 392572 152154 392624
rect 47854 392096 47860 392148
rect 47912 392136 47918 392148
rect 110874 392136 110880 392148
rect 47912 392108 110880 392136
rect 47912 392096 47918 392108
rect 110874 392096 110880 392108
rect 110932 392096 110938 392148
rect 134058 392096 134064 392148
rect 134116 392136 134122 392148
rect 136818 392136 136824 392148
rect 134116 392108 136824 392136
rect 134116 392096 134122 392108
rect 136818 392096 136824 392108
rect 136876 392096 136882 392148
rect 106274 392028 106280 392080
rect 106332 392068 106338 392080
rect 360194 392068 360200 392080
rect 106332 392040 360200 392068
rect 106332 392028 106338 392040
rect 360194 392028 360200 392040
rect 360252 392028 360258 392080
rect 324314 392000 324320 392012
rect 67560 391972 324320 392000
rect 53558 391892 53564 391944
rect 53616 391932 53622 391944
rect 57330 391932 57336 391944
rect 53616 391904 57336 391932
rect 53616 391892 53622 391904
rect 57330 391892 57336 391904
rect 57388 391932 57394 391944
rect 67560 391932 67588 391972
rect 324314 391960 324320 391972
rect 324372 391960 324378 392012
rect 57388 391904 67588 391932
rect 57388 391892 57394 391904
rect 91002 391892 91008 391944
rect 91060 391932 91066 391944
rect 92566 391932 92572 391944
rect 91060 391904 92572 391932
rect 91060 391892 91066 391904
rect 92566 391892 92572 391904
rect 92624 391892 92630 391944
rect 47946 391280 47952 391332
rect 48004 391320 48010 391332
rect 76006 391320 76012 391332
rect 48004 391292 76012 391320
rect 48004 391280 48010 391292
rect 76006 391280 76012 391292
rect 76064 391280 76070 391332
rect 103330 391280 103336 391332
rect 103388 391320 103394 391332
rect 116118 391320 116124 391332
rect 103388 391292 116124 391320
rect 103388 391280 103394 391292
rect 116118 391280 116124 391292
rect 116176 391280 116182 391332
rect 55122 391212 55128 391264
rect 55180 391252 55186 391264
rect 88978 391252 88984 391264
rect 55180 391224 88984 391252
rect 55180 391212 55186 391224
rect 88978 391212 88984 391224
rect 89036 391212 89042 391264
rect 102042 391212 102048 391264
rect 102100 391252 102106 391264
rect 132678 391252 132684 391264
rect 102100 391224 132684 391252
rect 102100 391212 102106 391224
rect 132678 391212 132684 391224
rect 132736 391252 132742 391264
rect 133690 391252 133696 391264
rect 132736 391224 133696 391252
rect 132736 391212 132742 391224
rect 133690 391212 133696 391224
rect 133748 391212 133754 391264
rect 113910 390668 113916 390720
rect 113968 390708 113974 390720
rect 167638 390708 167644 390720
rect 113968 390680 167644 390708
rect 113968 390668 113974 390680
rect 167638 390668 167644 390680
rect 167696 390668 167702 390720
rect 67542 390600 67548 390652
rect 67600 390640 67606 390652
rect 136634 390640 136640 390652
rect 67600 390612 136640 390640
rect 67600 390600 67606 390612
rect 136634 390600 136640 390612
rect 136692 390600 136698 390652
rect 137278 390600 137284 390652
rect 137336 390640 137342 390652
rect 140774 390640 140780 390652
rect 137336 390612 140780 390640
rect 137336 390600 137342 390612
rect 140774 390600 140780 390612
rect 140832 390600 140838 390652
rect 52270 390532 52276 390584
rect 52328 390572 52334 390584
rect 79318 390572 79324 390584
rect 52328 390544 79324 390572
rect 52328 390532 52334 390544
rect 79318 390532 79324 390544
rect 79376 390532 79382 390584
rect 133690 390532 133696 390584
rect 133748 390572 133754 390584
rect 313274 390572 313280 390584
rect 133748 390544 313280 390572
rect 133748 390532 133754 390544
rect 313274 390532 313280 390544
rect 313332 390532 313338 390584
rect 56502 390464 56508 390516
rect 56560 390504 56566 390516
rect 67542 390504 67548 390516
rect 56560 390476 67548 390504
rect 56560 390464 56566 390476
rect 67542 390464 67548 390476
rect 67600 390464 67606 390516
rect 111058 390056 111064 390108
rect 111116 390096 111122 390108
rect 114922 390096 114928 390108
rect 111116 390068 114928 390096
rect 111116 390056 111122 390068
rect 114922 390056 114928 390068
rect 114980 390056 114986 390108
rect 92566 389920 92572 389972
rect 92624 389960 92630 389972
rect 121454 389960 121460 389972
rect 92624 389932 121460 389960
rect 92624 389920 92630 389932
rect 121454 389920 121460 389932
rect 121512 389920 121518 389972
rect 39942 389852 39948 389904
rect 40000 389892 40006 389904
rect 69566 389892 69572 389904
rect 40000 389864 69572 389892
rect 40000 389852 40006 389864
rect 69566 389852 69572 389864
rect 69624 389852 69630 389904
rect 102594 389852 102600 389904
rect 102652 389892 102658 389904
rect 135346 389892 135352 389904
rect 102652 389864 135352 389892
rect 102652 389852 102658 389864
rect 135346 389852 135352 389864
rect 135404 389892 135410 389904
rect 136542 389892 136548 389904
rect 135404 389864 136548 389892
rect 135404 389852 135410 389864
rect 136542 389852 136548 389864
rect 136600 389852 136606 389904
rect 38470 389784 38476 389836
rect 38528 389824 38534 389836
rect 109034 389824 109040 389836
rect 38528 389796 109040 389824
rect 38528 389784 38534 389796
rect 109034 389784 109040 389796
rect 109092 389784 109098 389836
rect 119430 389784 119436 389836
rect 119488 389824 119494 389836
rect 143810 389824 143816 389836
rect 119488 389796 143816 389824
rect 119488 389784 119494 389796
rect 143810 389784 143816 389796
rect 143868 389784 143874 389836
rect 115842 389444 115848 389496
rect 115900 389484 115906 389496
rect 119430 389484 119436 389496
rect 115900 389456 119436 389484
rect 115900 389444 115906 389456
rect 119430 389444 119436 389456
rect 119488 389444 119494 389496
rect 69566 389376 69572 389428
rect 69624 389416 69630 389428
rect 84470 389416 84476 389428
rect 69624 389388 84476 389416
rect 69624 389376 69630 389388
rect 84470 389376 84476 389388
rect 84528 389376 84534 389428
rect 120718 389376 120724 389428
rect 120776 389416 120782 389428
rect 121638 389416 121644 389428
rect 120776 389388 121644 389416
rect 120776 389376 120782 389388
rect 121638 389376 121644 389388
rect 121696 389376 121702 389428
rect 54754 389308 54760 389360
rect 54812 389348 54818 389360
rect 57882 389348 57888 389360
rect 54812 389320 57888 389348
rect 54812 389308 54818 389320
rect 57882 389308 57888 389320
rect 57940 389348 57946 389360
rect 80606 389348 80612 389360
rect 57940 389320 80612 389348
rect 57940 389308 57946 389320
rect 80606 389308 80612 389320
rect 80664 389308 80670 389360
rect 89714 389308 89720 389360
rect 89772 389348 89778 389360
rect 90358 389348 90364 389360
rect 89772 389320 90364 389348
rect 89772 389308 89778 389320
rect 90358 389308 90364 389320
rect 90416 389308 90422 389360
rect 110322 389308 110328 389360
rect 110380 389348 110386 389360
rect 137278 389348 137284 389360
rect 110380 389320 137284 389348
rect 110380 389308 110386 389320
rect 137278 389308 137284 389320
rect 137336 389308 137342 389360
rect 48958 389240 48964 389292
rect 49016 389280 49022 389292
rect 120718 389280 120724 389292
rect 49016 389252 120724 389280
rect 49016 389240 49022 389252
rect 120718 389240 120724 389252
rect 120776 389240 120782 389292
rect 121454 389240 121460 389292
rect 121512 389280 121518 389292
rect 122098 389280 122104 389292
rect 121512 389252 122104 389280
rect 121512 389240 121518 389252
rect 122098 389240 122104 389252
rect 122156 389280 122162 389292
rect 222838 389280 222844 389292
rect 122156 389252 222844 389280
rect 122156 389240 122162 389252
rect 222838 389240 222844 389252
rect 222896 389240 222902 389292
rect 56318 389172 56324 389224
rect 56376 389212 56382 389224
rect 56502 389212 56508 389224
rect 56376 389184 56508 389212
rect 56376 389172 56382 389184
rect 56502 389172 56508 389184
rect 56560 389172 56566 389224
rect 63218 389172 63224 389224
rect 63276 389212 63282 389224
rect 253198 389212 253204 389224
rect 63276 389184 253204 389212
rect 63276 389172 63282 389184
rect 253198 389172 253204 389184
rect 253256 389172 253262 389224
rect 102778 389104 102784 389156
rect 102836 389144 102842 389156
rect 103606 389144 103612 389156
rect 102836 389116 103612 389144
rect 102836 389104 102842 389116
rect 103606 389104 103612 389116
rect 103664 389144 103670 389156
rect 104802 389144 104808 389156
rect 103664 389116 104808 389144
rect 103664 389104 103670 389116
rect 104802 389104 104808 389116
rect 104860 389104 104866 389156
rect 77294 388832 77300 388884
rect 77352 388872 77358 388884
rect 77570 388872 77576 388884
rect 77352 388844 77576 388872
rect 77352 388832 77358 388844
rect 77570 388832 77576 388844
rect 77628 388832 77634 388884
rect 100018 388764 100024 388816
rect 100076 388804 100082 388816
rect 101398 388804 101404 388816
rect 100076 388776 101404 388804
rect 100076 388764 100082 388776
rect 101398 388764 101404 388776
rect 101456 388764 101462 388816
rect 50798 388560 50804 388612
rect 50856 388600 50862 388612
rect 54846 388600 54852 388612
rect 50856 388572 54852 388600
rect 50856 388560 50862 388572
rect 54846 388560 54852 388572
rect 54904 388600 54910 388612
rect 69750 388600 69756 388612
rect 54904 388572 69756 388600
rect 54904 388560 54910 388572
rect 69750 388560 69756 388572
rect 69808 388560 69814 388612
rect 58618 388492 58624 388544
rect 58676 388532 58682 388544
rect 81434 388532 81440 388544
rect 58676 388504 81440 388532
rect 58676 388492 58682 388504
rect 81434 388492 81440 388504
rect 81492 388492 81498 388544
rect 48222 388424 48228 388476
rect 48280 388464 48286 388476
rect 78214 388464 78220 388476
rect 48280 388436 78220 388464
rect 48280 388424 48286 388436
rect 78214 388424 78220 388436
rect 78272 388424 78278 388476
rect 95878 388220 95884 388272
rect 95936 388260 95942 388272
rect 102134 388260 102140 388272
rect 95936 388232 102140 388260
rect 95936 388220 95942 388232
rect 102134 388220 102140 388232
rect 102192 388220 102198 388272
rect 104802 388220 104808 388272
rect 104860 388260 104866 388272
rect 266998 388260 267004 388272
rect 104860 388232 267004 388260
rect 104860 388220 104866 388232
rect 266998 388220 267004 388232
rect 267056 388220 267062 388272
rect 109126 388152 109132 388204
rect 109184 388192 109190 388204
rect 117958 388192 117964 388204
rect 109184 388164 117964 388192
rect 109184 388152 109190 388164
rect 117958 388152 117964 388164
rect 118016 388152 118022 388204
rect 119448 388164 122834 388192
rect 94866 388084 94872 388136
rect 94924 388124 94930 388136
rect 109034 388124 109040 388136
rect 94924 388096 109040 388124
rect 94924 388084 94930 388096
rect 109034 388084 109040 388096
rect 109092 388084 109098 388136
rect 112162 388084 112168 388136
rect 112220 388124 112226 388136
rect 119448 388124 119476 388164
rect 112220 388096 119476 388124
rect 122806 388124 122834 388164
rect 122806 388096 142154 388124
rect 112220 388084 112226 388096
rect 4798 388016 4804 388068
rect 4856 388056 4862 388068
rect 72418 388056 72424 388068
rect 4856 388028 72424 388056
rect 4856 388016 4862 388028
rect 72418 388016 72424 388028
rect 72476 388016 72482 388068
rect 81434 388016 81440 388068
rect 81492 388056 81498 388068
rect 82354 388056 82360 388068
rect 81492 388028 82360 388056
rect 81492 388016 81498 388028
rect 82354 388016 82360 388028
rect 82412 388056 82418 388068
rect 119430 388056 119436 388068
rect 82412 388028 119436 388056
rect 82412 388016 82418 388028
rect 119430 388016 119436 388028
rect 119488 388016 119494 388068
rect 142126 388056 142154 388096
rect 143902 388056 143908 388068
rect 142126 388028 143908 388056
rect 143902 388016 143908 388028
rect 143960 388056 143966 388068
rect 159450 388056 159456 388068
rect 143960 388028 159456 388056
rect 143960 388016 143966 388028
rect 159450 388016 159456 388028
rect 159508 388016 159514 388068
rect 53650 387948 53656 388000
rect 53708 387988 53714 388000
rect 77570 387988 77576 388000
rect 53708 387960 77576 387988
rect 53708 387948 53714 387960
rect 77570 387948 77576 387960
rect 77628 387948 77634 388000
rect 93302 387948 93308 388000
rect 93360 387988 93366 388000
rect 119522 387988 119528 388000
rect 93360 387960 119528 387988
rect 93360 387948 93366 387960
rect 119522 387948 119528 387960
rect 119580 387948 119586 388000
rect 39942 387880 39948 387932
rect 40000 387920 40006 387932
rect 73338 387920 73344 387932
rect 40000 387892 73344 387920
rect 40000 387880 40006 387892
rect 73338 387880 73344 387892
rect 73396 387880 73402 387932
rect 108942 387880 108948 387932
rect 109000 387920 109006 387932
rect 115750 387920 115756 387932
rect 109000 387892 115756 387920
rect 109000 387880 109006 387892
rect 115750 387880 115756 387892
rect 115808 387880 115814 387932
rect 117958 387880 117964 387932
rect 118016 387920 118022 387932
rect 178678 387920 178684 387932
rect 118016 387892 178684 387920
rect 118016 387880 118022 387892
rect 178678 387880 178684 387892
rect 178736 387880 178742 387932
rect 70394 387812 70400 387864
rect 70452 387852 70458 387864
rect 80054 387852 80060 387864
rect 70452 387824 80060 387852
rect 70452 387812 70458 387824
rect 80054 387812 80060 387824
rect 80112 387812 80118 387864
rect 91554 387812 91560 387864
rect 91612 387852 91618 387864
rect 103514 387852 103520 387864
rect 91612 387824 103520 387852
rect 91612 387812 91618 387824
rect 103514 387812 103520 387824
rect 103572 387852 103578 387864
rect 104802 387852 104808 387864
rect 103572 387824 104808 387852
rect 103572 387812 103578 387824
rect 104802 387812 104808 387824
rect 104860 387812 104866 387864
rect 106182 387812 106188 387864
rect 106240 387852 106246 387864
rect 111794 387852 111800 387864
rect 106240 387824 111800 387852
rect 106240 387812 106246 387824
rect 111794 387812 111800 387824
rect 111852 387812 111858 387864
rect 114922 387812 114928 387864
rect 114980 387852 114986 387864
rect 184198 387852 184204 387864
rect 114980 387824 184204 387852
rect 114980 387812 114986 387824
rect 184198 387812 184204 387824
rect 184256 387812 184262 387864
rect 54846 387132 54852 387184
rect 54904 387172 54910 387184
rect 83458 387172 83464 387184
rect 54904 387144 83464 387172
rect 54904 387132 54910 387144
rect 83458 387132 83464 387144
rect 83516 387132 83522 387184
rect 104802 387132 104808 387184
rect 104860 387172 104866 387184
rect 118694 387172 118700 387184
rect 104860 387144 118700 387172
rect 104860 387132 104866 387144
rect 118694 387132 118700 387144
rect 118752 387132 118758 387184
rect 46658 387064 46664 387116
rect 46716 387104 46722 387116
rect 78766 387104 78772 387116
rect 46716 387076 78772 387104
rect 46716 387064 46722 387076
rect 78766 387064 78772 387076
rect 78824 387064 78830 387116
rect 111150 387064 111156 387116
rect 111208 387104 111214 387116
rect 130010 387104 130016 387116
rect 111208 387076 130016 387104
rect 111208 387064 111214 387076
rect 130010 387064 130016 387076
rect 130068 387064 130074 387116
rect 107562 386588 107568 386640
rect 107620 386628 107626 386640
rect 126238 386628 126244 386640
rect 107620 386600 126244 386628
rect 107620 386588 107626 386600
rect 126238 386588 126244 386600
rect 126296 386588 126302 386640
rect 56502 386520 56508 386572
rect 56560 386560 56566 386572
rect 87046 386560 87052 386572
rect 56560 386532 87052 386560
rect 56560 386520 56566 386532
rect 87046 386520 87052 386532
rect 87104 386520 87110 386572
rect 104434 386520 104440 386572
rect 104492 386560 104498 386572
rect 104618 386560 104624 386572
rect 104492 386532 104624 386560
rect 104492 386520 104498 386532
rect 104618 386520 104624 386532
rect 104676 386560 104682 386572
rect 124398 386560 124404 386572
rect 104676 386532 124404 386560
rect 104676 386520 104682 386532
rect 124398 386520 124404 386532
rect 124456 386520 124462 386572
rect 34238 386452 34244 386504
rect 34296 386492 34302 386504
rect 80514 386492 80520 386504
rect 34296 386464 80520 386492
rect 34296 386452 34302 386464
rect 80514 386452 80520 386464
rect 80572 386452 80578 386504
rect 118694 386452 118700 386504
rect 118752 386492 118758 386504
rect 264238 386492 264244 386504
rect 118752 386464 264244 386492
rect 118752 386452 118758 386464
rect 264238 386452 264244 386464
rect 264296 386452 264302 386504
rect 78214 386384 78220 386436
rect 78272 386424 78278 386436
rect 126974 386424 126980 386436
rect 78272 386396 126980 386424
rect 78272 386384 78278 386396
rect 126974 386384 126980 386396
rect 127032 386424 127038 386436
rect 301498 386424 301504 386436
rect 127032 386396 301504 386424
rect 127032 386384 127038 386396
rect 301498 386384 301504 386396
rect 301556 386384 301562 386436
rect 38562 386316 38568 386368
rect 38620 386356 38626 386368
rect 58618 386356 58624 386368
rect 38620 386328 58624 386356
rect 38620 386316 38626 386328
rect 58618 386316 58624 386328
rect 58676 386316 58682 386368
rect 109034 386316 109040 386368
rect 109092 386356 109098 386368
rect 125594 386356 125600 386368
rect 109092 386328 125600 386356
rect 109092 386316 109098 386328
rect 125594 386316 125600 386328
rect 125652 386356 125658 386368
rect 126882 386356 126888 386368
rect 125652 386328 126888 386356
rect 125652 386316 125658 386328
rect 126882 386316 126888 386328
rect 126940 386316 126946 386368
rect 45370 385840 45376 385892
rect 45428 385880 45434 385892
rect 49602 385880 49608 385892
rect 45428 385852 49608 385880
rect 45428 385840 45434 385852
rect 49602 385840 49608 385852
rect 49660 385840 49666 385892
rect 49326 385704 49332 385756
rect 49384 385744 49390 385756
rect 81526 385744 81532 385756
rect 49384 385716 81532 385744
rect 49384 385704 49390 385716
rect 81526 385704 81532 385716
rect 81584 385704 81590 385756
rect 126882 385704 126888 385756
rect 126940 385744 126946 385756
rect 155218 385744 155224 385756
rect 126940 385716 155224 385744
rect 126940 385704 126946 385716
rect 155218 385704 155224 385716
rect 155276 385704 155282 385756
rect 52086 385636 52092 385688
rect 52144 385676 52150 385688
rect 86310 385676 86316 385688
rect 52144 385648 86316 385676
rect 52144 385636 52150 385648
rect 86310 385636 86316 385648
rect 86368 385636 86374 385688
rect 91738 385636 91744 385688
rect 91796 385676 91802 385688
rect 125686 385676 125692 385688
rect 91796 385648 125692 385676
rect 91796 385636 91802 385648
rect 125686 385636 125692 385648
rect 125744 385636 125750 385688
rect 71774 385336 71780 385348
rect 64846 385308 71780 385336
rect 35710 385092 35716 385144
rect 35768 385132 35774 385144
rect 64846 385132 64874 385308
rect 71774 385296 71780 385308
rect 71832 385296 71838 385348
rect 92934 385336 92940 385348
rect 84166 385308 92940 385336
rect 35768 385104 64874 385132
rect 35768 385092 35774 385104
rect 49602 385024 49608 385076
rect 49660 385064 49666 385076
rect 84166 385064 84194 385308
rect 92934 385296 92940 385308
rect 92992 385296 92998 385348
rect 101306 385296 101312 385348
rect 101364 385336 101370 385348
rect 101364 385308 103514 385336
rect 101364 385296 101370 385308
rect 49660 385036 84194 385064
rect 103486 385064 103514 385308
rect 122282 385092 122288 385144
rect 122340 385132 122346 385144
rect 123754 385132 123760 385144
rect 122340 385104 123760 385132
rect 122340 385092 122346 385104
rect 123754 385092 123760 385104
rect 123812 385092 123818 385144
rect 135898 385064 135904 385076
rect 103486 385036 135904 385064
rect 49660 385024 49666 385036
rect 135898 385024 135904 385036
rect 135956 385024 135962 385076
rect 60550 384276 60556 384328
rect 60608 384316 60614 384328
rect 67634 384316 67640 384328
rect 60608 384288 67640 384316
rect 60608 384276 60614 384288
rect 67634 384276 67640 384288
rect 67692 384276 67698 384328
rect 118510 384276 118516 384328
rect 118568 384316 118574 384328
rect 147582 384316 147588 384328
rect 118568 384288 147588 384316
rect 118568 384276 118574 384288
rect 147582 384276 147588 384288
rect 147640 384276 147646 384328
rect 118050 383664 118056 383716
rect 118108 383704 118114 383716
rect 139394 383704 139400 383716
rect 118108 383676 139400 383704
rect 118108 383664 118114 383676
rect 139394 383664 139400 383676
rect 139452 383664 139458 383716
rect 119522 382916 119528 382968
rect 119580 382956 119586 382968
rect 297358 382956 297364 382968
rect 119580 382928 297364 382956
rect 119580 382916 119586 382928
rect 297358 382916 297364 382928
rect 297416 382916 297422 382968
rect 126054 382304 126060 382356
rect 126112 382344 126118 382356
rect 129918 382344 129924 382356
rect 126112 382316 129924 382344
rect 126112 382304 126118 382316
rect 129918 382304 129924 382316
rect 129976 382304 129982 382356
rect 39850 382236 39856 382288
rect 39908 382276 39914 382288
rect 67634 382276 67640 382288
rect 39908 382248 67640 382276
rect 39908 382236 39914 382248
rect 67634 382236 67640 382248
rect 67692 382236 67698 382288
rect 118142 382236 118148 382288
rect 118200 382276 118206 382288
rect 127618 382276 127624 382288
rect 118200 382248 127624 382276
rect 118200 382236 118206 382248
rect 127618 382236 127624 382248
rect 127676 382236 127682 382288
rect 118602 382168 118608 382220
rect 118660 382208 118666 382220
rect 141050 382208 141056 382220
rect 118660 382180 141056 382208
rect 118660 382168 118666 382180
rect 141050 382168 141056 382180
rect 141108 382168 141114 382220
rect 141050 381556 141056 381608
rect 141108 381596 141114 381608
rect 181438 381596 181444 381608
rect 141108 381568 181444 381596
rect 141108 381556 141114 381568
rect 181438 381556 181444 381568
rect 181496 381556 181502 381608
rect 118602 381488 118608 381540
rect 118660 381528 118666 381540
rect 125594 381528 125600 381540
rect 118660 381500 125600 381528
rect 118660 381488 118666 381500
rect 125594 381488 125600 381500
rect 125652 381528 125658 381540
rect 126054 381528 126060 381540
rect 125652 381500 126060 381528
rect 125652 381488 125658 381500
rect 126054 381488 126060 381500
rect 126112 381488 126118 381540
rect 147582 381488 147588 381540
rect 147640 381528 147646 381540
rect 349798 381528 349804 381540
rect 147640 381500 349804 381528
rect 147640 381488 147646 381500
rect 349798 381488 349804 381500
rect 349856 381488 349862 381540
rect 118602 380332 118608 380384
rect 118660 380372 118666 380384
rect 122466 380372 122472 380384
rect 118660 380344 122472 380372
rect 118660 380332 118666 380344
rect 122466 380332 122472 380344
rect 122524 380332 122530 380384
rect 115290 380264 115296 380316
rect 115348 380304 115354 380316
rect 117314 380304 117320 380316
rect 115348 380276 117320 380304
rect 115348 380264 115354 380276
rect 117314 380264 117320 380276
rect 117372 380264 117378 380316
rect 117682 380128 117688 380180
rect 117740 380168 117746 380180
rect 118326 380168 118332 380180
rect 117740 380140 118332 380168
rect 117740 380128 117746 380140
rect 118326 380128 118332 380140
rect 118384 380168 118390 380180
rect 192478 380168 192484 380180
rect 118384 380140 192484 380168
rect 118384 380128 118390 380140
rect 192478 380128 192484 380140
rect 192536 380128 192542 380180
rect 65978 379652 65984 379704
rect 66036 379692 66042 379704
rect 67726 379692 67732 379704
rect 66036 379664 67732 379692
rect 66036 379652 66042 379664
rect 67726 379652 67732 379664
rect 67784 379652 67790 379704
rect 60642 379584 60648 379636
rect 60700 379624 60706 379636
rect 66162 379624 66168 379636
rect 60700 379596 66168 379624
rect 60700 379584 60706 379596
rect 66162 379584 66168 379596
rect 66220 379624 66226 379636
rect 67634 379624 67640 379636
rect 66220 379596 67640 379624
rect 66220 379584 66226 379596
rect 67634 379584 67640 379596
rect 67692 379584 67698 379636
rect 48038 379516 48044 379568
rect 48096 379556 48102 379568
rect 69658 379556 69664 379568
rect 48096 379528 69664 379556
rect 48096 379516 48102 379528
rect 69658 379516 69664 379528
rect 69716 379516 69722 379568
rect 263594 379516 263600 379568
rect 263652 379556 263658 379568
rect 264238 379556 264244 379568
rect 263652 379528 264244 379556
rect 263652 379516 263658 379528
rect 264238 379516 264244 379528
rect 264296 379556 264302 379568
rect 483658 379556 483664 379568
rect 264296 379528 483664 379556
rect 264296 379516 264302 379528
rect 483658 379516 483664 379528
rect 483716 379516 483722 379568
rect 35618 379448 35624 379500
rect 35676 379488 35682 379500
rect 65610 379488 65616 379500
rect 35676 379460 65616 379488
rect 35676 379448 35682 379460
rect 65610 379448 65616 379460
rect 65668 379488 65674 379500
rect 65978 379488 65984 379500
rect 65668 379460 65984 379488
rect 65668 379448 65674 379460
rect 65978 379448 65984 379460
rect 66036 379448 66042 379500
rect 42610 379380 42616 379432
rect 42668 379420 42674 379432
rect 69842 379420 69848 379432
rect 42668 379392 69848 379420
rect 42668 379380 42674 379392
rect 69842 379380 69848 379392
rect 69900 379380 69906 379432
rect 37182 378768 37188 378820
rect 37240 378808 37246 378820
rect 69198 378808 69204 378820
rect 37240 378780 69204 378808
rect 37240 378768 37246 378780
rect 69198 378768 69204 378780
rect 69256 378768 69262 378820
rect 118602 378700 118608 378752
rect 118660 378740 118666 378752
rect 124122 378740 124128 378752
rect 118660 378712 124128 378740
rect 118660 378700 118666 378712
rect 124122 378700 124128 378712
rect 124180 378700 124186 378752
rect 233878 378292 233884 378344
rect 233936 378332 233942 378344
rect 357434 378332 357440 378344
rect 233936 378304 357440 378332
rect 233936 378292 233942 378304
rect 357434 378292 357440 378304
rect 357492 378292 357498 378344
rect 118050 378224 118056 378276
rect 118108 378264 118114 378276
rect 244274 378264 244280 378276
rect 118108 378236 244280 378264
rect 118108 378224 118114 378236
rect 244274 378224 244280 378236
rect 244332 378224 244338 378276
rect 253198 378224 253204 378276
rect 253256 378264 253262 378276
rect 347774 378264 347780 378276
rect 253256 378236 347780 378264
rect 253256 378224 253262 378236
rect 347774 378224 347780 378236
rect 347832 378224 347838 378276
rect 174538 378156 174544 378208
rect 174596 378196 174602 378208
rect 323118 378196 323124 378208
rect 174596 378168 323124 378196
rect 174596 378156 174602 378168
rect 323118 378156 323124 378168
rect 323176 378156 323182 378208
rect 353938 378156 353944 378208
rect 353996 378196 354002 378208
rect 580166 378196 580172 378208
rect 353996 378168 580172 378196
rect 353996 378156 354002 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 57882 378088 57888 378140
rect 57940 378128 57946 378140
rect 61470 378128 61476 378140
rect 57940 378100 61476 378128
rect 57940 378088 57946 378100
rect 61470 378088 61476 378100
rect 61528 378128 61534 378140
rect 67634 378128 67640 378140
rect 61528 378100 67640 378128
rect 61528 378088 61534 378100
rect 67634 378088 67640 378100
rect 67692 378088 67698 378140
rect 244274 377408 244280 377460
rect 244332 377448 244338 377460
rect 265250 377448 265256 377460
rect 244332 377420 265256 377448
rect 244332 377408 244338 377420
rect 265250 377408 265256 377420
rect 265308 377408 265314 377460
rect 266998 377408 267004 377460
rect 267056 377448 267062 377460
rect 308398 377448 308404 377460
rect 267056 377420 308404 377448
rect 267056 377408 267062 377420
rect 308398 377408 308404 377420
rect 308456 377408 308462 377460
rect 249702 376796 249708 376848
rect 249760 376836 249766 376848
rect 358814 376836 358820 376848
rect 249760 376808 358820 376836
rect 249760 376796 249766 376808
rect 358814 376796 358820 376808
rect 358872 376796 358878 376848
rect 117866 376728 117872 376780
rect 117924 376768 117930 376780
rect 121454 376768 121460 376780
rect 117924 376740 121460 376768
rect 117924 376728 117930 376740
rect 121454 376728 121460 376740
rect 121512 376728 121518 376780
rect 197262 376728 197268 376780
rect 197320 376768 197326 376780
rect 511994 376768 512000 376780
rect 197320 376740 512000 376768
rect 197320 376728 197326 376740
rect 511994 376728 512000 376740
rect 512052 376728 512058 376780
rect 52178 376660 52184 376712
rect 52236 376700 52242 376712
rect 66898 376700 66904 376712
rect 52236 376672 66904 376700
rect 52236 376660 52242 376672
rect 66898 376660 66904 376672
rect 66956 376700 66962 376712
rect 67542 376700 67548 376712
rect 66956 376672 67548 376700
rect 66956 376660 66962 376672
rect 67542 376660 67548 376672
rect 67600 376660 67606 376712
rect 118602 376660 118608 376712
rect 118660 376700 118666 376712
rect 146294 376700 146300 376712
rect 118660 376672 146300 376700
rect 118660 376660 118666 376672
rect 146294 376660 146300 376672
rect 146352 376700 146358 376712
rect 149054 376700 149060 376712
rect 146352 376672 149060 376700
rect 146352 376660 146358 376672
rect 149054 376660 149060 376672
rect 149112 376660 149118 376712
rect 119430 376048 119436 376100
rect 119488 376088 119494 376100
rect 154574 376088 154580 376100
rect 119488 376060 154580 376088
rect 119488 376048 119494 376060
rect 154574 376048 154580 376060
rect 154632 376048 154638 376100
rect 120166 375980 120172 376032
rect 120224 376020 120230 376032
rect 143718 376020 143724 376032
rect 120224 375992 143724 376020
rect 120224 375980 120230 375992
rect 143718 375980 143724 375992
rect 143776 376020 143782 376032
rect 319530 376020 319536 376032
rect 143776 375992 319536 376020
rect 143776 375980 143782 375992
rect 319530 375980 319536 375992
rect 319588 375980 319594 376032
rect 61378 375368 61384 375420
rect 61436 375408 61442 375420
rect 64690 375408 64696 375420
rect 61436 375380 64696 375408
rect 61436 375368 61442 375380
rect 64690 375368 64696 375380
rect 64748 375408 64754 375420
rect 67634 375408 67640 375420
rect 64748 375380 67640 375408
rect 64748 375368 64754 375380
rect 67634 375368 67640 375380
rect 67692 375368 67698 375420
rect 118510 375368 118516 375420
rect 118568 375408 118574 375420
rect 120166 375408 120172 375420
rect 118568 375380 120172 375408
rect 118568 375368 118574 375380
rect 120166 375368 120172 375380
rect 120224 375368 120230 375420
rect 265250 375368 265256 375420
rect 265308 375408 265314 375420
rect 403618 375408 403624 375420
rect 265308 375380 403624 375408
rect 265308 375368 265314 375380
rect 403618 375368 403624 375380
rect 403676 375368 403682 375420
rect 61838 375300 61844 375352
rect 61896 375340 61902 375352
rect 63402 375340 63408 375352
rect 61896 375312 63408 375340
rect 61896 375300 61902 375312
rect 63402 375300 63408 375312
rect 63460 375300 63466 375352
rect 118602 375300 118608 375352
rect 118660 375340 118666 375352
rect 133874 375340 133880 375352
rect 118660 375312 133880 375340
rect 118660 375300 118666 375312
rect 133874 375300 133880 375312
rect 133932 375340 133938 375352
rect 135162 375340 135168 375352
rect 133932 375312 135168 375340
rect 133932 375300 133938 375312
rect 135162 375300 135168 375312
rect 135220 375300 135226 375352
rect 62022 374620 62028 374672
rect 62080 374660 62086 374672
rect 65886 374660 65892 374672
rect 62080 374632 65892 374660
rect 62080 374620 62086 374632
rect 65886 374620 65892 374632
rect 65944 374660 65950 374672
rect 67634 374660 67640 374672
rect 65944 374632 67640 374660
rect 65944 374620 65950 374632
rect 67634 374620 67640 374632
rect 67692 374620 67698 374672
rect 121454 374620 121460 374672
rect 121512 374660 121518 374672
rect 155954 374660 155960 374672
rect 121512 374632 155960 374660
rect 121512 374620 121518 374632
rect 155954 374620 155960 374632
rect 156012 374620 156018 374672
rect 140038 374280 140044 374332
rect 140096 374320 140102 374332
rect 140682 374320 140688 374332
rect 140096 374292 140688 374320
rect 140096 374280 140102 374292
rect 140682 374280 140688 374292
rect 140740 374280 140746 374332
rect 224218 374212 224224 374264
rect 224276 374252 224282 374264
rect 340874 374252 340880 374264
rect 224276 374224 340880 374252
rect 224276 374212 224282 374224
rect 340874 374212 340880 374224
rect 340932 374212 340938 374264
rect 155954 374144 155960 374196
rect 156012 374184 156018 374196
rect 320082 374184 320088 374196
rect 156012 374156 320088 374184
rect 156012 374144 156018 374156
rect 320082 374144 320088 374156
rect 320140 374144 320146 374196
rect 327166 374116 327172 374128
rect 142126 374088 327172 374116
rect 63402 374008 63408 374060
rect 63460 374048 63466 374060
rect 67634 374048 67640 374060
rect 63460 374020 67640 374048
rect 63460 374008 63466 374020
rect 67634 374008 67640 374020
rect 67692 374008 67698 374060
rect 140682 374008 140688 374060
rect 140740 374048 140746 374060
rect 142126 374048 142154 374088
rect 327166 374076 327172 374088
rect 327224 374076 327230 374128
rect 140740 374020 142154 374048
rect 140740 374008 140746 374020
rect 204898 374008 204904 374060
rect 204956 374048 204962 374060
rect 209774 374048 209780 374060
rect 204956 374020 209780 374048
rect 204956 374008 204962 374020
rect 209774 374008 209780 374020
rect 209832 374048 209838 374060
rect 471974 374048 471980 374060
rect 209832 374020 471980 374048
rect 209832 374008 209838 374020
rect 471974 374008 471980 374020
rect 472032 374008 472038 374060
rect 137370 373668 137376 373720
rect 137428 373708 137434 373720
rect 138290 373708 138296 373720
rect 137428 373680 138296 373708
rect 137428 373668 137434 373680
rect 138290 373668 138296 373680
rect 138348 373668 138354 373720
rect 59262 373260 59268 373312
rect 59320 373300 59326 373312
rect 67634 373300 67640 373312
rect 59320 373272 67640 373300
rect 59320 373260 59326 373272
rect 67634 373260 67640 373272
rect 67692 373260 67698 373312
rect 117314 373260 117320 373312
rect 117372 373300 117378 373312
rect 185578 373300 185584 373312
rect 117372 373272 185584 373300
rect 117372 373260 117378 373272
rect 185578 373260 185584 373272
rect 185636 373260 185642 373312
rect 193950 372784 193956 372836
rect 194008 372824 194014 372836
rect 282914 372824 282920 372836
rect 194008 372796 282920 372824
rect 194008 372784 194014 372796
rect 282914 372784 282920 372796
rect 282972 372784 282978 372836
rect 177390 372716 177396 372768
rect 177448 372756 177454 372768
rect 333974 372756 333980 372768
rect 177448 372728 333980 372756
rect 177448 372716 177454 372728
rect 333974 372716 333980 372728
rect 334032 372756 334038 372768
rect 334618 372756 334624 372768
rect 334032 372728 334624 372756
rect 334032 372716 334038 372728
rect 334618 372716 334624 372728
rect 334676 372716 334682 372768
rect 123478 372648 123484 372700
rect 123536 372688 123542 372700
rect 321738 372688 321744 372700
rect 123536 372660 321744 372688
rect 123536 372648 123542 372660
rect 321738 372648 321744 372660
rect 321796 372648 321802 372700
rect 118050 372580 118056 372632
rect 118108 372620 118114 372632
rect 121454 372620 121460 372632
rect 118108 372592 121460 372620
rect 118108 372580 118114 372592
rect 121454 372580 121460 372592
rect 121512 372580 121518 372632
rect 138290 372580 138296 372632
rect 138348 372620 138354 372632
rect 339494 372620 339500 372632
rect 138348 372592 339500 372620
rect 138348 372580 138354 372592
rect 339494 372580 339500 372592
rect 339552 372580 339558 372632
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 48958 372552 48964 372564
rect 3292 372524 48964 372552
rect 3292 372512 3298 372524
rect 48958 372512 48964 372524
rect 49016 372512 49022 372564
rect 61930 371832 61936 371884
rect 61988 371872 61994 371884
rect 67634 371872 67640 371884
rect 61988 371844 67640 371872
rect 61988 371832 61994 371844
rect 67634 371832 67640 371844
rect 67692 371832 67698 371884
rect 142798 371832 142804 371884
rect 142856 371872 142862 371884
rect 150618 371872 150624 371884
rect 142856 371844 150624 371872
rect 142856 371832 142862 371844
rect 150618 371832 150624 371844
rect 150676 371872 150682 371884
rect 212534 371872 212540 371884
rect 150676 371844 212540 371872
rect 150676 371832 150682 371844
rect 212534 371832 212540 371844
rect 212592 371872 212598 371884
rect 213822 371872 213828 371884
rect 212592 371844 213828 371872
rect 212592 371832 212598 371844
rect 213822 371832 213828 371844
rect 213880 371832 213886 371884
rect 276658 371424 276664 371476
rect 276716 371464 276722 371476
rect 354674 371464 354680 371476
rect 276716 371436 354680 371464
rect 276716 371424 276722 371436
rect 354674 371424 354680 371436
rect 354732 371424 354738 371476
rect 200758 371356 200764 371408
rect 200816 371396 200822 371408
rect 324498 371396 324504 371408
rect 200816 371368 324504 371396
rect 200816 371356 200822 371368
rect 324498 371356 324504 371368
rect 324556 371356 324562 371408
rect 213822 371288 213828 371340
rect 213880 371328 213886 371340
rect 417418 371328 417424 371340
rect 213880 371300 417424 371328
rect 213880 371288 213886 371300
rect 417418 371288 417424 371300
rect 417476 371288 417482 371340
rect 117866 371220 117872 371272
rect 117924 371260 117930 371272
rect 338758 371260 338764 371272
rect 117924 371232 338764 371260
rect 117924 371220 117930 371232
rect 338758 371220 338764 371232
rect 338816 371220 338822 371272
rect 41046 371152 41052 371204
rect 41104 371192 41110 371204
rect 69290 371192 69296 371204
rect 41104 371164 69296 371192
rect 41104 371152 41110 371164
rect 69290 371152 69296 371164
rect 69348 371152 69354 371204
rect 118602 370540 118608 370592
rect 118660 370580 118666 370592
rect 129826 370580 129832 370592
rect 118660 370552 129832 370580
rect 118660 370540 118666 370552
rect 129826 370540 129832 370552
rect 129884 370540 129890 370592
rect 121454 370472 121460 370524
rect 121512 370512 121518 370524
rect 337378 370512 337384 370524
rect 121512 370484 337384 370512
rect 121512 370472 121518 370484
rect 337378 370472 337384 370484
rect 337436 370472 337442 370524
rect 177482 369996 177488 370048
rect 177540 370036 177546 370048
rect 305086 370036 305092 370048
rect 177540 370008 305092 370036
rect 177540 369996 177546 370008
rect 305086 369996 305092 370008
rect 305144 369996 305150 370048
rect 118234 369928 118240 369980
rect 118292 369968 118298 369980
rect 121454 369968 121460 369980
rect 118292 369940 121460 369968
rect 118292 369928 118298 369940
rect 121454 369928 121460 369940
rect 121512 369928 121518 369980
rect 162210 369928 162216 369980
rect 162268 369968 162274 369980
rect 323210 369968 323216 369980
rect 162268 369940 323216 369968
rect 162268 369928 162274 369940
rect 323210 369928 323216 369940
rect 323268 369928 323274 369980
rect 166350 369860 166356 369912
rect 166408 369900 166414 369912
rect 242158 369900 242164 369912
rect 166408 369872 242164 369900
rect 166408 369860 166414 369872
rect 242158 369860 242164 369872
rect 242216 369860 242222 369912
rect 244642 369860 244648 369912
rect 244700 369900 244706 369912
rect 244918 369900 244924 369912
rect 244700 369872 244924 369900
rect 244700 369860 244706 369872
rect 244918 369860 244924 369872
rect 244976 369900 244982 369912
rect 517514 369900 517520 369912
rect 244976 369872 517520 369900
rect 244976 369860 244982 369872
rect 517514 369860 517520 369872
rect 517572 369860 517578 369912
rect 118602 369792 118608 369844
rect 118660 369832 118666 369844
rect 122650 369832 122656 369844
rect 118660 369804 122656 369832
rect 118660 369792 118666 369804
rect 122650 369792 122656 369804
rect 122708 369832 122714 369844
rect 124306 369832 124312 369844
rect 122708 369804 124312 369832
rect 122708 369792 122714 369804
rect 124306 369792 124312 369804
rect 124364 369792 124370 369844
rect 66070 369452 66076 369504
rect 66128 369492 66134 369504
rect 68370 369492 68376 369504
rect 66128 369464 68376 369492
rect 66128 369452 66134 369464
rect 68370 369452 68376 369464
rect 68428 369452 68434 369504
rect 121454 369112 121460 369164
rect 121512 369152 121518 369164
rect 255314 369152 255320 369164
rect 121512 369124 255320 369152
rect 121512 369112 121518 369124
rect 255314 369112 255320 369124
rect 255372 369112 255378 369164
rect 119430 368772 119436 368824
rect 119488 368812 119494 368824
rect 269850 368812 269856 368824
rect 119488 368784 269856 368812
rect 119488 368772 119494 368784
rect 269850 368772 269856 368784
rect 269908 368812 269914 368824
rect 352006 368812 352012 368824
rect 269908 368784 352012 368812
rect 269908 368772 269914 368784
rect 352006 368772 352012 368784
rect 352064 368772 352070 368824
rect 124950 368704 124956 368756
rect 125008 368744 125014 368756
rect 312538 368744 312544 368756
rect 125008 368716 312544 368744
rect 125008 368704 125014 368716
rect 312538 368704 312544 368716
rect 312596 368704 312602 368756
rect 255314 368636 255320 368688
rect 255372 368676 255378 368688
rect 464338 368676 464344 368688
rect 255372 368648 464344 368676
rect 255372 368636 255378 368648
rect 464338 368636 464344 368648
rect 464396 368636 464402 368688
rect 119338 368568 119344 368620
rect 119396 368608 119402 368620
rect 335354 368608 335360 368620
rect 119396 368580 335360 368608
rect 119396 368568 119402 368580
rect 335354 368568 335360 368580
rect 335412 368568 335418 368620
rect 50338 368500 50344 368552
rect 50396 368540 50402 368552
rect 55030 368540 55036 368552
rect 50396 368512 55036 368540
rect 50396 368500 50402 368512
rect 55030 368500 55036 368512
rect 55088 368540 55094 368552
rect 67634 368540 67640 368552
rect 55088 368512 67640 368540
rect 55088 368500 55094 368512
rect 67634 368500 67640 368512
rect 67692 368500 67698 368552
rect 223482 368500 223488 368552
rect 223540 368540 223546 368552
rect 468478 368540 468484 368552
rect 223540 368512 468484 368540
rect 223540 368500 223546 368512
rect 468478 368500 468484 368512
rect 468536 368500 468542 368552
rect 127618 368432 127624 368484
rect 127676 368472 127682 368484
rect 151814 368472 151820 368484
rect 127676 368444 151820 368472
rect 127676 368432 127682 368444
rect 151814 368432 151820 368444
rect 151872 368472 151878 368484
rect 197262 368472 197268 368484
rect 151872 368444 197268 368472
rect 151872 368432 151878 368444
rect 197262 368432 197268 368444
rect 197320 368472 197326 368484
rect 197998 368472 198004 368484
rect 197320 368444 198004 368472
rect 197320 368432 197326 368444
rect 197998 368432 198004 368444
rect 198056 368432 198062 368484
rect 118602 367888 118608 367940
rect 118660 367928 118666 367940
rect 122834 367928 122840 367940
rect 118660 367900 122840 367928
rect 118660 367888 118666 367900
rect 122834 367888 122840 367900
rect 122892 367888 122898 367940
rect 209038 367344 209044 367396
rect 209096 367384 209102 367396
rect 345014 367384 345020 367396
rect 209096 367356 345020 367384
rect 209096 367344 209102 367356
rect 345014 367344 345020 367356
rect 345072 367344 345078 367396
rect 180242 367276 180248 367328
rect 180300 367316 180306 367328
rect 325786 367316 325792 367328
rect 180300 367288 325792 367316
rect 180300 367276 180306 367288
rect 325786 367276 325792 367288
rect 325844 367276 325850 367328
rect 222838 367208 222844 367260
rect 222896 367248 222902 367260
rect 385678 367248 385684 367260
rect 222896 367220 385684 367248
rect 222896 367208 222902 367220
rect 385678 367208 385684 367220
rect 385736 367208 385742 367260
rect 160738 367140 160744 367192
rect 160796 367180 160802 367192
rect 238202 367180 238208 367192
rect 160796 367152 238208 367180
rect 160796 367140 160802 367152
rect 238202 367140 238208 367152
rect 238260 367140 238266 367192
rect 297358 367140 297364 367192
rect 297416 367180 297422 367192
rect 471238 367180 471244 367192
rect 297416 367152 471244 367180
rect 297416 367140 297422 367152
rect 471238 367140 471244 367152
rect 471296 367140 471302 367192
rect 123570 367072 123576 367124
rect 123628 367112 123634 367124
rect 321646 367112 321652 367124
rect 123628 367084 321652 367112
rect 123628 367072 123634 367084
rect 321646 367072 321652 367084
rect 321704 367072 321710 367124
rect 56318 367004 56324 367056
rect 56376 367044 56382 367056
rect 67634 367044 67640 367056
rect 56376 367016 67640 367044
rect 56376 367004 56382 367016
rect 67634 367004 67640 367016
rect 67692 367004 67698 367056
rect 118602 367004 118608 367056
rect 118660 367044 118666 367056
rect 142154 367044 142160 367056
rect 118660 367016 142160 367044
rect 118660 367004 118666 367016
rect 142154 367004 142160 367016
rect 142212 367044 142218 367056
rect 146294 367044 146300 367056
rect 142212 367016 146300 367044
rect 142212 367004 142218 367016
rect 146294 367004 146300 367016
rect 146352 367004 146358 367056
rect 261846 366052 261852 366104
rect 261904 366092 261910 366104
rect 320174 366092 320180 366104
rect 261904 366064 320180 366092
rect 261904 366052 261910 366064
rect 320174 366052 320180 366064
rect 320232 366052 320238 366104
rect 199378 365984 199384 366036
rect 199436 366024 199442 366036
rect 227714 366024 227720 366036
rect 199436 365996 227720 366024
rect 199436 365984 199442 365996
rect 227714 365984 227720 365996
rect 227772 365984 227778 366036
rect 259362 365984 259368 366036
rect 259420 366024 259426 366036
rect 349154 366024 349160 366036
rect 259420 365996 349160 366024
rect 259420 365984 259426 365996
rect 349154 365984 349160 365996
rect 349212 365984 349218 366036
rect 171778 365916 171784 365968
rect 171836 365956 171842 365968
rect 295334 365956 295340 365968
rect 171836 365928 295340 365956
rect 171836 365916 171842 365928
rect 295334 365916 295340 365928
rect 295392 365916 295398 365968
rect 304994 365916 305000 365968
rect 305052 365956 305058 365968
rect 350534 365956 350540 365968
rect 305052 365928 350540 365956
rect 305052 365916 305058 365928
rect 350534 365916 350540 365928
rect 350592 365916 350598 365968
rect 189718 365848 189724 365900
rect 189776 365888 189782 365900
rect 331306 365888 331312 365900
rect 189776 365860 331312 365888
rect 189776 365848 189782 365860
rect 331306 365848 331312 365860
rect 331364 365848 331370 365900
rect 125042 365780 125048 365832
rect 125100 365820 125106 365832
rect 293402 365820 293408 365832
rect 125100 365792 293408 365820
rect 125100 365780 125106 365792
rect 293402 365780 293408 365792
rect 293460 365780 293466 365832
rect 295334 365780 295340 365832
rect 295392 365820 295398 365832
rect 295978 365820 295984 365832
rect 295392 365792 295984 365820
rect 295392 365780 295398 365792
rect 295978 365780 295984 365792
rect 296036 365820 296042 365832
rect 346394 365820 346400 365832
rect 296036 365792 346400 365820
rect 296036 365780 296042 365792
rect 346394 365780 346400 365792
rect 346452 365780 346458 365832
rect 148410 365712 148416 365764
rect 148468 365752 148474 365764
rect 209038 365752 209044 365764
rect 148468 365724 209044 365752
rect 148468 365712 148474 365724
rect 209038 365712 209044 365724
rect 209096 365712 209102 365764
rect 216582 365712 216588 365764
rect 216640 365752 216646 365764
rect 510614 365752 510620 365764
rect 216640 365724 510620 365752
rect 216640 365712 216646 365724
rect 510614 365712 510620 365724
rect 510672 365712 510678 365764
rect 60366 365644 60372 365696
rect 60424 365684 60430 365696
rect 66070 365684 66076 365696
rect 60424 365656 66076 365684
rect 60424 365644 60430 365656
rect 66070 365644 66076 365656
rect 66128 365644 66134 365696
rect 117866 365644 117872 365696
rect 117924 365684 117930 365696
rect 138198 365684 138204 365696
rect 117924 365656 138204 365684
rect 117924 365644 117930 365656
rect 138198 365644 138204 365656
rect 138256 365644 138262 365696
rect 117406 364964 117412 365016
rect 117464 365004 117470 365016
rect 145006 365004 145012 365016
rect 117464 364976 145012 365004
rect 117464 364964 117470 364976
rect 145006 364964 145012 364976
rect 145064 364964 145070 365016
rect 163590 364760 163596 364812
rect 163648 364800 163654 364812
rect 258258 364800 258264 364812
rect 163648 364772 258264 364800
rect 163648 364760 163654 364772
rect 258258 364760 258264 364772
rect 258316 364800 258322 364812
rect 259362 364800 259368 364812
rect 258316 364772 259368 364800
rect 258316 364760 258322 364772
rect 259362 364760 259368 364772
rect 259420 364760 259426 364812
rect 176010 364692 176016 364744
rect 176068 364732 176074 364744
rect 224218 364732 224224 364744
rect 176068 364704 224224 364732
rect 176068 364692 176074 364704
rect 224218 364692 224224 364704
rect 224276 364692 224282 364744
rect 188430 364624 188436 364676
rect 188488 364664 188494 364676
rect 303522 364664 303528 364676
rect 188488 364636 303528 364664
rect 188488 364624 188494 364636
rect 303522 364624 303528 364636
rect 303580 364624 303586 364676
rect 305086 364624 305092 364676
rect 305144 364664 305150 364676
rect 305638 364664 305644 364676
rect 305144 364636 305644 364664
rect 305144 364624 305150 364636
rect 305638 364624 305644 364636
rect 305696 364664 305702 364676
rect 342346 364664 342352 364676
rect 305696 364636 342352 364664
rect 305696 364624 305702 364636
rect 342346 364624 342352 364636
rect 342404 364624 342410 364676
rect 123662 364556 123668 364608
rect 123720 364596 123726 364608
rect 214834 364596 214840 364608
rect 123720 364568 214840 364596
rect 123720 364556 123726 364568
rect 214834 364556 214840 364568
rect 214892 364596 214898 364608
rect 343634 364596 343640 364608
rect 214892 364568 343640 364596
rect 214892 364556 214898 364568
rect 343634 364556 343640 364568
rect 343692 364556 343698 364608
rect 146938 364488 146944 364540
rect 146996 364528 147002 364540
rect 324406 364528 324412 364540
rect 146996 364500 324412 364528
rect 146996 364488 147002 364500
rect 324406 364488 324412 364500
rect 324464 364488 324470 364540
rect 257338 364420 257344 364472
rect 257396 364460 257402 364472
rect 447778 364460 447784 364472
rect 257396 364432 447784 364460
rect 257396 364420 257402 364432
rect 447778 364420 447784 364432
rect 447836 364420 447842 364472
rect 41230 364352 41236 364404
rect 41288 364392 41294 364404
rect 69014 364392 69020 364404
rect 41288 364364 69020 364392
rect 41288 364352 41294 364364
rect 69014 364352 69020 364364
rect 69072 364352 69078 364404
rect 198642 364352 198648 364404
rect 198700 364392 198706 364404
rect 579798 364392 579804 364404
rect 198700 364364 511994 364392
rect 198700 364352 198706 364364
rect 508516 364336 508544 364364
rect 118142 364284 118148 364336
rect 118200 364324 118206 364336
rect 146386 364324 146392 364336
rect 118200 364296 146392 364324
rect 118200 364284 118206 364296
rect 146386 364284 146392 364296
rect 146444 364284 146450 364336
rect 508498 364284 508504 364336
rect 508556 364284 508562 364336
rect 511966 364256 511994 364364
rect 579586 364364 579804 364392
rect 579586 364336 579614 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 579586 364296 579620 364336
rect 579614 364284 579620 364296
rect 579672 364284 579678 364336
rect 511966 364228 518894 364256
rect 56318 363672 56324 363724
rect 56376 363712 56382 363724
rect 69382 363712 69388 363724
rect 56376 363684 69388 363712
rect 56376 363672 56382 363684
rect 69382 363672 69388 363684
rect 69440 363672 69446 363724
rect 43990 363604 43996 363656
rect 44048 363644 44054 363656
rect 67634 363644 67640 363656
rect 44048 363616 67640 363644
rect 44048 363604 44054 363616
rect 67634 363604 67640 363616
rect 67692 363604 67698 363656
rect 518866 363644 518894 364228
rect 579614 363644 579620 363656
rect 518866 363616 579620 363644
rect 579614 363604 579620 363616
rect 579672 363604 579678 363656
rect 195238 363264 195244 363316
rect 195296 363304 195302 363316
rect 206462 363304 206468 363316
rect 195296 363276 206468 363304
rect 195296 363264 195302 363276
rect 206462 363264 206468 363276
rect 206520 363264 206526 363316
rect 187050 363196 187056 363248
rect 187108 363236 187114 363248
rect 233878 363236 233884 363248
rect 187108 363208 233884 363236
rect 187108 363196 187114 363208
rect 233878 363196 233884 363208
rect 233936 363196 233942 363248
rect 242158 363196 242164 363248
rect 242216 363236 242222 363248
rect 242526 363236 242532 363248
rect 242216 363208 242532 363236
rect 242216 363196 242222 363208
rect 242526 363196 242532 363208
rect 242584 363236 242590 363248
rect 323302 363236 323308 363248
rect 242584 363208 323308 363236
rect 242584 363196 242590 363208
rect 323302 363196 323308 363208
rect 323360 363196 323366 363248
rect 195330 363128 195336 363180
rect 195388 363168 195394 363180
rect 285030 363168 285036 363180
rect 195388 363140 285036 363168
rect 195388 363128 195394 363140
rect 285030 363128 285036 363140
rect 285088 363128 285094 363180
rect 301498 363128 301504 363180
rect 301556 363168 301562 363180
rect 413278 363168 413284 363180
rect 301556 363140 413284 363168
rect 301556 363128 301562 363140
rect 413278 363128 413284 363140
rect 413336 363128 413342 363180
rect 178862 363060 178868 363112
rect 178920 363100 178926 363112
rect 236086 363100 236092 363112
rect 178920 363072 236092 363100
rect 178920 363060 178926 363072
rect 236086 363060 236092 363072
rect 236144 363100 236150 363112
rect 356054 363100 356060 363112
rect 236144 363072 356060 363100
rect 236144 363060 236150 363072
rect 356054 363060 356060 363072
rect 356112 363060 356118 363112
rect 196618 362992 196624 363044
rect 196676 363032 196682 363044
rect 322106 363032 322112 363044
rect 196676 363004 322112 363032
rect 196676 362992 196682 363004
rect 322106 362992 322112 363004
rect 322164 362992 322170 363044
rect 164878 362924 164884 362976
rect 164936 362964 164942 362976
rect 247034 362964 247040 362976
rect 164936 362936 247040 362964
rect 164936 362924 164942 362936
rect 247034 362924 247040 362936
rect 247092 362964 247098 362976
rect 247092 362936 248414 362964
rect 247092 362924 247098 362936
rect 118602 362856 118608 362908
rect 118660 362896 118666 362908
rect 140958 362896 140964 362908
rect 118660 362868 140964 362896
rect 118660 362856 118666 362868
rect 140958 362856 140964 362868
rect 141016 362856 141022 362908
rect 248386 362896 248414 362936
rect 268378 362924 268384 362976
rect 268436 362964 268442 362976
rect 466454 362964 466460 362976
rect 268436 362936 466460 362964
rect 268436 362924 268442 362936
rect 466454 362924 466460 362936
rect 466512 362924 466518 362976
rect 304994 362896 305000 362908
rect 248386 362868 305000 362896
rect 304994 362856 305000 362868
rect 305052 362856 305058 362908
rect 226978 362448 226984 362500
rect 227036 362488 227042 362500
rect 229646 362488 229652 362500
rect 227036 362460 229652 362488
rect 227036 362448 227042 362460
rect 229646 362448 229652 362460
rect 229704 362448 229710 362500
rect 199562 362244 199568 362296
rect 199620 362284 199626 362296
rect 223482 362284 223488 362296
rect 199620 362256 223488 362284
rect 199620 362244 199626 362256
rect 223482 362244 223488 362256
rect 223540 362244 223546 362296
rect 140958 362176 140964 362228
rect 141016 362216 141022 362228
rect 180150 362216 180156 362228
rect 141016 362188 180156 362216
rect 141016 362176 141022 362188
rect 180150 362176 180156 362188
rect 180208 362176 180214 362228
rect 196710 362176 196716 362228
rect 196768 362216 196774 362228
rect 249702 362216 249708 362228
rect 196768 362188 249708 362216
rect 196768 362176 196774 362188
rect 249702 362176 249708 362188
rect 249760 362216 249766 362228
rect 250898 362216 250904 362228
rect 249760 362188 250904 362216
rect 249760 362176 249766 362188
rect 250898 362176 250904 362188
rect 250956 362176 250962 362228
rect 313274 362176 313280 362228
rect 313332 362216 313338 362228
rect 406378 362216 406384 362228
rect 313332 362188 406384 362216
rect 313332 362176 313338 362188
rect 406378 362176 406384 362188
rect 406436 362176 406442 362228
rect 310790 361972 310796 362024
rect 310848 362012 310854 362024
rect 313274 362012 313280 362024
rect 310848 361984 313280 362012
rect 310848 361972 310854 361984
rect 313274 361972 313280 361984
rect 313332 361972 313338 362024
rect 258258 361904 258264 361956
rect 258316 361944 258322 361956
rect 259914 361944 259920 361956
rect 258316 361916 259920 361944
rect 258316 361904 258322 361916
rect 259914 361904 259920 361916
rect 259972 361904 259978 361956
rect 274726 361904 274732 361956
rect 274784 361944 274790 361956
rect 275922 361944 275928 361956
rect 274784 361916 275928 361944
rect 274784 361904 274790 361916
rect 275922 361904 275928 361916
rect 275980 361944 275986 361956
rect 514754 361944 514760 361956
rect 275980 361916 514760 361944
rect 275980 361904 275986 361916
rect 514754 361904 514760 361916
rect 514812 361904 514818 361956
rect 240594 361876 240600 361888
rect 122806 361848 240600 361876
rect 118602 361768 118608 361820
rect 118660 361808 118666 361820
rect 120074 361808 120080 361820
rect 118660 361780 120080 361808
rect 118660 361768 118666 361780
rect 120074 361768 120080 361780
rect 120132 361808 120138 361820
rect 122806 361808 122834 361848
rect 240594 361836 240600 361848
rect 240652 361836 240658 361888
rect 289538 361836 289544 361888
rect 289596 361876 289602 361888
rect 300762 361876 300768 361888
rect 289596 361848 300768 361876
rect 289596 361836 289602 361848
rect 300762 361836 300768 361848
rect 300820 361836 300826 361888
rect 120132 361780 122834 361808
rect 120132 361768 120138 361780
rect 193490 361768 193496 361820
rect 193548 361808 193554 361820
rect 204530 361808 204536 361820
rect 193548 361780 204536 361808
rect 193548 361768 193554 361780
rect 204530 361768 204536 361780
rect 204588 361768 204594 361820
rect 221274 361768 221280 361820
rect 221332 361808 221338 361820
rect 222838 361808 222844 361820
rect 221332 361780 222844 361808
rect 221332 361768 221338 361780
rect 222838 361768 222844 361780
rect 222896 361768 222902 361820
rect 224218 361768 224224 361820
rect 224276 361808 224282 361820
rect 225782 361808 225788 361820
rect 224276 361780 225788 361808
rect 224276 361768 224282 361780
rect 225782 361768 225788 361780
rect 225840 361768 225846 361820
rect 278130 361768 278136 361820
rect 278188 361808 278194 361820
rect 278590 361808 278596 361820
rect 278188 361780 278596 361808
rect 278188 361768 278194 361780
rect 278590 361768 278596 361780
rect 278648 361808 278654 361820
rect 320818 361808 320824 361820
rect 278648 361780 320824 361808
rect 278648 361768 278654 361780
rect 320818 361768 320824 361780
rect 320876 361768 320882 361820
rect 160830 361700 160836 361752
rect 160888 361740 160894 361752
rect 202598 361740 202604 361752
rect 160888 361712 202604 361740
rect 160888 361700 160894 361712
rect 202598 361700 202604 361712
rect 202656 361700 202662 361752
rect 249702 361700 249708 361752
rect 249760 361740 249766 361752
rect 316862 361740 316868 361752
rect 249760 361712 316868 361740
rect 249760 361700 249766 361712
rect 316862 361700 316868 361712
rect 316920 361700 316926 361752
rect 196802 361632 196808 361684
rect 196860 361672 196866 361684
rect 276658 361672 276664 361684
rect 196860 361644 276664 361672
rect 196860 361632 196866 361644
rect 276658 361632 276664 361644
rect 276716 361632 276722 361684
rect 281166 361672 281172 361684
rect 277366 361644 281172 361672
rect 252462 361564 252468 361616
rect 252520 361604 252526 361616
rect 277366 361604 277394 361644
rect 281166 361632 281172 361644
rect 281224 361672 281230 361684
rect 485038 361672 485044 361684
rect 281224 361644 485044 361672
rect 281224 361632 281230 361644
rect 485038 361632 485044 361644
rect 485096 361632 485102 361684
rect 252520 361576 277394 361604
rect 252520 361564 252526 361576
rect 303522 361564 303528 361616
rect 303580 361604 303586 361616
rect 304350 361604 304356 361616
rect 303580 361576 304356 361604
rect 303580 361564 303586 361576
rect 304350 361564 304356 361576
rect 304408 361564 304414 361616
rect 36998 361496 37004 361548
rect 37056 361536 37062 361548
rect 68002 361536 68008 361548
rect 37056 361508 68008 361536
rect 37056 361496 37062 361508
rect 68002 361496 68008 361508
rect 68060 361496 68066 361548
rect 130010 361496 130016 361548
rect 130068 361536 130074 361548
rect 289538 361536 289544 361548
rect 130068 361508 289544 361536
rect 130068 361496 130074 361508
rect 289538 361496 289544 361508
rect 289596 361496 289602 361548
rect 45462 361428 45468 361480
rect 45520 361468 45526 361480
rect 66990 361468 66996 361480
rect 45520 361440 66996 361468
rect 45520 361428 45526 361440
rect 66990 361428 66996 361440
rect 67048 361468 67054 361480
rect 67542 361468 67548 361480
rect 67048 361440 67548 361468
rect 67048 361428 67054 361440
rect 67542 361428 67548 361440
rect 67600 361428 67606 361480
rect 118050 361428 118056 361480
rect 118108 361468 118114 361480
rect 147858 361468 147864 361480
rect 118108 361440 147864 361468
rect 118108 361428 118114 361440
rect 147858 361428 147864 361440
rect 147916 361468 147922 361480
rect 252462 361468 252468 361480
rect 147916 361440 252468 361468
rect 147916 361428 147922 361440
rect 252462 361428 252468 361440
rect 252520 361428 252526 361480
rect 146478 361360 146484 361412
rect 146536 361400 146542 361412
rect 200758 361400 200764 361412
rect 146536 361372 200764 361400
rect 146536 361360 146542 361372
rect 200758 361360 200764 361372
rect 200816 361360 200822 361412
rect 119522 360952 119528 361004
rect 119580 360992 119586 361004
rect 120258 360992 120264 361004
rect 119580 360964 120264 360992
rect 119580 360952 119586 360964
rect 120258 360952 120264 360964
rect 120316 360992 120322 361004
rect 120316 360964 122834 360992
rect 120316 360952 120322 360964
rect 64782 360816 64788 360868
rect 64840 360856 64846 360868
rect 67634 360856 67640 360868
rect 64840 360828 67640 360856
rect 64840 360816 64846 360828
rect 67634 360816 67640 360828
rect 67692 360816 67698 360868
rect 122806 360856 122834 360964
rect 198182 360884 198188 360936
rect 198240 360924 198246 360936
rect 216582 360924 216588 360936
rect 198240 360896 216588 360924
rect 198240 360884 198246 360896
rect 216582 360884 216588 360896
rect 216640 360924 216646 360936
rect 217134 360924 217140 360936
rect 216640 360896 217140 360924
rect 216640 360884 216646 360896
rect 217134 360884 217140 360896
rect 217192 360884 217198 360936
rect 300762 360884 300768 360936
rect 300820 360924 300826 360936
rect 452654 360924 452660 360936
rect 300820 360896 452660 360924
rect 300820 360884 300826 360896
rect 452654 360884 452660 360896
rect 452712 360884 452718 360936
rect 314654 360856 314660 360868
rect 122806 360828 314660 360856
rect 314654 360816 314660 360828
rect 314712 360816 314718 360868
rect 312538 360408 312544 360460
rect 312596 360448 312602 360460
rect 323026 360448 323032 360460
rect 312596 360420 323032 360448
rect 312596 360408 312602 360420
rect 323026 360408 323032 360420
rect 323084 360408 323090 360460
rect 285030 360340 285036 360392
rect 285088 360380 285094 360392
rect 319438 360380 319444 360392
rect 285088 360352 319444 360380
rect 285088 360340 285094 360352
rect 319438 360340 319444 360352
rect 319496 360340 319502 360392
rect 145558 360272 145564 360324
rect 145616 360312 145622 360324
rect 146478 360312 146484 360324
rect 145616 360284 146484 360312
rect 145616 360272 145622 360284
rect 146478 360272 146484 360284
rect 146536 360272 146542 360324
rect 308214 360272 308220 360324
rect 308272 360312 308278 360324
rect 308398 360312 308404 360324
rect 308272 360284 308404 360312
rect 308272 360272 308278 360284
rect 308398 360272 308404 360284
rect 308456 360312 308462 360324
rect 359458 360312 359464 360324
rect 308456 360284 359464 360312
rect 308456 360272 308462 360284
rect 359458 360272 359464 360284
rect 359516 360272 359522 360324
rect 129090 360204 129096 360256
rect 129148 360244 129154 360256
rect 130010 360244 130016 360256
rect 129148 360216 130016 360244
rect 129148 360204 129154 360216
rect 130010 360204 130016 360216
rect 130068 360204 130074 360256
rect 196894 360204 196900 360256
rect 196952 360244 196958 360256
rect 257338 360244 257344 360256
rect 196952 360216 257344 360244
rect 196952 360204 196958 360216
rect 257338 360204 257344 360216
rect 257396 360204 257402 360256
rect 272150 360204 272156 360256
rect 272208 360244 272214 360256
rect 389818 360244 389824 360256
rect 272208 360216 389824 360244
rect 272208 360204 272214 360216
rect 389818 360204 389824 360216
rect 389876 360204 389882 360256
rect 118510 360136 118516 360188
rect 118568 360176 118574 360188
rect 149146 360176 149152 360188
rect 118568 360148 149152 360176
rect 118568 360136 118574 360148
rect 149146 360136 149152 360148
rect 149204 360176 149210 360188
rect 149698 360176 149704 360188
rect 149204 360148 149704 360176
rect 149204 360136 149210 360148
rect 149698 360136 149704 360148
rect 149756 360136 149762 360188
rect 118602 360068 118608 360120
rect 118660 360108 118666 360120
rect 133782 360108 133788 360120
rect 118660 360080 133788 360108
rect 118660 360068 118666 360080
rect 133782 360068 133788 360080
rect 133840 360068 133846 360120
rect 39758 359456 39764 359508
rect 39816 359496 39822 359508
rect 67634 359496 67640 359508
rect 39816 359468 67640 359496
rect 39816 359456 39822 359468
rect 67634 359456 67640 359468
rect 67692 359456 67698 359508
rect 68554 359456 68560 359508
rect 68612 359496 68618 359508
rect 68922 359496 68928 359508
rect 68612 359468 68928 359496
rect 68612 359456 68618 359468
rect 68922 359456 68928 359468
rect 68980 359456 68986 359508
rect 133782 359456 133788 359508
rect 133840 359496 133846 359508
rect 143718 359496 143724 359508
rect 133840 359468 143724 359496
rect 133840 359456 133846 359468
rect 143718 359456 143724 359468
rect 143776 359456 143782 359508
rect 317506 359456 317512 359508
rect 317564 359496 317570 359508
rect 319622 359496 319628 359508
rect 317564 359468 319628 359496
rect 317564 359456 317570 359468
rect 319622 359456 319628 359468
rect 319680 359456 319686 359508
rect 193858 358912 193864 358964
rect 193916 358952 193922 358964
rect 321554 358952 321560 358964
rect 193916 358924 321560 358952
rect 193916 358912 193922 358924
rect 321554 358912 321560 358924
rect 321612 358912 321618 358964
rect 169110 358844 169116 358896
rect 169168 358884 169174 358896
rect 324590 358884 324596 358896
rect 169168 358856 324596 358884
rect 169168 358844 169174 358856
rect 324590 358844 324596 358856
rect 324648 358844 324654 358896
rect 158162 358776 158168 358828
rect 158220 358816 158226 358828
rect 320358 358816 320364 358828
rect 158220 358788 320364 358816
rect 158220 358776 158226 358788
rect 320358 358776 320364 358788
rect 320416 358776 320422 358828
rect 64138 358708 64144 358760
rect 64196 358748 64202 358760
rect 67450 358748 67456 358760
rect 64196 358720 67456 358748
rect 64196 358708 64202 358720
rect 67450 358708 67456 358720
rect 67508 358748 67514 358760
rect 67634 358748 67640 358760
rect 67508 358720 67640 358748
rect 67508 358708 67514 358720
rect 67634 358708 67640 358720
rect 67692 358708 67698 358760
rect 122650 358096 122656 358148
rect 122708 358136 122714 358148
rect 146386 358136 146392 358148
rect 122708 358108 146392 358136
rect 122708 358096 122714 358108
rect 146386 358096 146392 358108
rect 146444 358096 146450 358148
rect 53558 358028 53564 358080
rect 53616 358068 53622 358080
rect 67634 358068 67640 358080
rect 53616 358040 67640 358068
rect 53616 358028 53622 358040
rect 67634 358028 67640 358040
rect 67692 358028 67698 358080
rect 118602 358028 118608 358080
rect 118660 358068 118666 358080
rect 120718 358068 120724 358080
rect 118660 358040 120724 358068
rect 118660 358028 118666 358040
rect 120718 358028 120724 358040
rect 120776 358068 120782 358080
rect 148318 358068 148324 358080
rect 120776 358040 148324 358068
rect 120776 358028 120782 358040
rect 148318 358028 148324 358040
rect 148376 358068 148382 358080
rect 193490 358068 193496 358080
rect 148376 358040 193496 358068
rect 148376 358028 148382 358040
rect 193490 358028 193496 358040
rect 193548 358028 193554 358080
rect 3418 357824 3424 357876
rect 3476 357864 3482 357876
rect 7558 357864 7564 357876
rect 3476 357836 7564 357864
rect 3476 357824 3482 357836
rect 7558 357824 7564 357836
rect 7616 357824 7622 357876
rect 146386 357416 146392 357468
rect 146444 357456 146450 357468
rect 198090 357456 198096 357468
rect 146444 357428 198096 357456
rect 146444 357416 146450 357428
rect 198090 357416 198096 357428
rect 198148 357416 198154 357468
rect 118602 357348 118608 357400
rect 118660 357388 118666 357400
rect 144914 357388 144920 357400
rect 118660 357360 144920 357388
rect 118660 357348 118666 357360
rect 144914 357348 144920 357360
rect 144972 357388 144978 357400
rect 146202 357388 146208 357400
rect 144972 357360 146208 357388
rect 144972 357348 144978 357360
rect 146202 357348 146208 357360
rect 146260 357348 146266 357400
rect 198734 356940 198740 356992
rect 198792 356980 198798 356992
rect 199654 356980 199660 356992
rect 198792 356952 199660 356980
rect 198792 356940 198798 356952
rect 199654 356940 199660 356952
rect 199712 356940 199718 356992
rect 118602 356668 118608 356720
rect 118660 356708 118666 356720
rect 142430 356708 142436 356720
rect 118660 356680 142436 356708
rect 118660 356668 118666 356680
rect 142430 356668 142436 356680
rect 142488 356708 142494 356720
rect 142798 356708 142804 356720
rect 142488 356680 142804 356708
rect 142488 356668 142494 356680
rect 142798 356668 142804 356680
rect 142856 356668 142862 356720
rect 151078 356668 151084 356720
rect 151136 356708 151142 356720
rect 193950 356708 193956 356720
rect 151136 356680 193956 356708
rect 151136 356668 151142 356680
rect 193950 356668 193956 356680
rect 194008 356668 194014 356720
rect 191098 356192 191104 356244
rect 191156 356232 191162 356244
rect 197354 356232 197360 356244
rect 191156 356204 197360 356232
rect 191156 356192 191162 356204
rect 197354 356192 197360 356204
rect 197412 356192 197418 356244
rect 42610 356056 42616 356108
rect 42668 356096 42674 356108
rect 67910 356096 67916 356108
rect 42668 356068 67916 356096
rect 42668 356056 42674 356068
rect 67910 356056 67916 356068
rect 67968 356056 67974 356108
rect 57790 355376 57796 355428
rect 57848 355416 57854 355428
rect 67634 355416 67640 355428
rect 57848 355388 67640 355416
rect 57848 355376 57854 355388
rect 67634 355376 67640 355388
rect 67692 355376 67698 355428
rect 52178 355308 52184 355360
rect 52236 355348 52242 355360
rect 54202 355348 54208 355360
rect 52236 355320 54208 355348
rect 52236 355308 52242 355320
rect 54202 355308 54208 355320
rect 54260 355348 54266 355360
rect 67726 355348 67732 355360
rect 54260 355320 67732 355348
rect 54260 355308 54266 355320
rect 67726 355308 67732 355320
rect 67784 355308 67790 355360
rect 118142 354696 118148 354748
rect 118200 354736 118206 354748
rect 182818 354736 182824 354748
rect 118200 354708 182824 354736
rect 118200 354696 118206 354708
rect 182818 354696 182824 354708
rect 182876 354696 182882 354748
rect 117774 354628 117780 354680
rect 117832 354668 117838 354680
rect 128630 354668 128636 354680
rect 117832 354640 128636 354668
rect 117832 354628 117838 354640
rect 128630 354628 128636 354640
rect 128688 354628 128694 354680
rect 128630 354016 128636 354068
rect 128688 354056 128694 354068
rect 128688 354028 142154 354056
rect 128688 354016 128694 354028
rect 142126 354000 142154 354028
rect 115934 353948 115940 354000
rect 115992 353988 115998 354000
rect 137278 353988 137284 354000
rect 115992 353960 137284 353988
rect 115992 353948 115998 353960
rect 137278 353948 137284 353960
rect 137336 353948 137342 354000
rect 142126 353960 142160 354000
rect 142154 353948 142160 353960
rect 142212 353988 142218 354000
rect 198182 353988 198188 354000
rect 142212 353960 198188 353988
rect 142212 353948 142218 353960
rect 198182 353948 198188 353960
rect 198240 353948 198246 354000
rect 49602 352588 49608 352640
rect 49660 352628 49666 352640
rect 68554 352628 68560 352640
rect 49660 352600 68560 352628
rect 49660 352588 49666 352600
rect 68554 352588 68560 352600
rect 68612 352588 68618 352640
rect 33042 352520 33048 352572
rect 33100 352560 33106 352572
rect 63494 352560 63500 352572
rect 33100 352532 63500 352560
rect 33100 352520 33106 352532
rect 63494 352520 63500 352532
rect 63552 352520 63558 352572
rect 118602 352520 118608 352572
rect 118660 352560 118666 352572
rect 118660 352532 142154 352560
rect 118660 352520 118666 352532
rect 142126 352492 142154 352532
rect 144914 352492 144920 352504
rect 142126 352464 144920 352492
rect 144914 352452 144920 352464
rect 144972 352492 144978 352504
rect 145558 352492 145564 352504
rect 144972 352464 145564 352492
rect 144972 352452 144978 352464
rect 145558 352452 145564 352464
rect 145616 352452 145622 352504
rect 15838 351908 15844 351960
rect 15896 351948 15902 351960
rect 49418 351948 49424 351960
rect 15896 351920 49424 351948
rect 15896 351908 15902 351920
rect 49418 351908 49424 351920
rect 49476 351948 49482 351960
rect 49602 351948 49608 351960
rect 49476 351920 49608 351948
rect 49476 351908 49482 351920
rect 49602 351908 49608 351920
rect 49660 351908 49666 351960
rect 63494 351908 63500 351960
rect 63552 351948 63558 351960
rect 64414 351948 64420 351960
rect 63552 351920 64420 351948
rect 63552 351908 63558 351920
rect 64414 351908 64420 351920
rect 64472 351948 64478 351960
rect 67634 351948 67640 351960
rect 64472 351920 67640 351948
rect 64472 351908 64478 351920
rect 67634 351908 67640 351920
rect 67692 351908 67698 351960
rect 118050 351840 118056 351892
rect 118108 351880 118114 351892
rect 147766 351880 147772 351892
rect 118108 351852 147772 351880
rect 118108 351840 118114 351852
rect 147766 351840 147772 351852
rect 147824 351840 147830 351892
rect 118602 351160 118608 351212
rect 118660 351200 118666 351212
rect 170398 351200 170404 351212
rect 118660 351172 170404 351200
rect 118660 351160 118666 351172
rect 170398 351160 170404 351172
rect 170456 351160 170462 351212
rect 177298 351160 177304 351212
rect 177356 351200 177362 351212
rect 198734 351200 198740 351212
rect 177356 351172 198740 351200
rect 177356 351160 177362 351172
rect 198734 351160 198740 351172
rect 198792 351160 198798 351212
rect 322106 351160 322112 351212
rect 322164 351200 322170 351212
rect 360838 351200 360844 351212
rect 322164 351172 360844 351200
rect 322164 351160 322170 351172
rect 360838 351160 360844 351172
rect 360896 351160 360902 351212
rect 504358 351160 504364 351212
rect 504416 351200 504422 351212
rect 580166 351200 580172 351212
rect 504416 351172 580172 351200
rect 504416 351160 504422 351172
rect 580166 351160 580172 351172
rect 580224 351160 580230 351212
rect 60458 350548 60464 350600
rect 60516 350588 60522 350600
rect 61838 350588 61844 350600
rect 60516 350560 61844 350588
rect 60516 350548 60522 350560
rect 61838 350548 61844 350560
rect 61896 350588 61902 350600
rect 67634 350588 67640 350600
rect 61896 350560 67640 350588
rect 61896 350548 61902 350560
rect 67634 350548 67640 350560
rect 67692 350548 67698 350600
rect 118602 350276 118608 350328
rect 118660 350316 118666 350328
rect 124214 350316 124220 350328
rect 118660 350288 124220 350316
rect 118660 350276 118666 350288
rect 124214 350276 124220 350288
rect 124272 350276 124278 350328
rect 117958 349800 117964 349852
rect 118016 349840 118022 349852
rect 118694 349840 118700 349852
rect 118016 349812 118700 349840
rect 118016 349800 118022 349812
rect 118694 349800 118700 349812
rect 118752 349800 118758 349852
rect 322750 349800 322756 349852
rect 322808 349840 322814 349852
rect 323210 349840 323216 349852
rect 322808 349812 323216 349840
rect 322808 349800 322814 349812
rect 323210 349800 323216 349812
rect 323268 349840 323274 349852
rect 489178 349840 489184 349852
rect 323268 349812 489184 349840
rect 323268 349800 323274 349812
rect 489178 349800 489184 349812
rect 489236 349800 489242 349852
rect 46566 349188 46572 349240
rect 46624 349228 46630 349240
rect 68002 349228 68008 349240
rect 46624 349200 68008 349228
rect 46624 349188 46630 349200
rect 68002 349188 68008 349200
rect 68060 349188 68066 349240
rect 35802 349120 35808 349172
rect 35860 349160 35866 349172
rect 62114 349160 62120 349172
rect 35860 349132 62120 349160
rect 35860 349120 35866 349132
rect 62114 349120 62120 349132
rect 62172 349120 62178 349172
rect 62132 349092 62160 349120
rect 67634 349092 67640 349104
rect 62132 349064 67640 349092
rect 67634 349052 67640 349064
rect 67692 349052 67698 349104
rect 118602 349052 118608 349104
rect 118660 349092 118666 349104
rect 151814 349092 151820 349104
rect 118660 349064 151820 349092
rect 118660 349052 118666 349064
rect 151814 349052 151820 349064
rect 151872 349092 151878 349104
rect 153102 349092 153108 349104
rect 151872 349064 153108 349092
rect 151872 349052 151878 349064
rect 153102 349052 153108 349064
rect 153160 349052 153166 349104
rect 117682 348984 117688 349036
rect 117740 349024 117746 349036
rect 151998 349024 152004 349036
rect 117740 348996 152004 349024
rect 117740 348984 117746 348996
rect 151998 348984 152004 348996
rect 152056 349024 152062 349036
rect 153010 349024 153016 349036
rect 152056 348996 153016 349024
rect 152056 348984 152062 348996
rect 153010 348984 153016 348996
rect 153068 348984 153074 349036
rect 153102 348372 153108 348424
rect 153160 348412 153166 348424
rect 188338 348412 188344 348424
rect 153160 348384 188344 348412
rect 153160 348372 153166 348384
rect 188338 348372 188344 348384
rect 188396 348372 188402 348424
rect 320818 348372 320824 348424
rect 320876 348412 320882 348424
rect 448514 348412 448520 348424
rect 320876 348384 448520 348412
rect 320876 348372 320882 348384
rect 448514 348372 448520 348384
rect 448572 348372 448578 348424
rect 65518 347692 65524 347744
rect 65576 347732 65582 347744
rect 66070 347732 66076 347744
rect 65576 347704 66076 347732
rect 65576 347692 65582 347704
rect 66070 347692 66076 347704
rect 66128 347692 66134 347744
rect 117406 347692 117412 347744
rect 117464 347732 117470 347744
rect 132494 347732 132500 347744
rect 117464 347704 132500 347732
rect 117464 347692 117470 347704
rect 132494 347692 132500 347704
rect 132552 347732 132558 347744
rect 133782 347732 133788 347744
rect 132552 347704 133788 347732
rect 132552 347692 132558 347704
rect 133782 347692 133788 347704
rect 133840 347692 133846 347744
rect 133782 347012 133788 347064
rect 133840 347052 133846 347064
rect 180058 347052 180064 347064
rect 133840 347024 180064 347052
rect 133840 347012 133846 347024
rect 180058 347012 180064 347024
rect 180116 347012 180122 347064
rect 319622 347012 319628 347064
rect 319680 347052 319686 347064
rect 469214 347052 469220 347064
rect 319680 347024 469220 347052
rect 319680 347012 319686 347024
rect 469214 347012 469220 347024
rect 469272 347012 469278 347064
rect 66070 346944 66076 346996
rect 66128 346984 66134 346996
rect 67634 346984 67640 346996
rect 66128 346956 67640 346984
rect 66128 346944 66134 346956
rect 67634 346944 67640 346956
rect 67692 346944 67698 346996
rect 183002 346400 183008 346452
rect 183060 346440 183066 346452
rect 197354 346440 197360 346452
rect 183060 346412 197360 346440
rect 183060 346400 183066 346412
rect 197354 346400 197360 346412
rect 197412 346400 197418 346452
rect 7558 346332 7564 346384
rect 7616 346372 7622 346384
rect 68554 346372 68560 346384
rect 7616 346344 68560 346372
rect 7616 346332 7622 346344
rect 68554 346332 68560 346344
rect 68612 346372 68618 346384
rect 68830 346372 68836 346384
rect 68612 346344 68836 346372
rect 68612 346332 68618 346344
rect 68830 346332 68836 346344
rect 68888 346332 68894 346384
rect 118602 346332 118608 346384
rect 118660 346372 118666 346384
rect 142246 346372 142252 346384
rect 118660 346344 142252 346372
rect 118660 346332 118666 346344
rect 142246 346332 142252 346344
rect 142304 346372 142310 346384
rect 143442 346372 143448 346384
rect 142304 346344 143448 346372
rect 142304 346332 142310 346344
rect 143442 346332 143448 346344
rect 143500 346332 143506 346384
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 143626 345692 143632 345704
rect 122806 345664 143632 345692
rect 118510 345584 118516 345636
rect 118568 345624 118574 345636
rect 119706 345624 119712 345636
rect 118568 345596 119712 345624
rect 118568 345584 118574 345596
rect 119706 345584 119712 345596
rect 119764 345624 119770 345636
rect 122806 345624 122834 345664
rect 143626 345652 143632 345664
rect 143684 345692 143690 345704
rect 144270 345692 144276 345704
rect 143684 345664 144276 345692
rect 143684 345652 143690 345664
rect 144270 345652 144276 345664
rect 144328 345652 144334 345704
rect 322474 345652 322480 345704
rect 322532 345692 322538 345704
rect 327074 345692 327080 345704
rect 322532 345664 327080 345692
rect 322532 345652 322538 345664
rect 327074 345652 327080 345664
rect 327132 345692 327138 345704
rect 461578 345692 461584 345704
rect 327132 345664 461584 345692
rect 327132 345652 327138 345664
rect 461578 345652 461584 345664
rect 461636 345652 461642 345704
rect 119764 345596 122834 345624
rect 119764 345584 119770 345596
rect 43898 345040 43904 345092
rect 43956 345080 43962 345092
rect 68646 345080 68652 345092
rect 43956 345052 68652 345080
rect 43956 345040 43962 345052
rect 68646 345040 68652 345052
rect 68704 345040 68710 345092
rect 118602 344972 118608 345024
rect 118660 345012 118666 345024
rect 138106 345012 138112 345024
rect 118660 344984 138112 345012
rect 118660 344972 118666 344984
rect 138106 344972 138112 344984
rect 138164 344972 138170 345024
rect 46842 344292 46848 344344
rect 46900 344332 46906 344344
rect 58986 344332 58992 344344
rect 46900 344304 58992 344332
rect 46900 344292 46906 344304
rect 58986 344292 58992 344304
rect 59044 344292 59050 344344
rect 138106 344292 138112 344344
rect 138164 344332 138170 344344
rect 186958 344332 186964 344344
rect 138164 344304 186964 344332
rect 138164 344292 138170 344304
rect 186958 344292 186964 344304
rect 187016 344292 187022 344344
rect 321646 344292 321652 344344
rect 321704 344332 321710 344344
rect 328454 344332 328460 344344
rect 321704 344304 328460 344332
rect 321704 344292 321710 344304
rect 328454 344292 328460 344304
rect 328512 344292 328518 344344
rect 58986 343680 58992 343732
rect 59044 343720 59050 343732
rect 67634 343720 67640 343732
rect 59044 343692 67640 343720
rect 59044 343680 59050 343692
rect 67634 343680 67640 343692
rect 67692 343680 67698 343732
rect 41322 343612 41328 343664
rect 41380 343652 41386 343664
rect 62758 343652 62764 343664
rect 41380 343624 62764 343652
rect 41380 343612 41386 343624
rect 62758 343612 62764 343624
rect 62816 343612 62822 343664
rect 62776 343584 62804 343612
rect 67634 343584 67640 343596
rect 62776 343556 67640 343584
rect 67634 343544 67640 343556
rect 67692 343544 67698 343596
rect 117866 343544 117872 343596
rect 117924 343584 117930 343596
rect 150526 343584 150532 343596
rect 117924 343556 150532 343584
rect 117924 343544 117930 343556
rect 150526 343544 150532 343556
rect 150584 343544 150590 343596
rect 117498 342932 117504 342984
rect 117556 342972 117562 342984
rect 126790 342972 126796 342984
rect 117556 342944 126796 342972
rect 117556 342932 117562 342944
rect 126790 342932 126796 342944
rect 126848 342932 126854 342984
rect 117682 342864 117688 342916
rect 117740 342904 117746 342916
rect 127158 342904 127164 342916
rect 117740 342876 127164 342904
rect 117740 342864 117746 342876
rect 127158 342864 127164 342876
rect 127216 342864 127222 342916
rect 322474 342864 322480 342916
rect 322532 342904 322538 342916
rect 327166 342904 327172 342916
rect 322532 342876 327172 342904
rect 322532 342864 322538 342876
rect 327166 342864 327172 342876
rect 327224 342904 327230 342916
rect 465074 342904 465080 342916
rect 327224 342876 465080 342904
rect 327224 342864 327230 342876
rect 465074 342864 465080 342876
rect 465132 342864 465138 342916
rect 34146 342184 34152 342236
rect 34204 342224 34210 342236
rect 68646 342224 68652 342236
rect 34204 342196 68652 342224
rect 34204 342184 34210 342196
rect 68646 342184 68652 342196
rect 68704 342184 68710 342236
rect 118602 342184 118608 342236
rect 118660 342224 118666 342236
rect 147674 342224 147680 342236
rect 118660 342196 147680 342224
rect 118660 342184 118666 342196
rect 147674 342184 147680 342196
rect 147732 342184 147738 342236
rect 328546 342184 328552 342236
rect 328604 342224 328610 342236
rect 370498 342224 370504 342236
rect 328604 342196 370504 342224
rect 328604 342184 328610 342196
rect 370498 342184 370504 342196
rect 370556 342184 370562 342236
rect 147674 341504 147680 341556
rect 147732 341544 147738 341556
rect 178770 341544 178776 341556
rect 147732 341516 178776 341544
rect 147732 341504 147738 341516
rect 178770 341504 178776 341516
rect 178828 341504 178834 341556
rect 322566 341504 322572 341556
rect 322624 341544 322630 341556
rect 322842 341544 322848 341556
rect 322624 341516 322848 341544
rect 322624 341504 322630 341516
rect 322842 341504 322848 341516
rect 322900 341544 322906 341556
rect 328546 341544 328552 341556
rect 322900 341516 328552 341544
rect 322900 341504 322906 341516
rect 328546 341504 328552 341516
rect 328604 341504 328610 341556
rect 61746 340892 61752 340944
rect 61804 340932 61810 340944
rect 63310 340932 63316 340944
rect 61804 340904 63316 340932
rect 61804 340892 61810 340904
rect 63310 340892 63316 340904
rect 63368 340932 63374 340944
rect 67634 340932 67640 340944
rect 63368 340904 67640 340932
rect 63368 340892 63374 340904
rect 67634 340892 67640 340904
rect 67692 340892 67698 340944
rect 117406 340824 117412 340876
rect 117464 340864 117470 340876
rect 138290 340864 138296 340876
rect 117464 340836 138296 340864
rect 117464 340824 117470 340836
rect 138290 340824 138296 340836
rect 138348 340824 138354 340876
rect 117314 340756 117320 340808
rect 117372 340796 117378 340808
rect 129090 340796 129096 340808
rect 117372 340768 129096 340796
rect 117372 340756 117378 340768
rect 129090 340756 129096 340768
rect 129148 340756 129154 340808
rect 43806 340212 43812 340264
rect 43864 340252 43870 340264
rect 43864 340224 64874 340252
rect 43864 340212 43870 340224
rect 64846 339912 64874 340224
rect 122742 340212 122748 340264
rect 122800 340252 122806 340264
rect 150526 340252 150532 340264
rect 122800 340224 150532 340252
rect 122800 340212 122806 340224
rect 150526 340212 150532 340224
rect 150584 340212 150590 340264
rect 69198 340144 69204 340196
rect 69256 340184 69262 340196
rect 132954 340184 132960 340196
rect 69256 340156 132960 340184
rect 69256 340144 69262 340156
rect 132954 340144 132960 340156
rect 133012 340144 133018 340196
rect 427814 340144 427820 340196
rect 427872 340184 427878 340196
rect 497458 340184 497464 340196
rect 427872 340156 497464 340184
rect 427872 340144 427878 340156
rect 497458 340144 497464 340156
rect 497516 340144 497522 340196
rect 73062 339912 73068 339924
rect 64846 339884 73068 339912
rect 73062 339872 73068 339884
rect 73120 339912 73126 339924
rect 73200 339912 73206 339924
rect 73120 339884 73206 339912
rect 73120 339872 73126 339884
rect 73200 339872 73206 339884
rect 73258 339872 73264 339924
rect 37090 339600 37096 339652
rect 37148 339640 37154 339652
rect 70394 339640 70400 339652
rect 37148 339612 70400 339640
rect 37148 339600 37154 339612
rect 70394 339600 70400 339612
rect 70452 339640 70458 339652
rect 71314 339640 71320 339652
rect 70452 339612 71320 339640
rect 70452 339600 70458 339612
rect 71314 339600 71320 339612
rect 71372 339600 71378 339652
rect 59078 339532 59084 339584
rect 59136 339572 59142 339584
rect 70486 339572 70492 339584
rect 59136 339544 70492 339572
rect 59136 339532 59142 339544
rect 70486 339532 70492 339544
rect 70544 339572 70550 339584
rect 70670 339572 70676 339584
rect 70544 339544 70676 339572
rect 70544 339532 70550 339544
rect 70670 339532 70676 339544
rect 70728 339532 70734 339584
rect 64506 339464 64512 339516
rect 64564 339504 64570 339516
rect 67174 339504 67180 339516
rect 64564 339476 67180 339504
rect 64564 339464 64570 339476
rect 67174 339464 67180 339476
rect 67232 339504 67238 339516
rect 67634 339504 67640 339516
rect 67232 339476 67640 339504
rect 67232 339464 67238 339476
rect 67634 339464 67640 339476
rect 67692 339464 67698 339516
rect 106918 339464 106924 339516
rect 106976 339504 106982 339516
rect 117314 339504 117320 339516
rect 106976 339476 117320 339504
rect 106976 339464 106982 339476
rect 117314 339464 117320 339476
rect 117372 339464 117378 339516
rect 132494 339464 132500 339516
rect 132552 339504 132558 339516
rect 132954 339504 132960 339516
rect 132552 339476 132960 339504
rect 132552 339464 132558 339476
rect 132954 339464 132960 339476
rect 133012 339504 133018 339516
rect 169662 339504 169668 339516
rect 133012 339476 169668 339504
rect 133012 339464 133018 339476
rect 169662 339464 169668 339476
rect 169720 339504 169726 339516
rect 197354 339504 197360 339516
rect 169720 339476 197360 339504
rect 169720 339464 169726 339476
rect 197354 339464 197360 339476
rect 197412 339464 197418 339516
rect 322382 339464 322388 339516
rect 322440 339504 322446 339516
rect 332870 339504 332876 339516
rect 322440 339476 332876 339504
rect 322440 339464 322446 339476
rect 332870 339464 332876 339476
rect 332928 339464 332934 339516
rect 113174 339396 113180 339448
rect 113232 339436 113238 339448
rect 113910 339436 113916 339448
rect 113232 339408 113916 339436
rect 113232 339396 113238 339408
rect 113910 339396 113916 339408
rect 113968 339436 113974 339448
rect 119338 339436 119344 339448
rect 113968 339408 119344 339436
rect 113968 339396 113974 339408
rect 119338 339396 119344 339408
rect 119396 339396 119402 339448
rect 55858 339328 55864 339380
rect 55916 339368 55922 339380
rect 73890 339368 73896 339380
rect 55916 339340 73896 339368
rect 55916 339328 55922 339340
rect 73890 339328 73896 339340
rect 73948 339328 73954 339380
rect 87414 339328 87420 339380
rect 87472 339368 87478 339380
rect 87598 339368 87604 339380
rect 87472 339340 87604 339368
rect 87472 339328 87478 339340
rect 87598 339328 87604 339340
rect 87656 339368 87662 339380
rect 191098 339368 191104 339380
rect 87656 339340 191104 339368
rect 87656 339328 87662 339340
rect 191098 339328 191104 339340
rect 191156 339328 191162 339380
rect 54846 339260 54852 339312
rect 54904 339300 54910 339312
rect 79686 339300 79692 339312
rect 54904 339272 79692 339300
rect 54904 339260 54910 339272
rect 79686 339260 79692 339272
rect 79744 339260 79750 339312
rect 104802 339260 104808 339312
rect 104860 339300 104866 339312
rect 132678 339300 132684 339312
rect 104860 339272 132684 339300
rect 104860 339260 104866 339272
rect 132678 339260 132684 339272
rect 132736 339260 132742 339312
rect 135254 339232 135260 339244
rect 122806 339204 135260 339232
rect 97718 339124 97724 339176
rect 97776 339164 97782 339176
rect 97902 339164 97908 339176
rect 97776 339136 97908 339164
rect 97776 339124 97782 339136
rect 97902 339124 97908 339136
rect 97960 339164 97966 339176
rect 117682 339164 117688 339176
rect 97960 339136 117688 339164
rect 97960 339124 97966 339136
rect 117682 339124 117688 339136
rect 117740 339124 117746 339176
rect 122806 339164 122834 339204
rect 135254 339192 135260 339204
rect 135312 339192 135318 339244
rect 117976 339136 122834 339164
rect 84838 339056 84844 339108
rect 84896 339096 84902 339108
rect 84896 339068 103514 339096
rect 84896 339056 84902 339068
rect 103486 338960 103514 339068
rect 110598 338988 110604 339040
rect 110656 339028 110662 339040
rect 111702 339028 111708 339040
rect 110656 339000 111708 339028
rect 110656 338988 110662 339000
rect 111702 338988 111708 339000
rect 111760 339028 111766 339040
rect 117976 339028 118004 339136
rect 199562 339096 199568 339108
rect 111760 339000 118004 339028
rect 122806 339068 199568 339096
rect 111760 338988 111766 339000
rect 122806 338960 122834 339068
rect 199562 339056 199568 339068
rect 199620 339056 199626 339108
rect 103486 338932 122834 338960
rect 68554 338852 68560 338904
rect 68612 338892 68618 338904
rect 98638 338892 98644 338904
rect 68612 338864 98644 338892
rect 68612 338852 68618 338864
rect 98638 338852 98644 338864
rect 98696 338852 98702 338904
rect 55122 338784 55128 338836
rect 55180 338824 55186 338836
rect 91002 338824 91008 338836
rect 55180 338796 91008 338824
rect 55180 338784 55186 338796
rect 91002 338784 91008 338796
rect 91060 338824 91066 338836
rect 91922 338824 91928 338836
rect 91060 338796 91928 338824
rect 91060 338784 91066 338796
rect 91922 338784 91928 338796
rect 91980 338784 91986 338836
rect 54846 338716 54852 338768
rect 54904 338756 54910 338768
rect 104802 338756 104808 338768
rect 54904 338728 104808 338756
rect 54904 338716 54910 338728
rect 104802 338716 104808 338728
rect 104860 338716 104866 338768
rect 79686 338172 79692 338224
rect 79744 338212 79750 338224
rect 83458 338212 83464 338224
rect 79744 338184 83464 338212
rect 79744 338172 79750 338184
rect 83458 338172 83464 338184
rect 83516 338172 83522 338224
rect 49510 338036 49516 338088
rect 49568 338076 49574 338088
rect 53374 338076 53380 338088
rect 49568 338048 53380 338076
rect 49568 338036 49574 338048
rect 53374 338036 53380 338048
rect 53432 338036 53438 338088
rect 103514 338036 103520 338088
rect 103572 338076 103578 338088
rect 131206 338076 131212 338088
rect 103572 338048 131212 338076
rect 103572 338036 103578 338048
rect 131206 338036 131212 338048
rect 131264 338036 131270 338088
rect 57698 337968 57704 338020
rect 57756 338008 57762 338020
rect 91278 338008 91284 338020
rect 57756 337980 91284 338008
rect 57756 337968 57762 337980
rect 91278 337968 91284 337980
rect 91336 338008 91342 338020
rect 91738 338008 91744 338020
rect 91336 337980 91744 338008
rect 91336 337968 91342 337980
rect 91738 337968 91744 337980
rect 91796 337968 91802 338020
rect 115750 337968 115756 338020
rect 115808 338008 115814 338020
rect 142246 338008 142252 338020
rect 115808 337980 142252 338008
rect 115808 337968 115814 337980
rect 142246 337968 142252 337980
rect 142304 338008 142310 338020
rect 143442 338008 143448 338020
rect 142304 337980 143448 338008
rect 142304 337968 142310 337980
rect 143442 337968 143448 337980
rect 143500 337968 143506 338020
rect 43714 337900 43720 337952
rect 43772 337940 43778 337952
rect 74534 337940 74540 337952
rect 43772 337912 74540 337940
rect 43772 337900 43778 337912
rect 74534 337900 74540 337912
rect 74592 337940 74598 337952
rect 75270 337940 75276 337952
rect 74592 337912 75276 337940
rect 74592 337900 74598 337912
rect 75270 337900 75276 337912
rect 75328 337900 75334 337952
rect 115198 337900 115204 337952
rect 115256 337940 115262 337952
rect 140038 337940 140044 337952
rect 115256 337912 140044 337940
rect 115256 337900 115262 337912
rect 140038 337900 140044 337912
rect 140096 337900 140102 337952
rect 50890 337832 50896 337884
rect 50948 337872 50954 337884
rect 86126 337872 86132 337884
rect 50948 337844 86132 337872
rect 50948 337832 50954 337844
rect 86126 337832 86132 337844
rect 86184 337872 86190 337884
rect 86862 337872 86868 337884
rect 86184 337844 86868 337872
rect 86184 337832 86190 337844
rect 86862 337832 86868 337844
rect 86920 337832 86926 337884
rect 119522 337872 119528 337884
rect 103486 337844 119528 337872
rect 99650 337696 99656 337748
rect 99708 337736 99714 337748
rect 100662 337736 100668 337748
rect 99708 337708 100668 337736
rect 99708 337696 99714 337708
rect 100662 337696 100668 337708
rect 100720 337736 100726 337748
rect 103486 337736 103514 337844
rect 119522 337832 119528 337844
rect 119580 337832 119586 337884
rect 109954 337764 109960 337816
rect 110012 337804 110018 337816
rect 126330 337804 126336 337816
rect 110012 337776 126336 337804
rect 110012 337764 110018 337776
rect 126330 337764 126336 337776
rect 126388 337764 126394 337816
rect 100720 337708 103514 337736
rect 100720 337696 100726 337708
rect 115198 337696 115204 337748
rect 115256 337736 115262 337748
rect 115382 337736 115388 337748
rect 115256 337708 115388 337736
rect 115256 337696 115262 337708
rect 115382 337696 115388 337708
rect 115440 337696 115446 337748
rect 45462 337492 45468 337544
rect 45520 337532 45526 337544
rect 70026 337532 70032 337544
rect 45520 337504 70032 337532
rect 45520 337492 45526 337504
rect 70026 337492 70032 337504
rect 70084 337492 70090 337544
rect 101398 337492 101404 337544
rect 101456 337532 101462 337544
rect 101456 337504 103514 337532
rect 101456 337492 101462 337504
rect 53374 337424 53380 337476
rect 53432 337464 53438 337476
rect 82262 337464 82268 337476
rect 53432 337436 82268 337464
rect 53432 337424 53438 337436
rect 82262 337424 82268 337436
rect 82320 337424 82326 337476
rect 101950 337424 101956 337476
rect 102008 337464 102014 337476
rect 102870 337464 102876 337476
rect 102008 337436 102876 337464
rect 102008 337424 102014 337436
rect 102870 337424 102876 337436
rect 102928 337424 102934 337476
rect 103486 337464 103514 337504
rect 115106 337464 115112 337476
rect 103486 337436 115112 337464
rect 115106 337424 115112 337436
rect 115164 337424 115170 337476
rect 150526 337424 150532 337476
rect 150584 337464 150590 337476
rect 151722 337464 151728 337476
rect 150584 337436 151728 337464
rect 150584 337424 150590 337436
rect 151722 337424 151728 337436
rect 151780 337464 151786 337476
rect 197354 337464 197360 337476
rect 151780 337436 197360 337464
rect 151780 337424 151786 337436
rect 197354 337424 197360 337436
rect 197412 337424 197418 337476
rect 53742 337356 53748 337408
rect 53800 337396 53806 337408
rect 55122 337396 55128 337408
rect 53800 337368 55128 337396
rect 53800 337356 53806 337368
rect 55122 337356 55128 337368
rect 55180 337396 55186 337408
rect 84194 337396 84200 337408
rect 55180 337368 84200 337396
rect 55180 337356 55186 337368
rect 84194 337356 84200 337368
rect 84252 337356 84258 337408
rect 86862 337356 86868 337408
rect 86920 337396 86926 337408
rect 86920 337368 103514 337396
rect 86920 337356 86926 337368
rect 103486 337328 103514 337368
rect 131206 337356 131212 337408
rect 131264 337396 131270 337408
rect 133874 337396 133880 337408
rect 131264 337368 133880 337396
rect 131264 337356 131270 337368
rect 133874 337356 133880 337368
rect 133932 337396 133938 337408
rect 196894 337396 196900 337408
rect 133932 337368 196900 337396
rect 133932 337356 133938 337368
rect 196894 337356 196900 337368
rect 196952 337356 196958 337408
rect 107562 337328 107568 337340
rect 103486 337300 107568 337328
rect 107562 337288 107568 337300
rect 107620 337328 107626 337340
rect 122190 337328 122196 337340
rect 107620 337300 122196 337328
rect 107620 337288 107626 337300
rect 122190 337288 122196 337300
rect 122248 337288 122254 337340
rect 91094 336812 91100 336864
rect 91152 336852 91158 336864
rect 94498 336852 94504 336864
rect 91152 336824 94504 336852
rect 91152 336812 91158 336824
rect 94498 336812 94504 336824
rect 94556 336812 94562 336864
rect 126330 336812 126336 336864
rect 126388 336852 126394 336864
rect 129734 336852 129740 336864
rect 126388 336824 129740 336852
rect 126388 336812 126394 336824
rect 129734 336812 129740 336824
rect 129792 336812 129798 336864
rect 75822 336744 75828 336796
rect 75880 336784 75886 336796
rect 97258 336784 97264 336796
rect 75880 336756 97264 336784
rect 75880 336744 75886 336756
rect 97258 336744 97264 336756
rect 97316 336744 97322 336796
rect 128998 336784 129004 336796
rect 128326 336756 129004 336784
rect 49602 336676 49608 336728
rect 49660 336716 49666 336728
rect 57238 336716 57244 336728
rect 49660 336688 57244 336716
rect 49660 336676 49666 336688
rect 57238 336676 57244 336688
rect 57296 336716 57302 336728
rect 91094 336716 91100 336728
rect 57296 336688 91100 336716
rect 57296 336676 57302 336688
rect 91094 336676 91100 336688
rect 91152 336676 91158 336728
rect 100294 336676 100300 336728
rect 100352 336716 100358 336728
rect 128326 336716 128354 336756
rect 128998 336744 129004 336756
rect 129056 336784 129062 336796
rect 138106 336784 138112 336796
rect 129056 336756 138112 336784
rect 129056 336744 129062 336756
rect 138106 336744 138112 336756
rect 138164 336744 138170 336796
rect 143442 336744 143448 336796
rect 143500 336784 143506 336796
rect 175918 336784 175924 336796
rect 143500 336756 175924 336784
rect 143500 336744 143506 336756
rect 175918 336744 175924 336756
rect 175976 336744 175982 336796
rect 100352 336688 128354 336716
rect 100352 336676 100358 336688
rect 54938 336608 54944 336660
rect 54996 336648 55002 336660
rect 89070 336648 89076 336660
rect 54996 336620 89076 336648
rect 54996 336608 55002 336620
rect 89070 336608 89076 336620
rect 89128 336608 89134 336660
rect 106182 336608 106188 336660
rect 106240 336648 106246 336660
rect 133966 336648 133972 336660
rect 106240 336620 133972 336648
rect 106240 336608 106246 336620
rect 133966 336608 133972 336620
rect 134024 336608 134030 336660
rect 56410 336540 56416 336592
rect 56468 336580 56474 336592
rect 86402 336580 86408 336592
rect 56468 336552 86408 336580
rect 56468 336540 56474 336552
rect 86402 336540 86408 336552
rect 86460 336540 86466 336592
rect 113818 336540 113824 336592
rect 113876 336580 113882 336592
rect 131114 336580 131120 336592
rect 113876 336552 131120 336580
rect 113876 336540 113882 336552
rect 131114 336540 131120 336552
rect 131172 336540 131178 336592
rect 48130 336472 48136 336524
rect 48188 336512 48194 336524
rect 76558 336512 76564 336524
rect 48188 336484 76564 336512
rect 48188 336472 48194 336484
rect 76558 336472 76564 336484
rect 76616 336472 76622 336524
rect 46750 336404 46756 336456
rect 46808 336444 46814 336456
rect 71958 336444 71964 336456
rect 46808 336416 71964 336444
rect 46808 336404 46814 336416
rect 71958 336404 71964 336416
rect 72016 336444 72022 336456
rect 72418 336444 72424 336456
rect 72016 336416 72424 336444
rect 72016 336404 72022 336416
rect 72418 336404 72424 336416
rect 72476 336404 72482 336456
rect 86218 336064 86224 336116
rect 86276 336104 86282 336116
rect 117958 336104 117964 336116
rect 86276 336076 117964 336104
rect 86276 336064 86282 336076
rect 117958 336064 117964 336076
rect 118016 336064 118022 336116
rect 66990 335996 66996 336048
rect 67048 336036 67054 336048
rect 121454 336036 121460 336048
rect 67048 336008 121460 336036
rect 67048 335996 67054 336008
rect 121454 335996 121460 336008
rect 121512 335996 121518 336048
rect 322474 335996 322480 336048
rect 322532 336036 322538 336048
rect 333974 336036 333980 336048
rect 322532 336008 333980 336036
rect 322532 335996 322538 336008
rect 333974 335996 333980 336008
rect 334032 335996 334038 336048
rect 195422 335588 195428 335640
rect 195480 335628 195486 335640
rect 197722 335628 197728 335640
rect 195480 335600 197728 335628
rect 195480 335588 195486 335600
rect 197722 335588 197728 335600
rect 197780 335588 197786 335640
rect 52086 335248 52092 335300
rect 52144 335288 52150 335300
rect 88702 335288 88708 335300
rect 52144 335260 88708 335288
rect 52144 335248 52150 335260
rect 88702 335248 88708 335260
rect 88760 335248 88766 335300
rect 92566 335248 92572 335300
rect 92624 335288 92630 335300
rect 93762 335288 93768 335300
rect 92624 335260 93768 335288
rect 92624 335248 92630 335260
rect 93762 335248 93768 335260
rect 93820 335288 93826 335300
rect 125686 335288 125692 335300
rect 93820 335260 125692 335288
rect 93820 335248 93826 335260
rect 125686 335248 125692 335260
rect 125744 335248 125750 335300
rect 46658 335180 46664 335232
rect 46716 335220 46722 335232
rect 80698 335220 80704 335232
rect 46716 335192 80704 335220
rect 46716 335180 46722 335192
rect 80698 335180 80704 335192
rect 80756 335180 80762 335232
rect 98362 335180 98368 335232
rect 98420 335220 98426 335232
rect 127342 335220 127348 335232
rect 98420 335192 127348 335220
rect 98420 335180 98426 335192
rect 127342 335180 127348 335192
rect 127400 335180 127406 335232
rect 42702 335112 42708 335164
rect 42760 335152 42766 335164
rect 75914 335152 75920 335164
rect 42760 335124 75920 335152
rect 42760 335112 42766 335124
rect 75914 335112 75920 335124
rect 75972 335112 75978 335164
rect 108022 335112 108028 335164
rect 108080 335152 108086 335164
rect 135438 335152 135444 335164
rect 108080 335124 135444 335152
rect 108080 335112 108086 335124
rect 135438 335112 135444 335124
rect 135496 335112 135502 335164
rect 52362 335044 52368 335096
rect 52420 335084 52426 335096
rect 84838 335084 84844 335096
rect 52420 335056 84844 335084
rect 52420 335044 52426 335056
rect 84838 335044 84844 335056
rect 84896 335044 84902 335096
rect 97810 335044 97816 335096
rect 97868 335084 97874 335096
rect 120258 335084 120264 335096
rect 97868 335056 120264 335084
rect 97868 335044 97874 335056
rect 120258 335044 120264 335056
rect 120316 335044 120322 335096
rect 121454 334568 121460 334620
rect 121512 334608 121518 334620
rect 131206 334608 131212 334620
rect 121512 334580 131212 334608
rect 121512 334568 121518 334580
rect 131206 334568 131212 334580
rect 131264 334608 131270 334620
rect 188430 334608 188436 334620
rect 131264 334580 188436 334608
rect 131264 334568 131270 334580
rect 188430 334568 188436 334580
rect 188488 334568 188494 334620
rect 322474 334568 322480 334620
rect 322532 334608 322538 334620
rect 325786 334608 325792 334620
rect 322532 334580 325792 334608
rect 322532 334568 322538 334580
rect 325786 334568 325792 334580
rect 325844 334608 325850 334620
rect 329834 334608 329840 334620
rect 325844 334580 329840 334608
rect 325844 334568 325850 334580
rect 329834 334568 329840 334580
rect 329892 334568 329898 334620
rect 97074 334500 97080 334552
rect 97132 334540 97138 334552
rect 97810 334540 97816 334552
rect 97132 334512 97816 334540
rect 97132 334500 97138 334512
rect 97810 334500 97816 334512
rect 97868 334500 97874 334552
rect 75914 334364 75920 334416
rect 75972 334404 75978 334416
rect 77110 334404 77116 334416
rect 75972 334376 77116 334404
rect 75972 334364 75978 334376
rect 77110 334364 77116 334376
rect 77168 334364 77174 334416
rect 50706 333956 50712 334008
rect 50764 333996 50770 334008
rect 52362 333996 52368 334008
rect 50764 333968 52368 333996
rect 50764 333956 50770 333968
rect 52362 333956 52368 333968
rect 52420 333956 52426 334008
rect 88702 333956 88708 334008
rect 88760 333996 88766 334008
rect 89162 333996 89168 334008
rect 88760 333968 89168 333996
rect 88760 333956 88766 333968
rect 89162 333956 89168 333968
rect 89220 333956 89226 334008
rect 127342 333956 127348 334008
rect 127400 333996 127406 334008
rect 128354 333996 128360 334008
rect 127400 333968 128360 333996
rect 127400 333956 127406 333968
rect 128354 333956 128360 333968
rect 128412 333956 128418 334008
rect 45278 333888 45284 333940
rect 45336 333928 45342 333940
rect 81618 333928 81624 333940
rect 45336 333900 81624 333928
rect 45336 333888 45342 333900
rect 81618 333888 81624 333900
rect 81676 333888 81682 333940
rect 95142 333888 95148 333940
rect 95200 333928 95206 333940
rect 128538 333928 128544 333940
rect 95200 333900 128544 333928
rect 95200 333888 95206 333900
rect 128538 333888 128544 333900
rect 128596 333928 128602 333940
rect 189718 333928 189724 333940
rect 128596 333900 189724 333928
rect 128596 333888 128602 333900
rect 189718 333888 189724 333900
rect 189776 333888 189782 333940
rect 53466 333820 53472 333872
rect 53524 333860 53530 333872
rect 87598 333860 87604 333872
rect 53524 333832 87604 333860
rect 53524 333820 53530 333832
rect 87598 333820 87604 333832
rect 87656 333820 87662 333872
rect 100938 333820 100944 333872
rect 100996 333860 101002 333872
rect 102042 333860 102048 333872
rect 100996 333832 102048 333860
rect 100996 333820 101002 333832
rect 102042 333820 102048 333832
rect 102100 333860 102106 333872
rect 132586 333860 132592 333872
rect 102100 333832 132592 333860
rect 102100 333820 102106 333832
rect 132586 333820 132592 333832
rect 132644 333820 132650 333872
rect 49326 333752 49332 333804
rect 49384 333792 49390 333804
rect 83550 333792 83556 333804
rect 49384 333764 83556 333792
rect 49384 333752 49390 333764
rect 83550 333752 83556 333764
rect 83608 333752 83614 333804
rect 189074 333208 189080 333260
rect 189132 333248 189138 333260
rect 190362 333248 190368 333260
rect 189132 333220 190368 333248
rect 189132 333208 189138 333220
rect 190362 333208 190368 333220
rect 190420 333248 190426 333260
rect 199470 333248 199476 333260
rect 190420 333220 199476 333248
rect 190420 333208 190426 333220
rect 199470 333208 199476 333220
rect 199528 333208 199534 333260
rect 333974 333208 333980 333260
rect 334032 333248 334038 333260
rect 371878 333248 371884 333260
rect 334032 333220 371884 333248
rect 334032 333208 334038 333220
rect 371878 333208 371884 333220
rect 371936 333208 371942 333260
rect 81618 332664 81624 332716
rect 81676 332704 81682 332716
rect 82078 332704 82084 332716
rect 81676 332676 82084 332704
rect 81676 332664 81682 332676
rect 82078 332664 82084 332676
rect 82136 332664 82142 332716
rect 48130 332596 48136 332648
rect 48188 332636 48194 332648
rect 53466 332636 53472 332648
rect 48188 332608 53472 332636
rect 48188 332596 48194 332608
rect 53466 332596 53472 332608
rect 53524 332596 53530 332648
rect 74626 332596 74632 332648
rect 74684 332636 74690 332648
rect 189074 332636 189080 332648
rect 74684 332608 189080 332636
rect 74684 332596 74690 332608
rect 189074 332596 189080 332608
rect 189132 332596 189138 332648
rect 47946 332528 47952 332580
rect 48004 332568 48010 332580
rect 78398 332568 78404 332580
rect 48004 332540 78404 332568
rect 48004 332528 48010 332540
rect 78398 332528 78404 332540
rect 78456 332528 78462 332580
rect 107378 332528 107384 332580
rect 107436 332568 107442 332580
rect 125502 332568 125508 332580
rect 107436 332540 125508 332568
rect 107436 332528 107442 332540
rect 125502 332528 125508 332540
rect 125560 332528 125566 332580
rect 104894 331984 104900 332036
rect 104952 332024 104958 332036
rect 127618 332024 127624 332036
rect 104952 331996 127624 332024
rect 104952 331984 104958 331996
rect 127618 331984 127624 331996
rect 127676 331984 127682 332036
rect 56410 331916 56416 331968
rect 56468 331956 56474 331968
rect 124306 331956 124312 331968
rect 56468 331928 124312 331956
rect 56468 331916 56474 331928
rect 124306 331916 124312 331928
rect 124364 331956 124370 331968
rect 159542 331956 159548 331968
rect 124364 331928 159548 331956
rect 124364 331916 124370 331928
rect 159542 331916 159548 331928
rect 159600 331916 159606 331968
rect 37090 331848 37096 331900
rect 37148 331888 37154 331900
rect 108022 331888 108028 331900
rect 37148 331860 108028 331888
rect 37148 331848 37154 331860
rect 108022 331848 108028 331860
rect 108080 331848 108086 331900
rect 122190 331848 122196 331900
rect 122248 331888 122254 331900
rect 124398 331888 124404 331900
rect 122248 331860 124404 331888
rect 122248 331848 122254 331860
rect 124398 331848 124404 331860
rect 124456 331888 124462 331900
rect 175182 331888 175188 331900
rect 124456 331860 175188 331888
rect 124456 331848 124462 331860
rect 175182 331848 175188 331860
rect 175240 331848 175246 331900
rect 322198 331712 322204 331764
rect 322256 331752 322262 331764
rect 327442 331752 327448 331764
rect 322256 331724 327448 331752
rect 322256 331712 322262 331724
rect 327442 331712 327448 331724
rect 327500 331712 327506 331764
rect 4798 331236 4804 331288
rect 4856 331276 4862 331288
rect 37090 331276 37096 331288
rect 4856 331248 37096 331276
rect 4856 331236 4862 331248
rect 37090 331236 37096 331248
rect 37148 331236 37154 331288
rect 77938 331236 77944 331288
rect 77996 331276 78002 331288
rect 78398 331276 78404 331288
rect 77996 331248 78404 331276
rect 77996 331236 78002 331248
rect 78398 331236 78404 331248
rect 78456 331236 78462 331288
rect 175182 331236 175188 331288
rect 175240 331276 175246 331288
rect 197354 331276 197360 331288
rect 175240 331248 197360 331276
rect 175240 331236 175246 331248
rect 197354 331236 197360 331248
rect 197412 331236 197418 331288
rect 93210 331168 93216 331220
rect 93268 331208 93274 331220
rect 122098 331208 122104 331220
rect 93268 331180 122104 331208
rect 93268 331168 93274 331180
rect 122098 331168 122104 331180
rect 122156 331208 122162 331220
rect 124306 331208 124312 331220
rect 122156 331180 124312 331208
rect 122156 331168 122162 331180
rect 124306 331168 124312 331180
rect 124364 331168 124370 331220
rect 322750 331032 322756 331084
rect 322808 331072 322814 331084
rect 324314 331072 324320 331084
rect 322808 331044 324320 331072
rect 322808 331032 322814 331044
rect 324314 331032 324320 331044
rect 324372 331032 324378 331084
rect 52086 330556 52092 330608
rect 52144 330596 52150 330608
rect 95050 330596 95056 330608
rect 52144 330568 95056 330596
rect 52144 330556 52150 330568
rect 95050 330556 95056 330568
rect 95108 330556 95114 330608
rect 95142 330556 95148 330608
rect 95200 330596 95206 330608
rect 113818 330596 113824 330608
rect 95200 330568 113824 330596
rect 95200 330556 95206 330568
rect 113818 330556 113824 330568
rect 113876 330556 113882 330608
rect 57790 330488 57796 330540
rect 57848 330528 57854 330540
rect 131114 330528 131120 330540
rect 57848 330500 131120 330528
rect 57848 330488 57854 330500
rect 131114 330488 131120 330500
rect 131172 330528 131178 330540
rect 160738 330528 160744 330540
rect 131172 330500 160744 330528
rect 131172 330488 131178 330500
rect 160738 330488 160744 330500
rect 160796 330488 160802 330540
rect 84286 329196 84292 329248
rect 84344 329236 84350 329248
rect 116026 329236 116032 329248
rect 84344 329208 116032 329236
rect 84344 329196 84350 329208
rect 116026 329196 116032 329208
rect 116084 329196 116090 329248
rect 103514 329128 103520 329180
rect 103572 329168 103578 329180
rect 151078 329168 151084 329180
rect 103572 329140 151084 329168
rect 103572 329128 103578 329140
rect 151078 329128 151084 329140
rect 151136 329128 151142 329180
rect 68738 329060 68744 329112
rect 68796 329100 68802 329112
rect 177390 329100 177396 329112
rect 68796 329072 177396 329100
rect 68796 329060 68802 329072
rect 177390 329060 177396 329072
rect 177448 329060 177454 329112
rect 123754 328448 123760 328500
rect 123812 328488 123818 328500
rect 124122 328488 124128 328500
rect 123812 328460 124128 328488
rect 123812 328448 123818 328460
rect 124122 328448 124128 328460
rect 124180 328488 124186 328500
rect 165522 328488 165528 328500
rect 124180 328460 165528 328488
rect 124180 328448 124186 328460
rect 165522 328448 165528 328460
rect 165580 328488 165586 328500
rect 197354 328488 197360 328500
rect 165580 328460 197360 328488
rect 165580 328448 165586 328460
rect 197354 328448 197360 328460
rect 197412 328448 197418 328500
rect 86310 327904 86316 327956
rect 86368 327944 86374 327956
rect 124122 327944 124128 327956
rect 86368 327916 124128 327944
rect 86368 327904 86374 327916
rect 124122 327904 124128 327916
rect 124180 327904 124186 327956
rect 111794 327836 111800 327888
rect 111852 327876 111858 327888
rect 174538 327876 174544 327888
rect 111852 327848 174544 327876
rect 111852 327836 111858 327848
rect 174538 327836 174544 327848
rect 174596 327836 174602 327888
rect 70486 327768 70492 327820
rect 70544 327808 70550 327820
rect 141418 327808 141424 327820
rect 70544 327780 141424 327808
rect 70544 327768 70550 327780
rect 141418 327768 141424 327780
rect 141476 327768 141482 327820
rect 88334 327700 88340 327752
rect 88392 327740 88398 327752
rect 178862 327740 178868 327752
rect 88392 327712 178868 327740
rect 88392 327700 88398 327712
rect 178862 327700 178868 327712
rect 178920 327700 178926 327752
rect 322750 327700 322756 327752
rect 322808 327740 322814 327752
rect 324314 327740 324320 327752
rect 322808 327712 324320 327740
rect 322808 327700 322814 327712
rect 324314 327700 324320 327712
rect 324372 327740 324378 327752
rect 482278 327740 482284 327752
rect 324372 327712 482284 327740
rect 324372 327700 324378 327712
rect 482278 327700 482284 327712
rect 482336 327700 482342 327752
rect 107470 327088 107476 327140
rect 107528 327128 107534 327140
rect 115290 327128 115296 327140
rect 107528 327100 115296 327128
rect 107528 327088 107534 327100
rect 115290 327088 115296 327100
rect 115348 327088 115354 327140
rect 185670 327088 185676 327140
rect 185728 327128 185734 327140
rect 197354 327128 197360 327140
rect 185728 327100 197360 327128
rect 185728 327088 185734 327100
rect 197354 327088 197360 327100
rect 197412 327088 197418 327140
rect 108666 327020 108672 327072
rect 108724 327060 108730 327072
rect 140866 327060 140872 327072
rect 108724 327032 140872 327060
rect 108724 327020 108730 327032
rect 140866 327020 140872 327032
rect 140924 327020 140930 327072
rect 93118 326544 93124 326596
rect 93176 326584 93182 326596
rect 115382 326584 115388 326596
rect 93176 326556 115388 326584
rect 93176 326544 93182 326556
rect 115382 326544 115388 326556
rect 115440 326544 115446 326596
rect 54938 326476 54944 326528
rect 54996 326516 55002 326528
rect 106918 326516 106924 326528
rect 54996 326488 106924 326516
rect 54996 326476 55002 326488
rect 106918 326476 106924 326488
rect 106976 326476 106982 326528
rect 115290 326476 115296 326528
rect 115348 326516 115354 326528
rect 162210 326516 162216 326528
rect 115348 326488 162216 326516
rect 115348 326476 115354 326488
rect 162210 326476 162216 326488
rect 162268 326476 162274 326528
rect 57698 326408 57704 326460
rect 57756 326448 57762 326460
rect 120166 326448 120172 326460
rect 57756 326420 120172 326448
rect 57756 326408 57762 326420
rect 120166 326408 120172 326420
rect 120224 326408 120230 326460
rect 140866 326408 140872 326460
rect 140924 326448 140930 326460
rect 152642 326448 152648 326460
rect 140924 326420 152648 326448
rect 140924 326408 140930 326420
rect 152642 326408 152648 326420
rect 152700 326408 152706 326460
rect 88978 326340 88984 326392
rect 89036 326380 89042 326392
rect 176010 326380 176016 326392
rect 89036 326352 176016 326380
rect 89036 326340 89042 326352
rect 176010 326340 176016 326352
rect 176068 326340 176074 326392
rect 322842 326340 322848 326392
rect 322900 326380 322906 326392
rect 494146 326380 494152 326392
rect 322900 326352 494152 326380
rect 322900 326340 322906 326352
rect 494146 326340 494152 326352
rect 494204 326340 494210 326392
rect 106182 325048 106188 325100
rect 106240 325088 106246 325100
rect 113818 325088 113824 325100
rect 106240 325060 113824 325088
rect 106240 325048 106246 325060
rect 113818 325048 113824 325060
rect 113876 325048 113882 325100
rect 71774 324980 71780 325032
rect 71832 325020 71838 325032
rect 166350 325020 166356 325032
rect 71832 324992 166356 325020
rect 71832 324980 71838 324992
rect 166350 324980 166356 324992
rect 166408 324980 166414 325032
rect 96614 324912 96620 324964
rect 96672 324952 96678 324964
rect 196802 324952 196808 324964
rect 96672 324924 196808 324952
rect 96672 324912 96678 324924
rect 196802 324912 196808 324924
rect 196860 324912 196866 324964
rect 360838 324912 360844 324964
rect 360896 324952 360902 324964
rect 380894 324952 380900 324964
rect 360896 324924 380900 324952
rect 360896 324912 360902 324924
rect 380894 324912 380900 324924
rect 380952 324912 380958 324964
rect 320358 324300 320364 324352
rect 320416 324340 320422 324352
rect 322842 324340 322848 324352
rect 320416 324312 322848 324340
rect 320416 324300 320422 324312
rect 322842 324300 322848 324312
rect 322900 324300 322906 324352
rect 380894 324300 380900 324352
rect 380952 324340 380958 324352
rect 382182 324340 382188 324352
rect 380952 324312 382188 324340
rect 380952 324300 380958 324312
rect 382182 324300 382188 324312
rect 382240 324340 382246 324352
rect 580166 324340 580172 324352
rect 382240 324312 580172 324340
rect 382240 324300 382246 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 49418 323688 49424 323740
rect 49476 323728 49482 323740
rect 117958 323728 117964 323740
rect 49476 323700 117964 323728
rect 49476 323688 49482 323700
rect 117958 323688 117964 323700
rect 118016 323688 118022 323740
rect 89162 323620 89168 323672
rect 89220 323660 89226 323672
rect 160738 323660 160744 323672
rect 89220 323632 160744 323660
rect 89220 323620 89226 323632
rect 160738 323620 160744 323632
rect 160796 323620 160802 323672
rect 73154 323552 73160 323604
rect 73212 323592 73218 323604
rect 164878 323592 164884 323604
rect 73212 323564 164884 323592
rect 73212 323552 73218 323564
rect 164878 323552 164884 323564
rect 164936 323552 164942 323604
rect 322474 322940 322480 322992
rect 322532 322980 322538 322992
rect 331214 322980 331220 322992
rect 322532 322952 331220 322980
rect 322532 322940 322538 322952
rect 331214 322940 331220 322952
rect 331272 322940 331278 322992
rect 128262 322872 128268 322924
rect 128320 322912 128326 322924
rect 134150 322912 134156 322924
rect 128320 322884 134156 322912
rect 128320 322872 128326 322884
rect 134150 322872 134156 322884
rect 134208 322912 134214 322924
rect 197354 322912 197360 322924
rect 134208 322884 197360 322912
rect 134208 322872 134214 322884
rect 197354 322872 197360 322884
rect 197412 322872 197418 322924
rect 70394 322192 70400 322244
rect 70452 322232 70458 322244
rect 170490 322232 170496 322244
rect 70452 322204 170496 322232
rect 70452 322192 70458 322204
rect 170490 322192 170496 322204
rect 170548 322192 170554 322244
rect 77938 320900 77944 320952
rect 77996 320940 78002 320952
rect 134518 320940 134524 320952
rect 77996 320912 134524 320940
rect 77996 320900 78002 320912
rect 134518 320900 134524 320912
rect 134576 320900 134582 320952
rect 49510 320832 49516 320884
rect 49568 320872 49574 320884
rect 148410 320872 148416 320884
rect 49568 320844 148416 320872
rect 49568 320832 49574 320844
rect 148410 320832 148416 320844
rect 148468 320832 148474 320884
rect 167822 320832 167828 320884
rect 167880 320872 167886 320884
rect 198182 320872 198188 320884
rect 167880 320844 198188 320872
rect 167880 320832 167886 320844
rect 198182 320832 198188 320844
rect 198240 320832 198246 320884
rect 172330 320152 172336 320204
rect 172388 320192 172394 320204
rect 197354 320192 197360 320204
rect 172388 320164 197360 320192
rect 172388 320152 172394 320164
rect 197354 320152 197360 320164
rect 197412 320152 197418 320204
rect 322842 320152 322848 320204
rect 322900 320192 322906 320204
rect 324314 320192 324320 320204
rect 322900 320164 324320 320192
rect 322900 320152 322906 320164
rect 324314 320152 324320 320164
rect 324372 320192 324378 320204
rect 499666 320192 499672 320204
rect 324372 320164 499672 320192
rect 324372 320152 324378 320164
rect 499666 320152 499672 320164
rect 499724 320152 499730 320204
rect 67450 319608 67456 319660
rect 67508 319648 67514 319660
rect 122098 319648 122104 319660
rect 67508 319620 122104 319648
rect 67508 319608 67514 319620
rect 122098 319608 122104 319620
rect 122156 319608 122162 319660
rect 117314 319540 117320 319592
rect 117372 319580 117378 319592
rect 180242 319580 180248 319592
rect 117372 319552 180248 319580
rect 117372 319540 117378 319552
rect 180242 319540 180248 319552
rect 180300 319540 180306 319592
rect 75178 319472 75184 319524
rect 75236 319512 75242 319524
rect 108666 319512 108672 319524
rect 75236 319484 108672 319512
rect 75236 319472 75242 319484
rect 108666 319472 108672 319484
rect 108724 319472 108730 319524
rect 111058 319472 111064 319524
rect 111116 319512 111122 319524
rect 177482 319512 177488 319524
rect 111116 319484 177488 319512
rect 111116 319472 111122 319484
rect 177482 319472 177488 319484
rect 177540 319472 177546 319524
rect 95326 319404 95332 319456
rect 95384 319444 95390 319456
rect 171778 319444 171784 319456
rect 95384 319416 171784 319444
rect 95384 319404 95390 319416
rect 171778 319404 171784 319416
rect 171836 319404 171842 319456
rect 3418 319064 3424 319116
rect 3476 319104 3482 319116
rect 7558 319104 7564 319116
rect 3476 319076 7564 319104
rect 3476 319064 3482 319076
rect 7558 319064 7564 319076
rect 7616 319064 7622 319116
rect 112530 318724 112536 318776
rect 112588 318764 112594 318776
rect 143534 318764 143540 318776
rect 112588 318736 143540 318764
rect 112588 318724 112594 318736
rect 143534 318724 143540 318736
rect 143592 318764 143598 318776
rect 144822 318764 144828 318776
rect 143592 318736 144828 318764
rect 143592 318724 143598 318736
rect 144822 318724 144828 318736
rect 144880 318724 144886 318776
rect 84378 318112 84384 318164
rect 84436 318152 84442 318164
rect 113910 318152 113916 318164
rect 84436 318124 113916 318152
rect 84436 318112 84442 318124
rect 113910 318112 113916 318124
rect 113968 318112 113974 318164
rect 65610 318044 65616 318096
rect 65668 318084 65674 318096
rect 115198 318084 115204 318096
rect 65668 318056 115204 318084
rect 65668 318044 65674 318056
rect 115198 318044 115204 318056
rect 115256 318044 115262 318096
rect 144822 318044 144828 318096
rect 144880 318084 144886 318096
rect 171778 318084 171784 318096
rect 144880 318056 171784 318084
rect 144880 318044 144886 318056
rect 171778 318044 171784 318056
rect 171836 318044 171842 318096
rect 115842 317500 115848 317552
rect 115900 317540 115906 317552
rect 128630 317540 128636 317552
rect 115900 317512 128636 317540
rect 115900 317500 115906 317512
rect 128630 317500 128636 317512
rect 128688 317540 128694 317552
rect 155310 317540 155316 317552
rect 128688 317512 155316 317540
rect 128688 317500 128694 317512
rect 155310 317500 155316 317512
rect 155368 317500 155374 317552
rect 116670 317432 116676 317484
rect 116728 317472 116734 317484
rect 193122 317472 193128 317484
rect 116728 317444 193128 317472
rect 116728 317432 116734 317444
rect 193122 317432 193128 317444
rect 193180 317472 193186 317484
rect 197354 317472 197360 317484
rect 193180 317444 197360 317472
rect 193180 317432 193186 317444
rect 197354 317432 197360 317444
rect 197412 317432 197418 317484
rect 101950 317364 101956 317416
rect 102008 317404 102014 317416
rect 131298 317404 131304 317416
rect 102008 317376 131304 317404
rect 102008 317364 102014 317376
rect 131298 317364 131304 317376
rect 131356 317404 131362 317416
rect 131482 317404 131488 317416
rect 131356 317376 131488 317404
rect 131356 317364 131362 317376
rect 131482 317364 131488 317376
rect 131540 317364 131546 317416
rect 322474 317364 322480 317416
rect 322532 317404 322538 317416
rect 335446 317404 335452 317416
rect 322532 317376 335452 317404
rect 322532 317364 322538 317376
rect 335446 317364 335452 317376
rect 335504 317404 335510 317416
rect 336642 317404 336648 317416
rect 335504 317376 336648 317404
rect 335504 317364 335510 317376
rect 336642 317364 336648 317376
rect 336700 317364 336706 317416
rect 93946 316820 93952 316872
rect 94004 316860 94010 316872
rect 115842 316860 115848 316872
rect 94004 316832 115848 316860
rect 94004 316820 94010 316832
rect 115842 316820 115848 316832
rect 115900 316820 115906 316872
rect 131482 316820 131488 316872
rect 131540 316860 131546 316872
rect 151078 316860 151084 316872
rect 131540 316832 151084 316860
rect 131540 316820 131546 316832
rect 151078 316820 151084 316832
rect 151136 316820 151142 316872
rect 69474 316752 69480 316804
rect 69532 316792 69538 316804
rect 107102 316792 107108 316804
rect 69532 316764 107108 316792
rect 69532 316752 69538 316764
rect 107102 316752 107108 316764
rect 107160 316752 107166 316804
rect 111610 316752 111616 316804
rect 111668 316792 111674 316804
rect 177482 316792 177488 316804
rect 111668 316764 177488 316792
rect 111668 316752 111674 316764
rect 177482 316752 177488 316764
rect 177540 316752 177546 316804
rect 80698 316684 80704 316736
rect 80756 316724 80762 316736
rect 191098 316724 191104 316736
rect 80756 316696 191104 316724
rect 80756 316684 80762 316696
rect 191098 316684 191104 316696
rect 191156 316684 191162 316736
rect 336642 316684 336648 316736
rect 336700 316724 336706 316736
rect 454678 316724 454684 316736
rect 336700 316696 454684 316724
rect 336700 316684 336706 316696
rect 454678 316684 454684 316696
rect 454736 316684 454742 316736
rect 75270 315936 75276 315988
rect 75328 315976 75334 315988
rect 114646 315976 114652 315988
rect 75328 315948 114652 315976
rect 75328 315936 75334 315948
rect 114646 315936 114652 315948
rect 114704 315936 114710 315988
rect 114646 315324 114652 315376
rect 114704 315364 114710 315376
rect 115290 315364 115296 315376
rect 114704 315336 115296 315364
rect 114704 315324 114710 315336
rect 115290 315324 115296 315336
rect 115348 315324 115354 315376
rect 79410 315256 79416 315308
rect 79468 315296 79474 315308
rect 136818 315296 136824 315308
rect 79468 315268 136824 315296
rect 79468 315256 79474 315268
rect 136818 315256 136824 315268
rect 136876 315296 136882 315308
rect 166534 315296 166540 315308
rect 136876 315268 166540 315296
rect 136876 315256 136882 315268
rect 166534 315256 166540 315268
rect 166592 315256 166598 315308
rect 102778 314644 102784 314696
rect 102836 314684 102842 314696
rect 184842 314684 184848 314696
rect 102836 314656 184848 314684
rect 102836 314644 102842 314656
rect 184842 314644 184848 314656
rect 184900 314684 184906 314696
rect 197354 314684 197360 314696
rect 184900 314656 197360 314684
rect 184900 314644 184906 314656
rect 197354 314644 197360 314656
rect 197412 314644 197418 314696
rect 7558 314576 7564 314628
rect 7616 314616 7622 314628
rect 48038 314616 48044 314628
rect 7616 314588 48044 314616
rect 7616 314576 7622 314588
rect 48038 314576 48044 314588
rect 48096 314576 48102 314628
rect 105446 314576 105452 314628
rect 105504 314616 105510 314628
rect 136726 314616 136732 314628
rect 105504 314588 136732 314616
rect 105504 314576 105510 314588
rect 136726 314576 136732 314588
rect 136784 314576 136790 314628
rect 322474 314576 322480 314628
rect 322532 314616 322538 314628
rect 331306 314616 331312 314628
rect 322532 314588 331312 314616
rect 322532 314576 322538 314588
rect 331306 314576 331312 314588
rect 331364 314576 331370 314628
rect 82078 314032 82084 314084
rect 82136 314072 82142 314084
rect 144178 314072 144184 314084
rect 82136 314044 144184 314072
rect 82136 314032 82142 314044
rect 144178 314032 144184 314044
rect 144236 314032 144242 314084
rect 90910 313964 90916 314016
rect 90968 314004 90974 314016
rect 153930 314004 153936 314016
rect 90968 313976 153936 314004
rect 90968 313964 90974 313976
rect 153930 313964 153936 313976
rect 153988 313964 153994 314016
rect 48038 313896 48044 313948
rect 48096 313936 48102 313948
rect 116578 313936 116584 313948
rect 48096 313908 116584 313936
rect 48096 313896 48102 313908
rect 116578 313896 116584 313908
rect 116636 313896 116642 313948
rect 136726 313896 136732 313948
rect 136784 313936 136790 313948
rect 163498 313936 163504 313948
rect 136784 313908 163504 313936
rect 136784 313896 136790 313908
rect 163498 313896 163504 313908
rect 163556 313896 163562 313948
rect 331306 313896 331312 313948
rect 331364 313936 331370 313948
rect 500954 313936 500960 313948
rect 331364 313908 500960 313936
rect 331364 313896 331370 313908
rect 500954 313896 500960 313908
rect 501012 313896 501018 313948
rect 129090 313284 129096 313336
rect 129148 313324 129154 313336
rect 197354 313324 197360 313336
rect 129148 313296 197360 313324
rect 129148 313284 129154 313296
rect 197354 313284 197360 313296
rect 197412 313284 197418 313336
rect 60458 312672 60464 312724
rect 60516 312712 60522 312724
rect 122190 312712 122196 312724
rect 60516 312684 122196 312712
rect 60516 312672 60522 312684
rect 122190 312672 122196 312684
rect 122248 312672 122254 312724
rect 97258 312604 97264 312656
rect 97316 312644 97322 312656
rect 164878 312644 164884 312656
rect 97316 312616 164884 312644
rect 97316 312604 97322 312616
rect 164878 312604 164884 312616
rect 164936 312604 164942 312656
rect 81434 312536 81440 312588
rect 81492 312576 81498 312588
rect 163590 312576 163596 312588
rect 81492 312548 163596 312576
rect 81492 312536 81498 312548
rect 163590 312536 163596 312548
rect 163648 312536 163654 312588
rect 181530 312536 181536 312588
rect 181588 312576 181594 312588
rect 195422 312576 195428 312588
rect 181588 312548 195428 312576
rect 181588 312536 181594 312548
rect 195422 312536 195428 312548
rect 195480 312536 195486 312588
rect 322842 312536 322848 312588
rect 322900 312576 322906 312588
rect 324498 312576 324504 312588
rect 322900 312548 324504 312576
rect 322900 312536 322906 312548
rect 324498 312536 324504 312548
rect 324556 312576 324562 312588
rect 395338 312576 395344 312588
rect 324556 312548 395344 312576
rect 324556 312536 324562 312548
rect 395338 312536 395344 312548
rect 395396 312536 395402 312588
rect 97810 311176 97816 311228
rect 97868 311216 97874 311228
rect 156598 311216 156604 311228
rect 97868 311188 156604 311216
rect 97868 311176 97874 311188
rect 156598 311176 156604 311188
rect 156656 311176 156662 311228
rect 72418 311108 72424 311160
rect 72476 311148 72482 311160
rect 148410 311148 148416 311160
rect 72476 311120 148416 311148
rect 72476 311108 72482 311120
rect 148410 311108 148416 311120
rect 148468 311108 148474 311160
rect 186314 311108 186320 311160
rect 186372 311148 186378 311160
rect 187602 311148 187608 311160
rect 186372 311120 187608 311148
rect 186372 311108 186378 311120
rect 187602 311108 187608 311120
rect 187660 311148 187666 311160
rect 198090 311148 198096 311160
rect 187660 311120 198096 311148
rect 187660 311108 187666 311120
rect 198090 311108 198096 311120
rect 198148 311108 198154 311160
rect 89714 310564 89720 310616
rect 89772 310604 89778 310616
rect 188982 310604 188988 310616
rect 89772 310576 188988 310604
rect 89772 310564 89778 310576
rect 188982 310564 188988 310576
rect 189040 310604 189046 310616
rect 197354 310604 197360 310616
rect 189040 310576 197360 310604
rect 189040 310564 189046 310576
rect 197354 310564 197360 310576
rect 197412 310564 197418 310616
rect 66162 310496 66168 310548
rect 66220 310536 66226 310548
rect 186314 310536 186320 310548
rect 66220 310508 186320 310536
rect 66220 310496 66226 310508
rect 186314 310496 186320 310508
rect 186372 310496 186378 310548
rect 107102 310428 107108 310480
rect 107160 310468 107166 310480
rect 125778 310468 125784 310480
rect 107160 310440 125784 310468
rect 107160 310428 107166 310440
rect 125778 310428 125784 310440
rect 125836 310468 125842 310480
rect 172330 310468 172336 310480
rect 125836 310440 172336 310468
rect 125836 310428 125842 310440
rect 172330 310428 172336 310440
rect 172388 310468 172394 310480
rect 173342 310468 173348 310480
rect 172388 310440 173348 310468
rect 172388 310428 172394 310440
rect 173342 310428 173348 310440
rect 173400 310428 173406 310480
rect 89070 309748 89076 309800
rect 89128 309788 89134 309800
rect 152458 309788 152464 309800
rect 89128 309760 152464 309788
rect 89128 309748 89134 309760
rect 152458 309748 152464 309760
rect 152516 309748 152522 309800
rect 322474 309748 322480 309800
rect 322532 309788 322538 309800
rect 325694 309788 325700 309800
rect 322532 309760 325700 309788
rect 322532 309748 322538 309760
rect 325694 309748 325700 309760
rect 325752 309788 325758 309800
rect 377398 309788 377404 309800
rect 325752 309760 377404 309788
rect 325752 309748 325758 309760
rect 377398 309748 377404 309760
rect 377456 309748 377462 309800
rect 178862 309204 178868 309256
rect 178920 309244 178926 309256
rect 197354 309244 197360 309256
rect 178920 309216 197360 309244
rect 178920 309204 178926 309216
rect 197354 309204 197360 309216
rect 197412 309204 197418 309256
rect 73890 309136 73896 309188
rect 73948 309176 73954 309188
rect 185670 309176 185676 309188
rect 73948 309148 185676 309176
rect 73948 309136 73954 309148
rect 185670 309136 185676 309148
rect 185728 309136 185734 309188
rect 126882 309068 126888 309120
rect 126940 309108 126946 309120
rect 131298 309108 131304 309120
rect 126940 309080 131304 309108
rect 126940 309068 126946 309080
rect 131298 309068 131304 309080
rect 131356 309068 131362 309120
rect 96522 308524 96528 308576
rect 96580 308564 96586 308576
rect 138658 308564 138664 308576
rect 96580 308536 138664 308564
rect 96580 308524 96586 308536
rect 138658 308524 138664 308536
rect 138716 308524 138722 308576
rect 73798 308456 73804 308508
rect 73856 308496 73862 308508
rect 119890 308496 119896 308508
rect 73856 308468 119896 308496
rect 73856 308456 73862 308468
rect 119890 308456 119896 308468
rect 119948 308456 119954 308508
rect 83550 308388 83556 308440
rect 83608 308428 83614 308440
rect 146938 308428 146944 308440
rect 83608 308400 146944 308428
rect 83608 308388 83614 308400
rect 146938 308388 146944 308400
rect 146996 308388 147002 308440
rect 165430 308388 165436 308440
rect 165488 308428 165494 308440
rect 198274 308428 198280 308440
rect 165488 308400 198280 308428
rect 165488 308388 165494 308400
rect 198274 308388 198280 308400
rect 198332 308388 198338 308440
rect 73062 307096 73068 307148
rect 73120 307136 73126 307148
rect 135990 307136 135996 307148
rect 73120 307108 135996 307136
rect 73120 307096 73126 307108
rect 135990 307096 135996 307108
rect 136048 307096 136054 307148
rect 85574 307028 85580 307080
rect 85632 307068 85638 307080
rect 196710 307068 196716 307080
rect 85632 307040 196716 307068
rect 85632 307028 85638 307040
rect 196710 307028 196716 307040
rect 196768 307028 196774 307080
rect 321738 307028 321744 307080
rect 321796 307068 321802 307080
rect 475378 307068 475384 307080
rect 321796 307040 475384 307068
rect 321796 307028 321802 307040
rect 475378 307028 475384 307040
rect 475436 307028 475442 307080
rect 70394 306484 70400 306536
rect 70452 306524 70458 306536
rect 70452 306496 196664 306524
rect 70452 306484 70458 306496
rect 87598 306416 87604 306468
rect 87656 306456 87662 306468
rect 162210 306456 162216 306468
rect 87656 306428 162216 306456
rect 87656 306416 87662 306428
rect 162210 306416 162216 306428
rect 162268 306416 162274 306468
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 15838 306320 15844 306332
rect 3476 306292 15844 306320
rect 3476 306280 3482 306292
rect 15838 306280 15844 306292
rect 15896 306280 15902 306332
rect 196636 306320 196664 306496
rect 197446 306320 197452 306332
rect 196636 306292 197452 306320
rect 197446 306280 197452 306292
rect 197504 306320 197510 306332
rect 199378 306320 199384 306332
rect 197504 306292 199384 306320
rect 197504 306280 197510 306292
rect 199378 306280 199384 306292
rect 199436 306280 199442 306332
rect 91002 305736 91008 305788
rect 91060 305776 91066 305788
rect 136726 305776 136732 305788
rect 91060 305748 136732 305776
rect 91060 305736 91066 305748
rect 136726 305736 136732 305748
rect 136784 305736 136790 305788
rect 79318 305668 79324 305720
rect 79376 305708 79382 305720
rect 142798 305708 142804 305720
rect 79376 305680 142804 305708
rect 79376 305668 79382 305680
rect 142798 305668 142804 305680
rect 142856 305668 142862 305720
rect 102042 305600 102048 305652
rect 102100 305640 102106 305652
rect 166350 305640 166356 305652
rect 102100 305612 166356 305640
rect 102100 305600 102106 305612
rect 166350 305600 166356 305612
rect 166408 305600 166414 305652
rect 111150 304988 111156 305040
rect 111208 305028 111214 305040
rect 167822 305028 167828 305040
rect 111208 305000 167828 305028
rect 111208 304988 111214 305000
rect 167822 304988 167828 305000
rect 167880 304988 167886 305040
rect 322474 304988 322480 305040
rect 322532 305028 322538 305040
rect 327166 305028 327172 305040
rect 322532 305000 327172 305028
rect 322532 304988 322538 305000
rect 327166 304988 327172 305000
rect 327224 304988 327230 305040
rect 91738 304308 91744 304360
rect 91796 304348 91802 304360
rect 149698 304348 149704 304360
rect 91796 304320 149704 304348
rect 91796 304308 91802 304320
rect 149698 304308 149704 304320
rect 149756 304308 149762 304360
rect 55030 304240 55036 304292
rect 55088 304280 55094 304292
rect 134610 304280 134616 304292
rect 55088 304252 134616 304280
rect 55088 304240 55094 304252
rect 134610 304240 134616 304252
rect 134668 304240 134674 304292
rect 119890 303968 119896 304020
rect 119948 304008 119954 304020
rect 123754 304008 123760 304020
rect 119948 303980 123760 304008
rect 119948 303968 119954 303980
rect 123754 303968 123760 303980
rect 123812 303968 123818 304020
rect 69198 303628 69204 303680
rect 69256 303668 69262 303680
rect 197722 303668 197728 303680
rect 69256 303640 197728 303668
rect 69256 303628 69262 303640
rect 197722 303628 197728 303640
rect 197780 303668 197786 303680
rect 198642 303668 198648 303680
rect 197780 303640 198648 303668
rect 197780 303628 197786 303640
rect 198642 303628 198648 303640
rect 198700 303628 198706 303680
rect 99282 303016 99288 303068
rect 99340 303056 99346 303068
rect 140038 303056 140044 303068
rect 99340 303028 140044 303056
rect 99340 303016 99346 303028
rect 140038 303016 140044 303028
rect 140096 303016 140102 303068
rect 66070 302948 66076 303000
rect 66128 302988 66134 303000
rect 130562 302988 130568 303000
rect 66128 302960 130568 302988
rect 66128 302948 66134 302960
rect 130562 302948 130568 302960
rect 130620 302948 130626 303000
rect 79318 302880 79324 302932
rect 79376 302920 79382 302932
rect 147030 302920 147036 302932
rect 79376 302892 147036 302920
rect 79376 302880 79382 302892
rect 147030 302880 147036 302892
rect 147088 302880 147094 302932
rect 186222 302880 186228 302932
rect 186280 302920 186286 302932
rect 197998 302920 198004 302932
rect 186280 302892 198004 302920
rect 186280 302880 186286 302892
rect 197998 302880 198004 302892
rect 198056 302880 198062 302932
rect 113266 302336 113272 302388
rect 113324 302376 113330 302388
rect 116670 302376 116676 302388
rect 113324 302348 116676 302376
rect 113324 302336 113330 302348
rect 116670 302336 116676 302348
rect 116728 302336 116734 302388
rect 48038 302268 48044 302320
rect 48096 302308 48102 302320
rect 69106 302308 69112 302320
rect 48096 302280 69112 302308
rect 48096 302268 48102 302280
rect 69106 302268 69112 302280
rect 69164 302308 69170 302320
rect 69474 302308 69480 302320
rect 69164 302280 69480 302308
rect 69164 302268 69170 302280
rect 69474 302268 69480 302280
rect 69532 302268 69538 302320
rect 86954 302268 86960 302320
rect 87012 302308 87018 302320
rect 163590 302308 163596 302320
rect 87012 302280 163596 302308
rect 87012 302268 87018 302280
rect 163590 302268 163596 302280
rect 163648 302268 163654 302320
rect 64506 302200 64512 302252
rect 64564 302240 64570 302252
rect 193030 302240 193036 302252
rect 64564 302212 193036 302240
rect 64564 302200 64570 302212
rect 193030 302200 193036 302212
rect 193088 302240 193094 302252
rect 197354 302240 197360 302252
rect 193088 302212 197360 302240
rect 193088 302200 193094 302212
rect 197354 302200 197360 302212
rect 197412 302200 197418 302252
rect 322474 302200 322480 302252
rect 322532 302240 322538 302252
rect 325694 302240 325700 302252
rect 322532 302212 325700 302240
rect 322532 302200 322538 302212
rect 325694 302200 325700 302212
rect 325752 302200 325758 302252
rect 58986 301656 58992 301708
rect 59044 301696 59050 301708
rect 101398 301696 101404 301708
rect 59044 301668 101404 301696
rect 59044 301656 59050 301668
rect 101398 301656 101404 301668
rect 101456 301656 101462 301708
rect 93762 301588 93768 301640
rect 93820 301628 93826 301640
rect 137278 301628 137284 301640
rect 93820 301600 137284 301628
rect 93820 301588 93826 301600
rect 137278 301588 137284 301600
rect 137336 301588 137342 301640
rect 87690 301520 87696 301572
rect 87748 301560 87754 301572
rect 143810 301560 143816 301572
rect 87748 301532 143816 301560
rect 87748 301520 87754 301532
rect 143810 301520 143816 301532
rect 143868 301560 143874 301572
rect 162302 301560 162308 301572
rect 143868 301532 162308 301560
rect 143868 301520 143874 301532
rect 162302 301520 162308 301532
rect 162360 301520 162366 301572
rect 69474 301452 69480 301504
rect 69532 301492 69538 301504
rect 184750 301492 184756 301504
rect 69532 301464 184756 301492
rect 69532 301452 69538 301464
rect 184750 301452 184756 301464
rect 184808 301452 184814 301504
rect 66898 301316 66904 301368
rect 66956 301356 66962 301368
rect 68830 301356 68836 301368
rect 66956 301328 68836 301356
rect 66956 301316 66962 301328
rect 68830 301316 68836 301328
rect 68888 301316 68894 301368
rect 102134 300908 102140 300960
rect 102192 300948 102198 300960
rect 133230 300948 133236 300960
rect 102192 300920 133236 300948
rect 102192 300908 102198 300920
rect 133230 300908 133236 300920
rect 133288 300908 133294 300960
rect 68830 300840 68836 300892
rect 68888 300880 68894 300892
rect 162394 300880 162400 300892
rect 68888 300852 162400 300880
rect 68888 300840 68894 300852
rect 162394 300840 162400 300852
rect 162452 300840 162458 300892
rect 98546 300636 98552 300688
rect 98604 300676 98610 300688
rect 102778 300676 102784 300688
rect 98604 300648 102784 300676
rect 98604 300636 98610 300648
rect 102778 300636 102784 300648
rect 102836 300636 102842 300688
rect 117866 300228 117872 300280
rect 117924 300268 117930 300280
rect 125594 300268 125600 300280
rect 117924 300240 125600 300268
rect 117924 300228 117930 300240
rect 125594 300228 125600 300240
rect 125652 300268 125658 300280
rect 148502 300268 148508 300280
rect 125652 300240 148508 300268
rect 125652 300228 125658 300240
rect 148502 300228 148508 300240
rect 148560 300228 148566 300280
rect 104986 300160 104992 300212
rect 105044 300200 105050 300212
rect 139394 300200 139400 300212
rect 105044 300172 139400 300200
rect 105044 300160 105050 300172
rect 139394 300160 139400 300172
rect 139452 300200 139458 300212
rect 170582 300200 170588 300212
rect 139452 300172 170588 300200
rect 139452 300160 139458 300172
rect 170582 300160 170588 300172
rect 170640 300160 170646 300212
rect 184750 300160 184756 300212
rect 184808 300200 184814 300212
rect 197354 300200 197360 300212
rect 184808 300172 197360 300200
rect 184808 300160 184814 300172
rect 197354 300160 197360 300172
rect 197412 300160 197418 300212
rect 146386 300132 146392 300144
rect 103486 300104 146392 300132
rect 100754 300024 100760 300076
rect 100812 300064 100818 300076
rect 101214 300064 101220 300076
rect 100812 300036 101220 300064
rect 100812 300024 100818 300036
rect 101214 300024 101220 300036
rect 101272 300064 101278 300076
rect 103486 300064 103514 300104
rect 146386 300092 146392 300104
rect 146444 300092 146450 300144
rect 176562 300092 176568 300144
rect 176620 300132 176626 300144
rect 197262 300132 197268 300144
rect 176620 300104 197268 300132
rect 176620 300092 176626 300104
rect 197262 300092 197268 300104
rect 197320 300092 197326 300144
rect 322566 300092 322572 300144
rect 322624 300132 322630 300144
rect 322750 300132 322756 300144
rect 322624 300104 322756 300132
rect 322624 300092 322630 300104
rect 322750 300092 322756 300104
rect 322808 300132 322814 300144
rect 356698 300132 356704 300144
rect 322808 300104 356704 300132
rect 322808 300092 322814 300104
rect 356698 300092 356704 300104
rect 356756 300092 356762 300144
rect 361482 300092 361488 300144
rect 361540 300132 361546 300144
rect 580258 300132 580264 300144
rect 361540 300104 580264 300132
rect 361540 300092 361546 300104
rect 580258 300092 580264 300104
rect 580316 300092 580322 300144
rect 101272 300036 103514 300064
rect 101272 300024 101278 300036
rect 82814 299684 82820 299736
rect 82872 299724 82878 299736
rect 136082 299724 136088 299736
rect 82872 299696 136088 299724
rect 82872 299684 82878 299696
rect 136082 299684 136088 299696
rect 136140 299684 136146 299736
rect 52362 299616 52368 299668
rect 52420 299656 52426 299668
rect 100754 299656 100760 299668
rect 52420 299628 100760 299656
rect 52420 299616 52426 299628
rect 100754 299616 100760 299628
rect 100812 299616 100818 299668
rect 109678 299616 109684 299668
rect 109736 299656 109742 299668
rect 115566 299656 115572 299668
rect 109736 299628 115572 299656
rect 109736 299616 109742 299628
rect 115566 299616 115572 299628
rect 115624 299656 115630 299668
rect 176562 299656 176568 299668
rect 115624 299628 176568 299656
rect 115624 299616 115630 299628
rect 176562 299616 176568 299628
rect 176620 299616 176626 299668
rect 81894 299548 81900 299600
rect 81952 299588 81958 299600
rect 169018 299588 169024 299600
rect 81952 299560 169024 299588
rect 81952 299548 81958 299560
rect 169018 299548 169024 299560
rect 169076 299548 169082 299600
rect 11698 299480 11704 299532
rect 11756 299520 11762 299532
rect 117866 299520 117872 299532
rect 11756 299492 117872 299520
rect 11756 299480 11762 299492
rect 117866 299480 117872 299492
rect 117924 299480 117930 299532
rect 94498 299072 94504 299124
rect 94556 299112 94562 299124
rect 95142 299112 95148 299124
rect 94556 299084 95148 299112
rect 94556 299072 94562 299084
rect 95142 299072 95148 299084
rect 95200 299072 95206 299124
rect 111702 298800 111708 298852
rect 111760 298840 111766 298852
rect 133138 298840 133144 298852
rect 111760 298812 133144 298840
rect 111760 298800 111766 298812
rect 133138 298800 133144 298812
rect 133196 298800 133202 298852
rect 83458 298732 83464 298784
rect 83516 298772 83522 298784
rect 129734 298772 129740 298784
rect 83516 298744 129740 298772
rect 83516 298732 83522 298744
rect 129734 298732 129740 298744
rect 129792 298732 129798 298784
rect 94498 298324 94504 298376
rect 94556 298364 94562 298376
rect 152734 298364 152740 298376
rect 94556 298336 152740 298364
rect 94556 298324 94562 298336
rect 152734 298324 152740 298336
rect 152792 298324 152798 298376
rect 99650 298256 99656 298308
rect 99708 298296 99714 298308
rect 189718 298296 189724 298308
rect 99708 298268 189724 298296
rect 99708 298256 99714 298268
rect 189718 298256 189724 298268
rect 189776 298256 189782 298308
rect 65518 298228 65524 298240
rect 64846 298200 65524 298228
rect 53650 298052 53656 298104
rect 53708 298092 53714 298104
rect 64846 298092 64874 298200
rect 65518 298188 65524 298200
rect 65576 298228 65582 298240
rect 167914 298228 167920 298240
rect 65576 298200 167920 298228
rect 65576 298188 65582 298200
rect 167914 298188 167920 298200
rect 167972 298188 167978 298240
rect 75270 298120 75276 298172
rect 75328 298160 75334 298172
rect 182910 298160 182916 298172
rect 75328 298132 182916 298160
rect 75328 298120 75334 298132
rect 182910 298120 182916 298132
rect 182968 298120 182974 298172
rect 53708 298064 64874 298092
rect 53708 298052 53714 298064
rect 50798 297508 50804 297560
rect 50856 297548 50862 297560
rect 56226 297548 56232 297560
rect 50856 297520 56232 297548
rect 50856 297508 50862 297520
rect 56226 297508 56232 297520
rect 56284 297548 56290 297560
rect 67542 297548 67548 297560
rect 56284 297520 67548 297548
rect 56284 297508 56290 297520
rect 67542 297508 67548 297520
rect 67600 297508 67606 297560
rect 25498 297372 25504 297424
rect 25556 297412 25562 297424
rect 56318 297412 56324 297424
rect 25556 297384 56324 297412
rect 25556 297372 25562 297384
rect 56318 297372 56324 297384
rect 56376 297412 56382 297424
rect 97074 297412 97080 297424
rect 56376 297384 97080 297412
rect 56376 297372 56382 297384
rect 97074 297372 97080 297384
rect 97132 297372 97138 297424
rect 97902 297372 97908 297424
rect 97960 297412 97966 297424
rect 145558 297412 145564 297424
rect 97960 297384 145564 297412
rect 97960 297372 97966 297384
rect 145558 297372 145564 297384
rect 145616 297372 145622 297424
rect 319530 297372 319536 297424
rect 319588 297412 319594 297424
rect 353938 297412 353944 297424
rect 319588 297384 353944 297412
rect 319588 297372 319594 297384
rect 353938 297372 353944 297384
rect 353996 297412 354002 297424
rect 388438 297412 388444 297424
rect 353996 297384 388444 297412
rect 353996 297372 354002 297384
rect 388438 297372 388444 297384
rect 388496 297372 388502 297424
rect 194502 297236 194508 297288
rect 194560 297276 194566 297288
rect 197354 297276 197360 297288
rect 194560 297248 197360 297276
rect 194560 297236 194566 297248
rect 197354 297236 197360 297248
rect 197412 297236 197418 297288
rect 112530 296964 112536 297016
rect 112588 297004 112594 297016
rect 124858 297004 124864 297016
rect 112588 296976 124864 297004
rect 112588 296964 112594 296976
rect 124858 296964 124864 296976
rect 124916 296964 124922 297016
rect 100662 296896 100668 296948
rect 100720 296936 100726 296948
rect 104802 296936 104808 296948
rect 100720 296908 104808 296936
rect 100720 296896 100726 296908
rect 104802 296896 104808 296908
rect 104860 296896 104866 296948
rect 116578 296896 116584 296948
rect 116636 296936 116642 296948
rect 144270 296936 144276 296948
rect 116636 296908 144276 296936
rect 116636 296896 116642 296908
rect 144270 296896 144276 296908
rect 144328 296896 144334 296948
rect 83550 296828 83556 296880
rect 83608 296868 83614 296880
rect 128998 296868 129004 296880
rect 83608 296840 129004 296868
rect 83608 296828 83614 296840
rect 128998 296828 129004 296840
rect 129056 296828 129062 296880
rect 90634 296760 90640 296812
rect 90692 296800 90698 296812
rect 147030 296800 147036 296812
rect 90692 296772 147036 296800
rect 90692 296760 90698 296772
rect 147030 296760 147036 296772
rect 147088 296760 147094 296812
rect 76466 296692 76472 296744
rect 76524 296732 76530 296744
rect 174630 296732 174636 296744
rect 76524 296704 174636 296732
rect 76524 296692 76530 296704
rect 174630 296692 174636 296704
rect 174688 296692 174694 296744
rect 59078 295944 59084 295996
rect 59136 295984 59142 295996
rect 73890 295984 73896 295996
rect 59136 295956 73896 295984
rect 59136 295944 59142 295956
rect 73890 295944 73896 295956
rect 73948 295944 73954 295996
rect 149790 295944 149796 295996
rect 149848 295984 149854 295996
rect 183002 295984 183008 295996
rect 149848 295956 183008 295984
rect 149848 295944 149854 295956
rect 183002 295944 183008 295956
rect 183060 295944 183066 295996
rect 107562 295672 107568 295724
rect 107620 295712 107626 295724
rect 140130 295712 140136 295724
rect 107620 295684 140136 295712
rect 107620 295672 107626 295684
rect 140130 295672 140136 295684
rect 140188 295672 140194 295724
rect 100938 295604 100944 295656
rect 100996 295644 101002 295656
rect 141510 295644 141516 295656
rect 100996 295616 141516 295644
rect 100996 295604 101002 295616
rect 141510 295604 141516 295616
rect 141568 295604 141574 295656
rect 113174 295536 113180 295588
rect 113232 295576 113238 295588
rect 113818 295576 113824 295588
rect 113232 295548 113824 295576
rect 113232 295536 113238 295548
rect 113818 295536 113824 295548
rect 113876 295576 113882 295588
rect 158070 295576 158076 295588
rect 113876 295548 158076 295576
rect 113876 295536 113882 295548
rect 158070 295536 158076 295548
rect 158128 295536 158134 295588
rect 115198 295468 115204 295520
rect 115256 295508 115262 295520
rect 115750 295508 115756 295520
rect 115256 295480 115756 295508
rect 115256 295468 115262 295480
rect 115750 295468 115756 295480
rect 115808 295508 115814 295520
rect 159634 295508 159640 295520
rect 115808 295480 159640 295508
rect 115808 295468 115814 295480
rect 159634 295468 159640 295480
rect 159692 295468 159698 295520
rect 68922 295400 68928 295452
rect 68980 295440 68986 295452
rect 134794 295440 134800 295452
rect 68980 295412 134800 295440
rect 68980 295400 68986 295412
rect 134794 295400 134800 295412
rect 134852 295400 134858 295452
rect 69106 295332 69112 295384
rect 69164 295372 69170 295384
rect 195698 295372 195704 295384
rect 69164 295344 195704 295372
rect 69164 295332 69170 295344
rect 195698 295332 195704 295344
rect 195756 295372 195762 295384
rect 197446 295372 197452 295384
rect 195756 295344 197452 295372
rect 195756 295332 195762 295344
rect 197446 295332 197452 295344
rect 197504 295332 197510 295384
rect 322474 295332 322480 295384
rect 322532 295372 322538 295384
rect 331306 295372 331312 295384
rect 322532 295344 331312 295372
rect 322532 295332 322538 295344
rect 331306 295332 331312 295344
rect 331364 295332 331370 295384
rect 71314 295264 71320 295316
rect 71372 295304 71378 295316
rect 75178 295304 75184 295316
rect 71372 295276 75184 295304
rect 71372 295264 71378 295276
rect 75178 295264 75184 295276
rect 75236 295264 75242 295316
rect 80330 295264 80336 295316
rect 80388 295304 80394 295316
rect 86218 295304 86224 295316
rect 80388 295276 86224 295304
rect 80388 295264 80394 295276
rect 86218 295264 86224 295276
rect 86276 295264 86282 295316
rect 117038 295264 117044 295316
rect 117096 295304 117102 295316
rect 123570 295304 123576 295316
rect 117096 295276 123576 295304
rect 117096 295264 117102 295276
rect 123570 295264 123576 295276
rect 123628 295264 123634 295316
rect 109310 294856 109316 294908
rect 109368 294896 109374 294908
rect 111058 294896 111064 294908
rect 109368 294868 111064 294896
rect 109368 294856 109374 294868
rect 111058 294856 111064 294868
rect 111116 294856 111122 294908
rect 111242 294856 111248 294908
rect 111300 294896 111306 294908
rect 124950 294896 124956 294908
rect 111300 294868 124956 294896
rect 111300 294856 111306 294868
rect 124950 294856 124956 294868
rect 125008 294856 125014 294908
rect 106734 294788 106740 294840
rect 106792 294828 106798 294840
rect 125042 294828 125048 294840
rect 106792 294800 125048 294828
rect 106792 294788 106798 294800
rect 125042 294788 125048 294800
rect 125100 294788 125106 294840
rect 72602 294720 72608 294772
rect 72660 294760 72666 294772
rect 87690 294760 87696 294772
rect 72660 294732 87696 294760
rect 72660 294720 72666 294732
rect 87690 294720 87696 294732
rect 87748 294720 87754 294772
rect 88702 294720 88708 294772
rect 88760 294760 88766 294772
rect 119430 294760 119436 294772
rect 88760 294732 119436 294760
rect 88760 294720 88766 294732
rect 119430 294720 119436 294732
rect 119488 294720 119494 294772
rect 56502 294652 56508 294704
rect 56560 294692 56566 294704
rect 111150 294692 111156 294704
rect 56560 294664 111156 294692
rect 56560 294652 56566 294664
rect 111150 294652 111156 294664
rect 111208 294652 111214 294704
rect 119614 294652 119620 294704
rect 119672 294692 119678 294704
rect 149238 294692 149244 294704
rect 119672 294664 149244 294692
rect 119672 294652 119678 294664
rect 149238 294652 149244 294664
rect 149296 294652 149302 294704
rect 88058 294584 88064 294636
rect 88116 294624 88122 294636
rect 107562 294624 107568 294636
rect 88116 294596 107568 294624
rect 88116 294584 88122 294596
rect 107562 294584 107568 294596
rect 107620 294584 107626 294636
rect 108022 294584 108028 294636
rect 108080 294624 108086 294636
rect 196618 294624 196624 294636
rect 108080 294596 196624 294624
rect 108080 294584 108086 294596
rect 196618 294584 196624 294596
rect 196676 294584 196682 294636
rect 322750 294584 322756 294636
rect 322808 294624 322814 294636
rect 420914 294624 420920 294636
rect 322808 294596 420920 294624
rect 322808 294584 322814 294596
rect 420914 294584 420920 294596
rect 420972 294584 420978 294636
rect 74626 294312 74632 294364
rect 74684 294352 74690 294364
rect 75454 294352 75460 294364
rect 74684 294324 75460 294352
rect 74684 294312 74690 294324
rect 75454 294312 75460 294324
rect 75512 294312 75518 294364
rect 77294 294312 77300 294364
rect 77352 294352 77358 294364
rect 78030 294352 78036 294364
rect 77352 294324 78036 294352
rect 77352 294312 77358 294324
rect 78030 294312 78036 294324
rect 78088 294312 78094 294364
rect 104894 294312 104900 294364
rect 104952 294352 104958 294364
rect 105814 294352 105820 294364
rect 104952 294324 105820 294352
rect 104952 294312 104958 294324
rect 105814 294312 105820 294324
rect 105872 294312 105878 294364
rect 77110 294244 77116 294296
rect 77168 294284 77174 294296
rect 79318 294284 79324 294296
rect 77168 294256 79324 294284
rect 77168 294244 77174 294256
rect 79318 294244 79324 294256
rect 79376 294244 79382 294296
rect 86126 294244 86132 294296
rect 86184 294284 86190 294296
rect 87598 294284 87604 294296
rect 86184 294256 87604 294284
rect 86184 294244 86190 294256
rect 87598 294244 87604 294256
rect 87656 294244 87662 294296
rect 55030 294108 55036 294160
rect 55088 294148 55094 294160
rect 74534 294148 74540 294160
rect 55088 294120 74540 294148
rect 55088 294108 55094 294120
rect 74534 294108 74540 294120
rect 74592 294108 74598 294160
rect 46750 294040 46756 294092
rect 46808 294080 46814 294092
rect 79686 294080 79692 294092
rect 46808 294052 79692 294080
rect 46808 294040 46814 294052
rect 79686 294040 79692 294052
rect 79744 294040 79750 294092
rect 110598 294040 110604 294092
rect 110656 294080 110662 294092
rect 117222 294080 117228 294092
rect 110656 294052 117228 294080
rect 110656 294040 110662 294052
rect 117222 294040 117228 294052
rect 117280 294040 117286 294092
rect 33778 293972 33784 294024
rect 33836 294012 33842 294024
rect 79410 294012 79416 294024
rect 33836 293984 79416 294012
rect 33836 293972 33842 293984
rect 79410 293972 79416 293984
rect 79468 293972 79474 294024
rect 84194 293972 84200 294024
rect 84252 294012 84258 294024
rect 180242 294012 180248 294024
rect 84252 293984 180248 294012
rect 84252 293972 84258 293984
rect 180242 293972 180248 293984
rect 180300 293972 180306 294024
rect 44082 293224 44088 293276
rect 44140 293264 44146 293276
rect 75914 293264 75920 293276
rect 44140 293236 75920 293264
rect 44140 293224 44146 293236
rect 75914 293224 75920 293236
rect 75972 293224 75978 293276
rect 322842 293224 322848 293276
rect 322900 293264 322906 293276
rect 324406 293264 324412 293276
rect 322900 293236 324412 293264
rect 322900 293224 322906 293236
rect 324406 293224 324412 293236
rect 324464 293264 324470 293276
rect 370498 293264 370504 293276
rect 324464 293236 370504 293264
rect 324464 293224 324470 293236
rect 370498 293224 370504 293236
rect 370556 293224 370562 293276
rect 2774 293156 2780 293208
rect 2832 293196 2838 293208
rect 4798 293196 4804 293208
rect 2832 293168 4804 293196
rect 2832 293156 2838 293168
rect 4798 293156 4804 293168
rect 4856 293156 4862 293208
rect 93210 292884 93216 292936
rect 93268 292924 93274 292936
rect 127618 292924 127624 292936
rect 93268 292896 127624 292924
rect 93268 292884 93274 292896
rect 127618 292884 127624 292896
rect 127676 292884 127682 292936
rect 53098 292816 53104 292868
rect 53156 292856 53162 292868
rect 92566 292856 92572 292868
rect 53156 292828 92572 292856
rect 53156 292816 53162 292828
rect 92566 292816 92572 292828
rect 92624 292856 92630 292868
rect 92934 292856 92940 292868
rect 92624 292828 92940 292856
rect 92624 292816 92630 292828
rect 92934 292816 92940 292828
rect 92992 292816 92998 292868
rect 93854 292816 93860 292868
rect 93912 292856 93918 292868
rect 130470 292856 130476 292868
rect 93912 292828 130476 292856
rect 93912 292816 93918 292828
rect 130470 292816 130476 292828
rect 130528 292816 130534 292868
rect 80974 292748 80980 292800
rect 81032 292788 81038 292800
rect 123478 292788 123484 292800
rect 81032 292760 123484 292788
rect 81032 292748 81038 292760
rect 123478 292748 123484 292760
rect 123536 292748 123542 292800
rect 73890 292680 73896 292732
rect 73948 292720 73954 292732
rect 124122 292720 124128 292732
rect 73948 292692 124128 292720
rect 73948 292680 73954 292692
rect 124122 292680 124128 292692
rect 124180 292680 124186 292732
rect 5442 292612 5448 292664
rect 5500 292652 5506 292664
rect 96430 292652 96436 292664
rect 5500 292624 96436 292652
rect 5500 292612 5506 292624
rect 96430 292612 96436 292624
rect 96488 292612 96494 292664
rect 98362 292612 98368 292664
rect 98420 292652 98426 292664
rect 98730 292652 98736 292664
rect 98420 292624 98736 292652
rect 98420 292612 98426 292624
rect 98730 292612 98736 292624
rect 98788 292652 98794 292664
rect 195330 292652 195336 292664
rect 98788 292624 195336 292652
rect 98788 292612 98794 292624
rect 195330 292612 195336 292624
rect 195388 292612 195394 292664
rect 68738 292544 68744 292596
rect 68796 292584 68802 292596
rect 196618 292584 196624 292596
rect 68796 292556 196624 292584
rect 68796 292544 68802 292556
rect 196618 292544 196624 292556
rect 196676 292544 196682 292596
rect 71682 292476 71688 292528
rect 71740 292516 71746 292528
rect 86402 292516 86408 292528
rect 71740 292488 86408 292516
rect 71740 292476 71746 292488
rect 86402 292476 86408 292488
rect 86460 292476 86466 292528
rect 121454 292476 121460 292528
rect 121512 292516 121518 292528
rect 152090 292516 152096 292528
rect 121512 292488 152096 292516
rect 121512 292476 121518 292488
rect 152090 292476 152096 292488
rect 152148 292516 152154 292528
rect 155402 292516 155408 292528
rect 152148 292488 155408 292516
rect 152148 292476 152154 292488
rect 155402 292476 155408 292488
rect 155460 292476 155466 292528
rect 118050 292408 118056 292460
rect 118108 292448 118114 292460
rect 124214 292448 124220 292460
rect 118108 292420 124220 292448
rect 118108 292408 118114 292420
rect 124214 292408 124220 292420
rect 124272 292408 124278 292460
rect 124122 292340 124128 292392
rect 124180 292380 124186 292392
rect 129826 292380 129832 292392
rect 124180 292352 129832 292380
rect 124180 292340 124186 292352
rect 129826 292340 129832 292352
rect 129884 292340 129890 292392
rect 89070 292108 89076 292120
rect 84166 292080 89076 292108
rect 66070 291796 66076 291848
rect 66128 291836 66134 291848
rect 84166 291836 84194 292080
rect 89070 292068 89076 292080
rect 89128 292068 89134 292120
rect 92290 291864 92296 291916
rect 92348 291904 92354 291916
rect 92348 291876 93854 291904
rect 92348 291864 92354 291876
rect 66128 291808 84194 291836
rect 66128 291796 66134 291808
rect 93826 291224 93854 291876
rect 117222 291864 117228 291916
rect 117280 291904 117286 291916
rect 117280 291876 122834 291904
rect 117280 291864 117286 291876
rect 122806 291836 122834 291876
rect 171870 291836 171876 291848
rect 122806 291808 171876 291836
rect 171870 291796 171876 291808
rect 171928 291796 171934 291848
rect 156690 291224 156696 291236
rect 93826 291196 156696 291224
rect 156690 291184 156696 291196
rect 156748 291184 156754 291236
rect 322474 291184 322480 291236
rect 322532 291224 322538 291236
rect 340138 291224 340144 291236
rect 322532 291196 340144 291224
rect 322532 291184 322538 291196
rect 340138 291184 340144 291196
rect 340196 291184 340202 291236
rect 38562 291116 38568 291168
rect 38620 291156 38626 291168
rect 67634 291156 67640 291168
rect 38620 291128 67640 291156
rect 38620 291116 38626 291128
rect 67634 291116 67640 291128
rect 67692 291116 67698 291168
rect 15838 290436 15844 290488
rect 15896 290476 15902 290488
rect 38562 290476 38568 290488
rect 15896 290448 38568 290476
rect 15896 290436 15902 290448
rect 38562 290436 38568 290448
rect 38620 290436 38626 290488
rect 129274 290436 129280 290488
rect 129332 290476 129338 290488
rect 142430 290476 142436 290488
rect 129332 290448 142436 290476
rect 129332 290436 129338 290448
rect 142430 290436 142436 290448
rect 142488 290436 142494 290488
rect 121546 289960 121552 290012
rect 121604 290000 121610 290012
rect 152550 290000 152556 290012
rect 121604 289972 152556 290000
rect 121604 289960 121610 289972
rect 152550 289960 152556 289972
rect 152608 289960 152614 290012
rect 121454 289892 121460 289944
rect 121512 289932 121518 289944
rect 173250 289932 173256 289944
rect 121512 289904 173256 289932
rect 121512 289892 121518 289904
rect 173250 289892 173256 289904
rect 173308 289892 173314 289944
rect 181622 289892 181628 289944
rect 181680 289932 181686 289944
rect 197446 289932 197452 289944
rect 181680 289904 197452 289932
rect 181680 289892 181686 289904
rect 197446 289892 197452 289904
rect 197504 289892 197510 289944
rect 42702 289824 42708 289876
rect 42760 289864 42766 289876
rect 67634 289864 67640 289876
rect 42760 289836 67640 289864
rect 42760 289824 42766 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 124030 289824 124036 289876
rect 124088 289864 124094 289876
rect 197998 289864 198004 289876
rect 124088 289836 198004 289864
rect 124088 289824 124094 289836
rect 197998 289824 198004 289836
rect 198056 289824 198062 289876
rect 121546 289756 121552 289808
rect 121604 289796 121610 289808
rect 195238 289796 195244 289808
rect 121604 289768 195244 289796
rect 121604 289756 121610 289768
rect 195238 289756 195244 289768
rect 195296 289756 195302 289808
rect 121454 289688 121460 289740
rect 121512 289728 121518 289740
rect 123754 289728 123760 289740
rect 121512 289700 123760 289728
rect 121512 289688 121518 289700
rect 123754 289688 123760 289700
rect 123812 289728 123818 289740
rect 124030 289728 124036 289740
rect 123812 289700 124036 289728
rect 123812 289688 123818 289700
rect 124030 289688 124036 289700
rect 124088 289688 124094 289740
rect 69014 289144 69020 289196
rect 69072 289184 69078 289196
rect 69750 289184 69756 289196
rect 69072 289156 69756 289184
rect 69072 289144 69078 289156
rect 69750 289144 69756 289156
rect 69808 289144 69814 289196
rect 123570 289076 123576 289128
rect 123628 289116 123634 289128
rect 128354 289116 128360 289128
rect 123628 289088 128360 289116
rect 123628 289076 123634 289088
rect 128354 289076 128360 289088
rect 128412 289116 128418 289128
rect 187694 289116 187700 289128
rect 128412 289088 187700 289116
rect 128412 289076 128418 289088
rect 187694 289076 187700 289088
rect 187752 289076 187758 289128
rect 187694 288396 187700 288448
rect 187752 288436 187758 288448
rect 188890 288436 188896 288448
rect 187752 288408 188896 288436
rect 187752 288396 187758 288408
rect 188890 288396 188896 288408
rect 188948 288436 188954 288448
rect 197446 288436 197452 288448
rect 188948 288408 197452 288436
rect 188948 288396 188954 288408
rect 197446 288396 197452 288408
rect 197504 288396 197510 288448
rect 340138 288396 340144 288448
rect 340196 288436 340202 288448
rect 495434 288436 495440 288448
rect 340196 288408 495440 288436
rect 340196 288396 340202 288408
rect 495434 288396 495440 288408
rect 495492 288396 495498 288448
rect 121454 288328 121460 288380
rect 121512 288368 121518 288380
rect 169110 288368 169116 288380
rect 121512 288340 169116 288368
rect 121512 288328 121518 288340
rect 169110 288328 169116 288340
rect 169168 288328 169174 288380
rect 121546 288260 121552 288312
rect 121604 288300 121610 288312
rect 142338 288300 142344 288312
rect 121604 288272 142344 288300
rect 121604 288260 121610 288272
rect 142338 288260 142344 288272
rect 142396 288300 142402 288312
rect 143442 288300 143448 288312
rect 142396 288272 143448 288300
rect 142396 288260 142402 288272
rect 143442 288260 143448 288272
rect 143500 288260 143506 288312
rect 143442 287648 143448 287700
rect 143500 287688 143506 287700
rect 163682 287688 163688 287700
rect 143500 287660 163688 287688
rect 143500 287648 143506 287660
rect 163682 287648 163688 287660
rect 163740 287648 163746 287700
rect 322750 287648 322756 287700
rect 322808 287688 322814 287700
rect 358722 287688 358728 287700
rect 322808 287660 358728 287688
rect 322808 287648 322814 287660
rect 358722 287648 358728 287660
rect 358780 287688 358786 287700
rect 506474 287688 506480 287700
rect 358780 287660 506480 287688
rect 358780 287648 358786 287660
rect 506474 287648 506480 287660
rect 506532 287648 506538 287700
rect 49418 287036 49424 287088
rect 49476 287076 49482 287088
rect 67634 287076 67640 287088
rect 49476 287048 67640 287076
rect 49476 287036 49482 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 52086 286968 52092 287020
rect 52144 287008 52150 287020
rect 67726 287008 67732 287020
rect 52144 286980 67732 287008
rect 52144 286968 52150 286980
rect 67726 286968 67732 286980
rect 67784 286968 67790 287020
rect 121546 286968 121552 287020
rect 121604 287008 121610 287020
rect 124214 287008 124220 287020
rect 121604 286980 124220 287008
rect 121604 286968 121610 286980
rect 124214 286968 124220 286980
rect 124272 286968 124278 287020
rect 121638 286900 121644 286952
rect 121696 286940 121702 286952
rect 124306 286940 124312 286952
rect 121696 286912 124312 286940
rect 121696 286900 121702 286912
rect 124306 286900 124312 286912
rect 124364 286900 124370 286952
rect 121454 286832 121460 286884
rect 121512 286872 121518 286884
rect 143718 286872 143724 286884
rect 121512 286844 143724 286872
rect 121512 286832 121518 286844
rect 143718 286832 143724 286844
rect 143776 286832 143782 286884
rect 66070 286288 66076 286340
rect 66128 286328 66134 286340
rect 68186 286328 68192 286340
rect 66128 286300 68192 286328
rect 66128 286288 66134 286300
rect 68186 286288 68192 286300
rect 68244 286288 68250 286340
rect 143718 286288 143724 286340
rect 143776 286328 143782 286340
rect 196802 286328 196808 286340
rect 143776 286300 196808 286328
rect 143776 286288 143782 286300
rect 196802 286288 196808 286300
rect 196860 286288 196866 286340
rect 52178 285676 52184 285728
rect 52236 285716 52242 285728
rect 67818 285716 67824 285728
rect 52236 285688 67824 285716
rect 52236 285676 52242 285688
rect 67818 285676 67824 285688
rect 67876 285676 67882 285728
rect 191190 285676 191196 285728
rect 191248 285716 191254 285728
rect 197446 285716 197452 285728
rect 191248 285688 197452 285716
rect 191248 285676 191254 285688
rect 197446 285676 197452 285688
rect 197504 285676 197510 285728
rect 322474 285676 322480 285728
rect 322532 285716 322538 285728
rect 329926 285716 329932 285728
rect 322532 285688 329932 285716
rect 322532 285676 322538 285688
rect 329926 285676 329932 285688
rect 329984 285676 329990 285728
rect 58986 285608 58992 285660
rect 59044 285648 59050 285660
rect 67634 285648 67640 285660
rect 59044 285620 67640 285648
rect 59044 285608 59050 285620
rect 67634 285608 67640 285620
rect 67692 285608 67698 285660
rect 121454 285608 121460 285660
rect 121512 285648 121518 285660
rect 193858 285648 193864 285660
rect 121512 285620 193864 285648
rect 121512 285608 121518 285620
rect 193858 285608 193864 285620
rect 193916 285608 193922 285660
rect 121546 285540 121552 285592
rect 121604 285580 121610 285592
rect 145006 285580 145012 285592
rect 121604 285552 145012 285580
rect 121604 285540 121610 285552
rect 145006 285540 145012 285552
rect 145064 285540 145070 285592
rect 121638 284996 121644 285048
rect 121696 285036 121702 285048
rect 158162 285036 158168 285048
rect 121696 285008 158168 285036
rect 121696 284996 121702 285008
rect 158162 284996 158168 285008
rect 158220 284996 158226 285048
rect 145006 284928 145012 284980
rect 145064 284968 145070 284980
rect 195974 284968 195980 284980
rect 145064 284940 195980 284968
rect 145064 284928 145070 284940
rect 195974 284928 195980 284940
rect 196032 284928 196038 284980
rect 38562 284316 38568 284368
rect 38620 284356 38626 284368
rect 67634 284356 67640 284368
rect 38620 284328 67640 284356
rect 38620 284316 38626 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 65518 284248 65524 284300
rect 65576 284288 65582 284300
rect 67726 284288 67732 284300
rect 65576 284260 67732 284288
rect 65576 284248 65582 284260
rect 67726 284248 67732 284260
rect 67784 284248 67790 284300
rect 121454 284248 121460 284300
rect 121512 284288 121518 284300
rect 131298 284288 131304 284300
rect 121512 284260 131304 284288
rect 121512 284248 121518 284260
rect 131298 284248 131304 284260
rect 131356 284248 131362 284300
rect 126238 284180 126244 284232
rect 126296 284220 126302 284232
rect 133598 284220 133604 284232
rect 126296 284192 133604 284220
rect 126296 284180 126302 284192
rect 133598 284180 133604 284192
rect 133656 284180 133662 284232
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 124950 282928 124956 282940
rect 121512 282900 124956 282928
rect 121512 282888 121518 282900
rect 124950 282888 124956 282900
rect 125008 282888 125014 282940
rect 132586 282888 132592 282940
rect 132644 282928 132650 282940
rect 133598 282928 133604 282940
rect 132644 282900 133604 282928
rect 132644 282888 132650 282900
rect 133598 282888 133604 282900
rect 133656 282928 133662 282940
rect 190270 282928 190276 282940
rect 133656 282900 190276 282928
rect 133656 282888 133662 282900
rect 190270 282888 190276 282900
rect 190328 282928 190334 282940
rect 197446 282928 197452 282940
rect 190328 282900 197452 282928
rect 190328 282888 190334 282900
rect 197446 282888 197452 282900
rect 197504 282888 197510 282940
rect 322474 282888 322480 282940
rect 322532 282928 322538 282940
rect 328546 282928 328552 282940
rect 322532 282900 328552 282928
rect 322532 282888 322538 282900
rect 328546 282888 328552 282900
rect 328604 282888 328610 282940
rect 41138 282820 41144 282872
rect 41196 282860 41202 282872
rect 67634 282860 67640 282872
rect 41196 282832 67640 282860
rect 41196 282820 41202 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 166442 281568 166448 281580
rect 121512 281540 166448 281568
rect 121512 281528 121518 281540
rect 166442 281528 166448 281540
rect 166500 281528 166506 281580
rect 180334 281528 180340 281580
rect 180392 281568 180398 281580
rect 197446 281568 197452 281580
rect 180392 281540 197452 281568
rect 180392 281528 180398 281540
rect 197446 281528 197452 281540
rect 197504 281528 197510 281580
rect 121546 281460 121552 281512
rect 121604 281500 121610 281512
rect 187050 281500 187056 281512
rect 121604 281472 187056 281500
rect 121604 281460 121610 281472
rect 187050 281460 187056 281472
rect 187108 281460 187114 281512
rect 178770 280780 178776 280832
rect 178828 280820 178834 280832
rect 186130 280820 186136 280832
rect 178828 280792 186136 280820
rect 178828 280780 178834 280792
rect 186130 280780 186136 280792
rect 186188 280780 186194 280832
rect 50890 280168 50896 280220
rect 50948 280208 50954 280220
rect 67634 280208 67640 280220
rect 50948 280180 67640 280208
rect 50948 280168 50954 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 129182 280208 129188 280220
rect 121512 280180 129188 280208
rect 121512 280168 121518 280180
rect 129182 280168 129188 280180
rect 129240 280168 129246 280220
rect 186130 280168 186136 280220
rect 186188 280208 186194 280220
rect 197446 280208 197452 280220
rect 186188 280180 197452 280208
rect 186188 280168 186194 280180
rect 197446 280168 197452 280180
rect 197504 280168 197510 280220
rect 322474 280168 322480 280220
rect 322532 280208 322538 280220
rect 335998 280208 336004 280220
rect 322532 280180 336004 280208
rect 322532 280168 322538 280180
rect 335998 280168 336004 280180
rect 336056 280168 336062 280220
rect 41414 280100 41420 280152
rect 41472 280140 41478 280152
rect 42610 280140 42616 280152
rect 41472 280112 42616 280140
rect 41472 280100 41478 280112
rect 42610 280100 42616 280112
rect 42668 280140 42674 280152
rect 67726 280140 67732 280152
rect 42668 280112 67732 280140
rect 42668 280100 42674 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 56226 280032 56232 280084
rect 56284 280072 56290 280084
rect 67634 280072 67640 280084
rect 56284 280044 67640 280072
rect 56284 280032 56290 280044
rect 67634 280032 67640 280044
rect 67692 280032 67698 280084
rect 29638 279420 29644 279472
rect 29696 279460 29702 279472
rect 41414 279460 41420 279472
rect 29696 279432 41420 279460
rect 29696 279420 29702 279432
rect 41414 279420 41420 279432
rect 41472 279420 41478 279472
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 192570 278780 192576 278792
rect 121512 278752 192576 278780
rect 121512 278740 121518 278752
rect 192570 278740 192576 278752
rect 192628 278740 192634 278792
rect 59078 278672 59084 278724
rect 59136 278712 59142 278724
rect 67634 278712 67640 278724
rect 59136 278684 67640 278712
rect 59136 278672 59142 278684
rect 67634 278672 67640 278684
rect 67692 278672 67698 278724
rect 152642 277992 152648 278044
rect 152700 278032 152706 278044
rect 183462 278032 183468 278044
rect 152700 278004 183468 278032
rect 152700 277992 152706 278004
rect 183462 277992 183468 278004
rect 183520 277992 183526 278044
rect 57790 277380 57796 277432
rect 57848 277420 57854 277432
rect 67634 277420 67640 277432
rect 57848 277392 67640 277420
rect 57848 277380 57854 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 121454 277380 121460 277432
rect 121512 277420 121518 277432
rect 142890 277420 142896 277432
rect 121512 277392 142896 277420
rect 121512 277380 121518 277392
rect 142890 277380 142896 277392
rect 142948 277380 142954 277432
rect 183462 277380 183468 277432
rect 183520 277420 183526 277432
rect 197446 277420 197452 277432
rect 183520 277392 197452 277420
rect 183520 277380 183526 277392
rect 197446 277380 197452 277392
rect 197504 277380 197510 277432
rect 122742 277312 122748 277364
rect 122800 277352 122806 277364
rect 160830 277352 160836 277364
rect 122800 277324 160836 277352
rect 122800 277312 122806 277324
rect 160830 277312 160836 277324
rect 160888 277312 160894 277364
rect 121454 277244 121460 277296
rect 121512 277284 121518 277296
rect 132494 277284 132500 277296
rect 121512 277256 132500 277284
rect 121512 277244 121518 277256
rect 132494 277244 132500 277256
rect 132552 277244 132558 277296
rect 321830 276632 321836 276684
rect 321888 276672 321894 276684
rect 493318 276672 493324 276684
rect 321888 276644 493324 276672
rect 321888 276632 321894 276644
rect 493318 276632 493324 276644
rect 493376 276632 493382 276684
rect 56134 276020 56140 276072
rect 56192 276060 56198 276072
rect 67726 276060 67732 276072
rect 56192 276032 67732 276060
rect 56192 276020 56198 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 160922 276060 160928 276072
rect 121512 276032 160928 276060
rect 121512 276020 121518 276032
rect 160922 276020 160928 276032
rect 160980 276020 160986 276072
rect 320818 276020 320824 276072
rect 320876 276060 320882 276072
rect 321830 276060 321836 276072
rect 320876 276032 321836 276060
rect 320876 276020 320882 276032
rect 321830 276020 321836 276032
rect 321888 276020 321894 276072
rect 56502 275952 56508 276004
rect 56560 275992 56566 276004
rect 67634 275992 67640 276004
rect 56560 275964 67640 275992
rect 56560 275952 56566 275964
rect 67634 275952 67640 275964
rect 67692 275952 67698 276004
rect 121546 274728 121552 274780
rect 121604 274768 121610 274780
rect 122098 274768 122104 274780
rect 121604 274740 122104 274768
rect 121604 274728 121610 274740
rect 122098 274728 122104 274740
rect 122156 274768 122162 274780
rect 144362 274768 144368 274780
rect 122156 274740 144368 274768
rect 122156 274728 122162 274740
rect 144362 274728 144368 274740
rect 144420 274728 144426 274780
rect 175090 274728 175096 274780
rect 175148 274768 175154 274780
rect 197446 274768 197452 274780
rect 175148 274740 197452 274768
rect 175148 274728 175154 274740
rect 197446 274728 197452 274740
rect 197504 274728 197510 274780
rect 53650 274660 53656 274712
rect 53708 274700 53714 274712
rect 67634 274700 67640 274712
rect 53708 274672 67640 274700
rect 53708 274660 53714 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121454 274660 121460 274712
rect 121512 274700 121518 274712
rect 187050 274700 187056 274712
rect 121512 274672 187056 274700
rect 121512 274660 121518 274672
rect 187050 274660 187056 274672
rect 187108 274660 187114 274712
rect 60458 274592 60464 274644
rect 60516 274632 60522 274644
rect 67726 274632 67732 274644
rect 60516 274604 67732 274632
rect 60516 274592 60522 274604
rect 67726 274592 67732 274604
rect 67784 274592 67790 274644
rect 322382 274592 322388 274644
rect 322440 274632 322446 274644
rect 339494 274632 339500 274644
rect 322440 274604 339500 274632
rect 322440 274592 322446 274604
rect 339494 274592 339500 274604
rect 339552 274592 339558 274644
rect 133230 273912 133236 273964
rect 133288 273952 133294 273964
rect 195238 273952 195244 273964
rect 133288 273924 195244 273952
rect 133288 273912 133294 273924
rect 195238 273912 195244 273924
rect 195296 273912 195302 273964
rect 339494 273912 339500 273964
rect 339552 273952 339558 273964
rect 382918 273952 382924 273964
rect 339552 273924 382924 273952
rect 339552 273912 339558 273924
rect 382918 273912 382924 273924
rect 382976 273912 382982 273964
rect 121454 273300 121460 273352
rect 121512 273340 121518 273352
rect 169110 273340 169116 273352
rect 121512 273312 169116 273340
rect 121512 273300 121518 273312
rect 169110 273300 169116 273312
rect 169168 273300 169174 273352
rect 43806 273232 43812 273284
rect 43864 273272 43870 273284
rect 67634 273272 67640 273284
rect 43864 273244 67640 273272
rect 43864 273232 43870 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 123754 273232 123760 273284
rect 123812 273272 123818 273284
rect 177942 273272 177948 273284
rect 123812 273244 177948 273272
rect 123812 273232 123818 273244
rect 177942 273232 177948 273244
rect 178000 273272 178006 273284
rect 197446 273272 197452 273284
rect 178000 273244 197452 273272
rect 178000 273232 178006 273244
rect 197446 273232 197452 273244
rect 197504 273232 197510 273284
rect 335998 273232 336004 273284
rect 336056 273272 336062 273284
rect 457438 273272 457444 273284
rect 336056 273244 457444 273272
rect 336056 273232 336062 273244
rect 457438 273232 457444 273244
rect 457496 273232 457502 273284
rect 121454 273164 121460 273216
rect 121512 273204 121518 273216
rect 133874 273204 133880 273216
rect 121512 273176 133880 273204
rect 121512 273164 121518 273176
rect 133874 273164 133880 273176
rect 133932 273164 133938 273216
rect 52086 271872 52092 271924
rect 52144 271912 52150 271924
rect 67634 271912 67640 271924
rect 52144 271884 67640 271912
rect 52144 271872 52150 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 417418 271872 417424 271924
rect 417476 271912 417482 271924
rect 419534 271912 419540 271924
rect 417476 271884 419540 271912
rect 417476 271872 417482 271884
rect 419534 271872 419540 271884
rect 419592 271912 419598 271924
rect 580166 271912 580172 271924
rect 419592 271884 580172 271912
rect 419592 271872 419598 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 53558 271804 53564 271856
rect 53616 271844 53622 271856
rect 67726 271844 67732 271856
rect 53616 271816 67732 271844
rect 53616 271804 53622 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 124950 271124 124956 271176
rect 125008 271164 125014 271176
rect 197446 271164 197452 271176
rect 125008 271136 197452 271164
rect 125008 271124 125014 271136
rect 197446 271124 197452 271136
rect 197504 271124 197510 271176
rect 65978 270512 65984 270564
rect 66036 270552 66042 270564
rect 68094 270552 68100 270564
rect 66036 270524 68100 270552
rect 66036 270512 66042 270524
rect 68094 270512 68100 270524
rect 68152 270512 68158 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 174538 270552 174544 270564
rect 121512 270524 174544 270552
rect 121512 270512 121518 270524
rect 174538 270512 174544 270524
rect 174596 270512 174602 270564
rect 121454 269628 121460 269680
rect 121512 269668 121518 269680
rect 124950 269668 124956 269680
rect 121512 269640 124956 269668
rect 121512 269628 121518 269640
rect 124950 269628 124956 269640
rect 125008 269628 125014 269680
rect 176010 269288 176016 269340
rect 176068 269328 176074 269340
rect 180334 269328 180340 269340
rect 176068 269300 180340 269328
rect 176068 269288 176074 269300
rect 180334 269288 180340 269300
rect 180392 269288 180398 269340
rect 59078 269084 59084 269136
rect 59136 269124 59142 269136
rect 67634 269124 67640 269136
rect 59136 269096 67640 269124
rect 59136 269084 59142 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121454 269084 121460 269136
rect 121512 269124 121518 269136
rect 133230 269124 133236 269136
rect 121512 269096 133236 269124
rect 121512 269084 121518 269096
rect 133230 269084 133236 269096
rect 133288 269084 133294 269136
rect 322842 269084 322848 269136
rect 322900 269124 322906 269136
rect 327258 269124 327264 269136
rect 322900 269096 327264 269124
rect 322900 269084 322906 269096
rect 327258 269084 327264 269096
rect 327316 269084 327322 269136
rect 47854 269016 47860 269068
rect 47912 269056 47918 269068
rect 48222 269056 48228 269068
rect 47912 269028 48228 269056
rect 47912 269016 47918 269028
rect 48222 269016 48228 269028
rect 48280 269016 48286 269068
rect 121546 269016 121552 269068
rect 121604 269056 121610 269068
rect 150434 269056 150440 269068
rect 121604 269028 150440 269056
rect 121604 269016 121610 269028
rect 150434 269016 150440 269028
rect 150492 269016 150498 269068
rect 43898 268404 43904 268456
rect 43956 268444 43962 268456
rect 55214 268444 55220 268456
rect 43956 268416 55220 268444
rect 43956 268404 43962 268416
rect 55214 268404 55220 268416
rect 55272 268404 55278 268456
rect 48222 268336 48228 268388
rect 48280 268376 48286 268388
rect 67634 268376 67640 268388
rect 48280 268348 67640 268376
rect 48280 268336 48286 268348
rect 67634 268336 67640 268348
rect 67692 268336 67698 268388
rect 134794 268336 134800 268388
rect 134852 268376 134858 268388
rect 134852 268348 180794 268376
rect 134852 268336 134858 268348
rect 180766 268240 180794 268348
rect 194318 268240 194324 268252
rect 180766 268212 194324 268240
rect 194318 268200 194324 268212
rect 194376 268240 194382 268252
rect 197446 268240 197452 268252
rect 194376 268212 197452 268240
rect 194376 268200 194382 268212
rect 197446 268200 197452 268212
rect 197504 268200 197510 268252
rect 121454 267724 121460 267776
rect 121512 267764 121518 267776
rect 134702 267764 134708 267776
rect 121512 267736 134708 267764
rect 121512 267724 121518 267736
rect 134702 267724 134708 267736
rect 134760 267724 134766 267776
rect 150434 267724 150440 267776
rect 150492 267764 150498 267776
rect 154022 267764 154028 267776
rect 150492 267736 154028 267764
rect 150492 267724 150498 267736
rect 154022 267724 154028 267736
rect 154080 267724 154086 267776
rect 45370 267656 45376 267708
rect 45428 267696 45434 267708
rect 67726 267696 67732 267708
rect 45428 267668 67732 267696
rect 45428 267656 45434 267668
rect 67726 267656 67732 267668
rect 67784 267656 67790 267708
rect 322474 267656 322480 267708
rect 322532 267696 322538 267708
rect 335354 267696 335360 267708
rect 322532 267668 335360 267696
rect 322532 267656 322538 267668
rect 335354 267656 335360 267668
rect 335412 267696 335418 267708
rect 336642 267696 336648 267708
rect 335412 267668 336648 267696
rect 335412 267656 335418 267668
rect 336642 267656 336648 267668
rect 336700 267656 336706 267708
rect 55214 266976 55220 267028
rect 55272 267016 55278 267028
rect 56318 267016 56324 267028
rect 55272 266988 56324 267016
rect 55272 266976 55278 266988
rect 56318 266976 56324 266988
rect 56376 267016 56382 267028
rect 67634 267016 67640 267028
rect 56376 266988 67640 267016
rect 56376 266976 56382 266988
rect 67634 266976 67640 266988
rect 67692 266976 67698 267028
rect 336642 266976 336648 267028
rect 336700 267016 336706 267028
rect 499758 267016 499764 267028
rect 336700 266988 499764 267016
rect 336700 266976 336706 266988
rect 499758 266976 499764 266988
rect 499816 266976 499822 267028
rect 121454 266432 121460 266484
rect 121512 266472 121518 266484
rect 144454 266472 144460 266484
rect 121512 266444 144460 266472
rect 121512 266432 121518 266444
rect 144454 266432 144460 266444
rect 144512 266432 144518 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 50338 266404 50344 266416
rect 3108 266376 50344 266404
rect 3108 266364 3114 266376
rect 50338 266364 50344 266376
rect 50396 266364 50402 266416
rect 121546 266364 121552 266416
rect 121604 266404 121610 266416
rect 158162 266404 158168 266416
rect 121604 266376 158168 266404
rect 121604 266364 121610 266376
rect 158162 266364 158168 266376
rect 158220 266364 158226 266416
rect 179414 266364 179420 266416
rect 179472 266404 179478 266416
rect 180702 266404 180708 266416
rect 179472 266376 180708 266404
rect 179472 266364 179478 266376
rect 180702 266364 180708 266376
rect 180760 266404 180766 266416
rect 197354 266404 197360 266416
rect 180760 266376 197360 266404
rect 180760 266364 180766 266376
rect 197354 266364 197360 266376
rect 197412 266364 197418 266416
rect 54846 266296 54852 266348
rect 54904 266336 54910 266348
rect 67634 266336 67640 266348
rect 54904 266308 67640 266336
rect 54904 266296 54910 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 145650 265044 145656 265056
rect 121512 265016 145656 265044
rect 121512 265004 121518 265016
rect 145650 265004 145656 265016
rect 145708 265004 145714 265056
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 151354 264976 151360 264988
rect 121604 264948 151360 264976
rect 121604 264936 121610 264948
rect 151354 264936 151360 264948
rect 151412 264936 151418 264988
rect 322474 264936 322480 264988
rect 322532 264976 322538 264988
rect 330018 264976 330024 264988
rect 322532 264948 330024 264976
rect 322532 264936 322538 264948
rect 330018 264936 330024 264948
rect 330076 264936 330082 264988
rect 121454 264868 121460 264920
rect 121512 264908 121518 264920
rect 125594 264908 125600 264920
rect 121512 264880 125600 264908
rect 121512 264868 121518 264880
rect 125594 264868 125600 264880
rect 125652 264868 125658 264920
rect 21358 264188 21364 264240
rect 21416 264228 21422 264240
rect 43990 264228 43996 264240
rect 21416 264200 43996 264228
rect 21416 264188 21422 264200
rect 43990 264188 43996 264200
rect 44048 264228 44054 264240
rect 53834 264228 53840 264240
rect 44048 264200 53840 264228
rect 44048 264188 44054 264200
rect 53834 264188 53840 264200
rect 53892 264188 53898 264240
rect 124122 264188 124128 264240
rect 124180 264228 124186 264240
rect 183370 264228 183376 264240
rect 124180 264200 183376 264228
rect 124180 264188 124186 264200
rect 183370 264188 183376 264200
rect 183428 264188 183434 264240
rect 60458 263644 60464 263696
rect 60516 263684 60522 263696
rect 67634 263684 67640 263696
rect 60516 263656 67640 263684
rect 60516 263644 60522 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 53834 263576 53840 263628
rect 53892 263616 53898 263628
rect 54846 263616 54852 263628
rect 53892 263588 54852 263616
rect 53892 263576 53898 263588
rect 54846 263576 54852 263588
rect 54904 263616 54910 263628
rect 67726 263616 67732 263628
rect 54904 263588 67732 263616
rect 54904 263576 54910 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121454 263576 121460 263628
rect 121512 263616 121518 263628
rect 138750 263616 138756 263628
rect 121512 263588 138756 263616
rect 121512 263576 121518 263588
rect 138750 263576 138756 263588
rect 138808 263576 138814 263628
rect 175090 263576 175096 263628
rect 175148 263616 175154 263628
rect 178770 263616 178776 263628
rect 175148 263588 178776 263616
rect 175148 263576 175154 263588
rect 178770 263576 178776 263588
rect 178828 263576 178834 263628
rect 183370 263576 183376 263628
rect 183428 263616 183434 263628
rect 197354 263616 197360 263628
rect 183428 263588 197360 263616
rect 183428 263576 183434 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 360286 263576 360292 263628
rect 360344 263616 360350 263628
rect 361482 263616 361488 263628
rect 360344 263588 361488 263616
rect 360344 263576 360350 263588
rect 361482 263576 361488 263588
rect 361540 263616 361546 263628
rect 490558 263616 490564 263628
rect 361540 263588 490564 263616
rect 361540 263576 361546 263588
rect 490558 263576 490564 263588
rect 490616 263576 490622 263628
rect 57698 263508 57704 263560
rect 57756 263548 57762 263560
rect 67634 263548 67640 263560
rect 57756 263520 67640 263548
rect 57756 263508 57762 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121546 263508 121552 263560
rect 121604 263548 121610 263560
rect 175108 263548 175136 263576
rect 121604 263520 175136 263548
rect 121604 263508 121610 263520
rect 121454 263440 121460 263492
rect 121512 263480 121518 263492
rect 138106 263480 138112 263492
rect 121512 263452 138112 263480
rect 121512 263440 121518 263452
rect 138106 263440 138112 263452
rect 138164 263440 138170 263492
rect 138106 263032 138112 263084
rect 138164 263072 138170 263084
rect 141602 263072 141608 263084
rect 138164 263044 141608 263072
rect 138164 263032 138170 263044
rect 141602 263032 141608 263044
rect 141660 263032 141666 263084
rect 334342 262828 334348 262880
rect 334400 262868 334406 262880
rect 360286 262868 360292 262880
rect 334400 262840 360292 262868
rect 334400 262828 334406 262840
rect 360286 262828 360292 262840
rect 360344 262828 360350 262880
rect 60366 262216 60372 262268
rect 60424 262256 60430 262268
rect 67634 262256 67640 262268
rect 60424 262228 67640 262256
rect 60424 262216 60430 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 128262 262256 128268 262268
rect 127820 262228 128268 262256
rect 64506 262148 64512 262200
rect 64564 262188 64570 262200
rect 67818 262188 67824 262200
rect 64564 262160 67824 262188
rect 64564 262148 64570 262160
rect 67818 262148 67824 262160
rect 67876 262148 67882 262200
rect 121546 262148 121552 262200
rect 121604 262188 121610 262200
rect 127820 262188 127848 262228
rect 128262 262216 128268 262228
rect 128320 262256 128326 262268
rect 152642 262256 152648 262268
rect 128320 262228 152648 262256
rect 128320 262216 128326 262228
rect 152642 262216 152648 262228
rect 152700 262216 152706 262268
rect 322474 262216 322480 262268
rect 322532 262256 322538 262268
rect 334066 262256 334072 262268
rect 322532 262228 334072 262256
rect 322532 262216 322538 262228
rect 334066 262216 334072 262228
rect 334124 262256 334130 262268
rect 334342 262256 334348 262268
rect 334124 262228 334348 262256
rect 334124 262216 334130 262228
rect 334342 262216 334348 262228
rect 334400 262216 334406 262268
rect 121604 262160 127848 262188
rect 121604 262148 121610 262160
rect 121454 262012 121460 262064
rect 121512 262052 121518 262064
rect 123754 262052 123760 262064
rect 121512 262024 123760 262052
rect 121512 262012 121518 262024
rect 123754 262012 123760 262024
rect 123812 262012 123818 262064
rect 123662 261468 123668 261520
rect 123720 261508 123726 261520
rect 138014 261508 138020 261520
rect 123720 261480 138020 261508
rect 123720 261468 123726 261480
rect 138014 261468 138020 261480
rect 138072 261508 138078 261520
rect 186314 261508 186320 261520
rect 138072 261480 186320 261508
rect 138072 261468 138078 261480
rect 186314 261468 186320 261480
rect 186372 261468 186378 261520
rect 56502 260856 56508 260908
rect 56560 260896 56566 260908
rect 67726 260896 67732 260908
rect 56560 260868 67732 260896
rect 56560 260856 56566 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 186314 260856 186320 260908
rect 186372 260896 186378 260908
rect 187510 260896 187516 260908
rect 186372 260868 187516 260896
rect 186372 260856 186378 260868
rect 187510 260856 187516 260868
rect 187568 260896 187574 260908
rect 197354 260896 197360 260908
rect 187568 260868 197360 260896
rect 187568 260856 187574 260868
rect 197354 260856 197360 260868
rect 197412 260856 197418 260908
rect 56410 260788 56416 260840
rect 56468 260828 56474 260840
rect 67634 260828 67640 260840
rect 56468 260800 67640 260828
rect 56468 260788 56474 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 150434 260828 150440 260840
rect 121512 260800 150440 260828
rect 121512 260788 121518 260800
rect 150434 260788 150440 260800
rect 150492 260788 150498 260840
rect 150434 260108 150440 260160
rect 150492 260148 150498 260160
rect 151722 260148 151728 260160
rect 150492 260120 151728 260148
rect 150492 260108 150498 260120
rect 151722 260108 151728 260120
rect 151780 260148 151786 260160
rect 160830 260148 160836 260160
rect 151780 260120 160836 260148
rect 151780 260108 151786 260120
rect 160830 260108 160836 260120
rect 160888 260108 160894 260160
rect 370498 260108 370504 260160
rect 370556 260148 370562 260160
rect 520918 260148 520924 260160
rect 370556 260120 520924 260148
rect 370556 260108 370562 260120
rect 520918 260108 520924 260120
rect 520976 260108 520982 260160
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 131758 259468 131764 259480
rect 121512 259440 131764 259468
rect 121512 259428 121518 259440
rect 131758 259428 131764 259440
rect 131816 259428 131822 259480
rect 194410 259428 194416 259480
rect 194468 259468 194474 259480
rect 197354 259468 197360 259480
rect 194468 259440 197360 259468
rect 194468 259428 194474 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 322474 259428 322480 259480
rect 322532 259468 322538 259480
rect 327350 259468 327356 259480
rect 322532 259440 327356 259468
rect 322532 259428 322538 259440
rect 327350 259428 327356 259440
rect 327408 259428 327414 259480
rect 121546 259360 121552 259412
rect 121604 259400 121610 259412
rect 136634 259400 136640 259412
rect 121604 259372 136640 259400
rect 121604 259360 121610 259372
rect 136634 259360 136640 259372
rect 136692 259400 136698 259412
rect 137094 259400 137100 259412
rect 136692 259372 137100 259400
rect 136692 259360 136698 259372
rect 137094 259360 137100 259372
rect 137152 259360 137158 259412
rect 137094 258680 137100 258732
rect 137152 258720 137158 258732
rect 161014 258720 161020 258732
rect 137152 258692 161020 258720
rect 137152 258680 137158 258692
rect 161014 258680 161020 258692
rect 161072 258680 161078 258732
rect 188798 258680 188804 258732
rect 188856 258720 188862 258732
rect 194410 258720 194416 258732
rect 188856 258692 194416 258720
rect 188856 258680 188862 258692
rect 194410 258680 194416 258692
rect 194468 258680 194474 258732
rect 520918 258680 520924 258732
rect 520976 258720 520982 258732
rect 579982 258720 579988 258732
rect 520976 258692 579988 258720
rect 520976 258680 520982 258692
rect 579982 258680 579988 258692
rect 580040 258680 580046 258732
rect 66070 258136 66076 258188
rect 66128 258176 66134 258188
rect 67634 258176 67640 258188
rect 66128 258148 67640 258176
rect 66128 258136 66134 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 322842 258136 322848 258188
rect 322900 258176 322906 258188
rect 324498 258176 324504 258188
rect 322900 258148 324504 258176
rect 322900 258136 322906 258148
rect 324498 258136 324504 258148
rect 324556 258176 324562 258188
rect 324556 258148 325694 258176
rect 324556 258136 324562 258148
rect 57698 258068 57704 258120
rect 57756 258108 57762 258120
rect 67726 258108 67732 258120
rect 57756 258080 67732 258108
rect 57756 258068 57762 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121638 258068 121644 258120
rect 121696 258108 121702 258120
rect 137462 258108 137468 258120
rect 121696 258080 137468 258108
rect 121696 258068 121702 258080
rect 137462 258068 137468 258080
rect 137520 258068 137526 258120
rect 325666 258108 325694 258148
rect 393958 258108 393964 258120
rect 325666 258080 393964 258108
rect 393958 258068 393964 258080
rect 394016 258068 394022 258120
rect 34238 258000 34244 258052
rect 34296 258040 34302 258052
rect 67634 258040 67640 258052
rect 34296 258012 67640 258040
rect 34296 258000 34302 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 121454 258000 121460 258052
rect 121512 258040 121518 258052
rect 154574 258040 154580 258052
rect 121512 258012 154580 258040
rect 121512 258000 121518 258012
rect 154574 258000 154580 258012
rect 154632 258000 154638 258052
rect 14458 257320 14464 257372
rect 14516 257360 14522 257372
rect 34238 257360 34244 257372
rect 14516 257332 34244 257360
rect 14516 257320 14522 257332
rect 34238 257320 34244 257332
rect 34296 257320 34302 257372
rect 53558 256708 53564 256760
rect 53616 256748 53622 256760
rect 67634 256748 67640 256760
rect 53616 256720 67640 256748
rect 53616 256708 53622 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 126238 256748 126244 256760
rect 121604 256720 126244 256748
rect 121604 256708 121610 256720
rect 126238 256708 126244 256720
rect 126296 256708 126302 256760
rect 133874 256708 133880 256760
rect 133932 256748 133938 256760
rect 197354 256748 197360 256760
rect 133932 256720 197360 256748
rect 133932 256708 133938 256720
rect 197354 256708 197360 256720
rect 197412 256708 197418 256760
rect 121454 256640 121460 256692
rect 121512 256680 121518 256692
rect 136726 256680 136732 256692
rect 121512 256652 136732 256680
rect 121512 256640 121518 256652
rect 136726 256640 136732 256652
rect 136784 256640 136790 256692
rect 136726 256028 136732 256080
rect 136784 256068 136790 256080
rect 169202 256068 169208 256080
rect 136784 256040 169208 256068
rect 136784 256028 136790 256040
rect 169202 256028 169208 256040
rect 169260 256028 169266 256080
rect 141602 255960 141608 256012
rect 141660 256000 141666 256012
rect 181806 256000 181812 256012
rect 141660 255972 181812 256000
rect 141660 255960 141666 255972
rect 181806 255960 181812 255972
rect 181864 255960 181870 256012
rect 63126 255280 63132 255332
rect 63184 255320 63190 255332
rect 67634 255320 67640 255332
rect 63184 255292 67640 255320
rect 63184 255280 63190 255292
rect 67634 255280 67640 255292
rect 67692 255280 67698 255332
rect 181806 255280 181812 255332
rect 181864 255320 181870 255332
rect 182082 255320 182088 255332
rect 181864 255292 182088 255320
rect 181864 255280 181870 255292
rect 182082 255280 182088 255292
rect 182140 255320 182146 255332
rect 197354 255320 197360 255332
rect 182140 255292 197360 255320
rect 182140 255280 182146 255292
rect 197354 255280 197360 255292
rect 197412 255280 197418 255332
rect 50706 255212 50712 255264
rect 50764 255252 50770 255264
rect 67726 255252 67732 255264
rect 50764 255224 67732 255252
rect 50764 255212 50770 255224
rect 67726 255212 67732 255224
rect 67784 255212 67790 255264
rect 52270 255144 52276 255196
rect 52328 255184 52334 255196
rect 67634 255184 67640 255196
rect 52328 255156 67640 255184
rect 52328 255144 52334 255156
rect 67634 255144 67640 255156
rect 67692 255144 67698 255196
rect 122098 254600 122104 254652
rect 122156 254640 122162 254652
rect 130378 254640 130384 254652
rect 122156 254612 130384 254640
rect 122156 254600 122162 254612
rect 130378 254600 130384 254612
rect 130436 254600 130442 254652
rect 122466 254532 122472 254584
rect 122524 254572 122530 254584
rect 167730 254572 167736 254584
rect 122524 254544 167736 254572
rect 122524 254532 122530 254544
rect 167730 254532 167736 254544
rect 167788 254532 167794 254584
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 142982 253960 142988 253972
rect 121512 253932 142988 253960
rect 121512 253920 121518 253932
rect 142982 253920 142988 253932
rect 143040 253920 143046 253972
rect 47670 253852 47676 253904
rect 47728 253892 47734 253904
rect 48038 253892 48044 253904
rect 47728 253864 48044 253892
rect 47728 253852 47734 253864
rect 48038 253852 48044 253864
rect 48096 253892 48102 253904
rect 67634 253892 67640 253904
rect 48096 253864 67640 253892
rect 48096 253852 48102 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 63218 253784 63224 253836
rect 63276 253824 63282 253836
rect 67726 253824 67732 253836
rect 63276 253796 67732 253824
rect 63276 253784 63282 253796
rect 67726 253784 67732 253796
rect 67784 253784 67790 253836
rect 32398 253172 32404 253224
rect 32456 253212 32462 253224
rect 47670 253212 47676 253224
rect 32456 253184 47676 253212
rect 32456 253172 32462 253184
rect 47670 253172 47676 253184
rect 47728 253172 47734 253224
rect 121454 252628 121460 252680
rect 121512 252668 121518 252680
rect 155494 252668 155500 252680
rect 121512 252640 155500 252668
rect 121512 252628 121518 252640
rect 155494 252628 155500 252640
rect 155552 252628 155558 252680
rect 120810 252560 120816 252612
rect 120868 252600 120874 252612
rect 191742 252600 191748 252612
rect 120868 252572 191748 252600
rect 120868 252560 120874 252572
rect 191742 252560 191748 252572
rect 191800 252600 191806 252612
rect 197354 252600 197360 252612
rect 191800 252572 197360 252600
rect 191800 252560 191806 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 322842 252560 322848 252612
rect 322900 252600 322906 252612
rect 324406 252600 324412 252612
rect 322900 252572 324412 252600
rect 322900 252560 322906 252572
rect 324406 252560 324412 252572
rect 324464 252560 324470 252612
rect 121454 252492 121460 252544
rect 121512 252532 121518 252544
rect 155954 252532 155960 252544
rect 121512 252504 155960 252532
rect 121512 252492 121518 252504
rect 155954 252492 155960 252504
rect 156012 252492 156018 252544
rect 192846 251608 192852 251660
rect 192904 251648 192910 251660
rect 196710 251648 196716 251660
rect 192904 251620 196716 251648
rect 192904 251608 192910 251620
rect 196710 251608 196716 251620
rect 196768 251608 196774 251660
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 184290 251240 184296 251252
rect 121512 251212 184296 251240
rect 121512 251200 121518 251212
rect 184290 251200 184296 251212
rect 184348 251200 184354 251252
rect 66162 251132 66168 251184
rect 66220 251172 66226 251184
rect 67634 251172 67640 251184
rect 66220 251144 67640 251172
rect 66220 251132 66226 251144
rect 67634 251132 67640 251144
rect 67692 251132 67698 251184
rect 167914 250452 167920 250504
rect 167972 250492 167978 250504
rect 194410 250492 194416 250504
rect 167972 250464 194416 250492
rect 167972 250452 167978 250464
rect 194410 250452 194416 250464
rect 194468 250452 194474 250504
rect 194410 249908 194416 249960
rect 194468 249948 194474 249960
rect 197354 249948 197360 249960
rect 194468 249920 197360 249948
rect 194468 249908 194474 249920
rect 197354 249908 197360 249920
rect 197412 249908 197418 249960
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 133322 249812 133328 249824
rect 121512 249784 133328 249812
rect 121512 249772 121518 249784
rect 133322 249772 133328 249784
rect 133380 249772 133386 249824
rect 140222 249812 140228 249824
rect 139412 249784 140228 249812
rect 121546 249704 121552 249756
rect 121604 249744 121610 249756
rect 139412 249744 139440 249784
rect 140222 249772 140228 249784
rect 140280 249812 140286 249824
rect 156782 249812 156788 249824
rect 140280 249784 156788 249812
rect 140280 249772 140286 249784
rect 156782 249772 156788 249784
rect 156840 249772 156846 249824
rect 121604 249716 139440 249744
rect 121604 249704 121610 249716
rect 121454 249636 121460 249688
rect 121512 249676 121518 249688
rect 129090 249676 129096 249688
rect 121512 249648 129096 249676
rect 121512 249636 121518 249648
rect 129090 249636 129096 249648
rect 129148 249636 129154 249688
rect 35710 249024 35716 249076
rect 35768 249064 35774 249076
rect 56226 249064 56232 249076
rect 35768 249036 56232 249064
rect 35768 249024 35774 249036
rect 56226 249024 56232 249036
rect 56284 249024 56290 249076
rect 195330 248956 195336 249008
rect 195388 248996 195394 249008
rect 197354 248996 197360 249008
rect 195388 248968 197360 248996
rect 195388 248956 195394 248968
rect 197354 248956 197360 248968
rect 197412 248956 197418 249008
rect 56226 248412 56232 248464
rect 56284 248452 56290 248464
rect 67634 248452 67640 248464
rect 56284 248424 67640 248452
rect 56284 248412 56290 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 322474 248412 322480 248464
rect 322532 248452 322538 248464
rect 335446 248452 335452 248464
rect 322532 248424 335452 248452
rect 322532 248412 322538 248424
rect 335446 248412 335452 248424
rect 335504 248452 335510 248464
rect 434714 248452 434720 248464
rect 335504 248424 434720 248452
rect 335504 248412 335510 248424
rect 434714 248412 434720 248424
rect 434772 248412 434778 248464
rect 121454 247120 121460 247172
rect 121512 247160 121518 247172
rect 137370 247160 137376 247172
rect 121512 247132 137376 247160
rect 121512 247120 121518 247132
rect 137370 247120 137376 247132
rect 137428 247120 137434 247172
rect 66162 247052 66168 247104
rect 66220 247092 66226 247104
rect 67634 247092 67640 247104
rect 66220 247064 67640 247092
rect 66220 247052 66226 247064
rect 67634 247052 67640 247064
rect 67692 247052 67698 247104
rect 121546 247052 121552 247104
rect 121604 247092 121610 247104
rect 178954 247092 178960 247104
rect 121604 247064 178960 247092
rect 121604 247052 121610 247064
rect 178954 247052 178960 247064
rect 179012 247052 179018 247104
rect 135898 246508 135904 246560
rect 135956 246548 135962 246560
rect 136634 246548 136640 246560
rect 135956 246520 136640 246548
rect 135956 246508 135962 246520
rect 136634 246508 136640 246520
rect 136692 246508 136698 246560
rect 121454 246168 121460 246220
rect 121512 246208 121518 246220
rect 125042 246208 125048 246220
rect 121512 246180 125048 246208
rect 121512 246168 121518 246180
rect 125042 246168 125048 246180
rect 125100 246168 125106 246220
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 151262 245732 151268 245744
rect 121604 245704 151268 245732
rect 121604 245692 121610 245704
rect 151262 245692 151268 245704
rect 151320 245692 151326 245744
rect 136634 245624 136640 245676
rect 136692 245664 136698 245676
rect 195882 245664 195888 245676
rect 136692 245636 195888 245664
rect 136692 245624 136698 245636
rect 195882 245624 195888 245636
rect 195940 245664 195946 245676
rect 198090 245664 198096 245676
rect 195940 245636 198096 245664
rect 195940 245624 195946 245636
rect 198090 245624 198096 245636
rect 198148 245624 198154 245676
rect 322474 245624 322480 245676
rect 322532 245664 322538 245676
rect 332686 245664 332692 245676
rect 322532 245636 332692 245664
rect 322532 245624 322538 245636
rect 332686 245624 332692 245636
rect 332744 245664 332750 245676
rect 374638 245664 374644 245676
rect 332744 245636 374644 245664
rect 332744 245624 332750 245636
rect 374638 245624 374644 245636
rect 374696 245624 374702 245676
rect 54938 245556 54944 245608
rect 54996 245596 55002 245608
rect 67634 245596 67640 245608
rect 54996 245568 67640 245596
rect 54996 245556 55002 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 53374 245488 53380 245540
rect 53432 245528 53438 245540
rect 67358 245528 67364 245540
rect 53432 245500 67364 245528
rect 53432 245488 53438 245500
rect 67358 245488 67364 245500
rect 67416 245488 67422 245540
rect 195330 245012 195336 245064
rect 195388 245052 195394 245064
rect 196710 245052 196716 245064
rect 195388 245024 196716 245052
rect 195388 245012 195394 245024
rect 196710 245012 196716 245024
rect 196768 245012 196774 245064
rect 137462 244876 137468 244928
rect 137520 244916 137526 244928
rect 189810 244916 189816 244928
rect 137520 244888 189816 244916
rect 137520 244876 137526 244888
rect 189810 244876 189816 244888
rect 189868 244876 189874 244928
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 123754 244304 123760 244316
rect 121604 244276 123760 244304
rect 121604 244264 121610 244276
rect 123754 244264 123760 244276
rect 123812 244264 123818 244316
rect 321738 244264 321744 244316
rect 321796 244304 321802 244316
rect 378778 244304 378784 244316
rect 321796 244276 378784 244304
rect 321796 244264 321802 244276
rect 378778 244264 378784 244276
rect 378836 244264 378842 244316
rect 37090 244196 37096 244248
rect 37148 244236 37154 244248
rect 67726 244236 67732 244248
rect 37148 244208 67732 244236
rect 37148 244196 37154 244208
rect 67726 244196 67732 244208
rect 67784 244196 67790 244248
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 131206 244236 131212 244248
rect 121512 244208 131212 244236
rect 121512 244196 121518 244208
rect 131206 244196 131212 244208
rect 131264 244196 131270 244248
rect 49510 244128 49516 244180
rect 49568 244168 49574 244180
rect 67634 244168 67640 244180
rect 49568 244140 67640 244168
rect 49568 244128 49574 244140
rect 67634 244128 67640 244140
rect 67692 244128 67698 244180
rect 194226 243788 194232 243840
rect 194284 243828 194290 243840
rect 195974 243828 195980 243840
rect 194284 243800 195980 243828
rect 194284 243788 194290 243800
rect 195974 243788 195980 243800
rect 196032 243828 196038 243840
rect 198274 243828 198280 243840
rect 196032 243800 198280 243828
rect 196032 243788 196038 243800
rect 198274 243788 198280 243800
rect 198332 243788 198338 243840
rect 194318 243652 194324 243704
rect 194376 243692 194382 243704
rect 195974 243692 195980 243704
rect 194376 243664 195980 243692
rect 194376 243652 194382 243664
rect 195974 243652 195980 243664
rect 196032 243652 196038 243704
rect 68554 243516 68560 243568
rect 68612 243556 68618 243568
rect 68922 243556 68928 243568
rect 68612 243528 68928 243556
rect 68612 243516 68618 243528
rect 68922 243516 68928 243528
rect 68980 243516 68986 243568
rect 145650 243516 145656 243568
rect 145708 243556 145714 243568
rect 195330 243556 195336 243568
rect 145708 243528 195336 243556
rect 145708 243516 145714 243528
rect 195330 243516 195336 243528
rect 195388 243516 195394 243568
rect 135162 242972 135168 243024
rect 135220 243012 135226 243024
rect 176102 243012 176108 243024
rect 135220 242984 176108 243012
rect 135220 242972 135226 242984
rect 176102 242972 176108 242984
rect 176160 242972 176166 243024
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 191650 242944 191656 242956
rect 121604 242916 191656 242944
rect 121604 242904 121610 242916
rect 191650 242904 191656 242916
rect 191708 242904 191714 242956
rect 321462 242904 321468 242956
rect 321520 242944 321526 242956
rect 443638 242944 443644 242956
rect 321520 242916 443644 242944
rect 321520 242904 321526 242916
rect 443638 242904 443644 242916
rect 443696 242904 443702 242956
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 134610 242876 134616 242888
rect 121512 242848 134616 242876
rect 121512 242836 121518 242848
rect 134610 242836 134616 242848
rect 134668 242876 134674 242888
rect 135162 242876 135168 242888
rect 134668 242848 135168 242876
rect 134668 242836 134674 242848
rect 135162 242836 135168 242848
rect 135220 242836 135226 242888
rect 155494 242156 155500 242208
rect 155552 242196 155558 242208
rect 193858 242196 193864 242208
rect 155552 242168 193864 242196
rect 155552 242156 155558 242168
rect 193858 242156 193864 242168
rect 193916 242156 193922 242208
rect 121454 241476 121460 241528
rect 121512 241516 121518 241528
rect 140682 241516 140688 241528
rect 121512 241488 140688 241516
rect 121512 241476 121518 241488
rect 140682 241476 140688 241488
rect 140740 241476 140746 241528
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 40862 241448 40868 241460
rect 3476 241420 40868 241448
rect 3476 241408 3482 241420
rect 40862 241408 40868 241420
rect 40920 241448 40926 241460
rect 41230 241448 41236 241460
rect 40920 241420 41236 241448
rect 40920 241408 40926 241420
rect 41230 241408 41236 241420
rect 41288 241408 41294 241460
rect 322198 241408 322204 241460
rect 322256 241448 322262 241460
rect 324590 241448 324596 241460
rect 322256 241420 324596 241448
rect 322256 241408 322262 241420
rect 324590 241408 324596 241420
rect 324648 241408 324654 241460
rect 162394 240796 162400 240848
rect 162452 240836 162458 240848
rect 195790 240836 195796 240848
rect 162452 240808 195796 240836
rect 162452 240796 162458 240808
rect 195790 240796 195796 240808
rect 195848 240796 195854 240848
rect 40862 240728 40868 240780
rect 40920 240768 40926 240780
rect 58710 240768 58716 240780
rect 40920 240740 58716 240768
rect 40920 240728 40926 240740
rect 58710 240728 58716 240740
rect 58768 240728 58774 240780
rect 144454 240728 144460 240780
rect 144512 240768 144518 240780
rect 196526 240768 196532 240780
rect 144512 240740 196532 240768
rect 144512 240728 144518 240740
rect 196526 240728 196532 240740
rect 196584 240728 196590 240780
rect 121454 240252 121460 240304
rect 121512 240292 121518 240304
rect 155494 240292 155500 240304
rect 121512 240264 155500 240292
rect 121512 240252 121518 240264
rect 155494 240252 155500 240264
rect 155552 240252 155558 240304
rect 120626 240184 120632 240236
rect 120684 240224 120690 240236
rect 191190 240224 191196 240236
rect 120684 240196 191196 240224
rect 120684 240184 120690 240196
rect 191190 240184 191196 240196
rect 191248 240184 191254 240236
rect 119982 240116 119988 240168
rect 120040 240156 120046 240168
rect 199654 240156 199660 240168
rect 120040 240128 199660 240156
rect 120040 240116 120046 240128
rect 199654 240116 199660 240128
rect 199712 240116 199718 240168
rect 324590 240116 324596 240168
rect 324648 240156 324654 240168
rect 502334 240156 502340 240168
rect 324648 240128 502340 240156
rect 324648 240116 324654 240128
rect 502334 240116 502340 240128
rect 502392 240116 502398 240168
rect 3510 240048 3516 240100
rect 3568 240088 3574 240100
rect 37182 240088 37188 240100
rect 3568 240060 37188 240088
rect 3568 240048 3574 240060
rect 37182 240048 37188 240060
rect 37240 240048 37246 240100
rect 194502 240048 194508 240100
rect 194560 240088 194566 240100
rect 196802 240088 196808 240100
rect 194560 240060 196808 240088
rect 194560 240048 194566 240060
rect 196802 240048 196808 240060
rect 196860 240048 196866 240100
rect 70394 239776 70400 239828
rect 70452 239816 70458 239828
rect 71302 239816 71308 239828
rect 70452 239788 71308 239816
rect 70452 239776 70458 239788
rect 71302 239776 71308 239788
rect 71360 239776 71366 239828
rect 76006 239776 76012 239828
rect 76064 239816 76070 239828
rect 77098 239816 77104 239828
rect 76064 239788 77104 239816
rect 76064 239776 76070 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 84286 239776 84292 239828
rect 84344 239816 84350 239828
rect 85470 239816 85476 239828
rect 84344 239788 85476 239816
rect 84344 239776 84350 239788
rect 85470 239776 85476 239788
rect 85528 239776 85534 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 89714 239776 89720 239828
rect 89772 239816 89778 239828
rect 90622 239816 90628 239828
rect 89772 239788 90628 239816
rect 89772 239776 89778 239788
rect 90622 239776 90628 239788
rect 90680 239776 90686 239828
rect 95234 239776 95240 239828
rect 95292 239816 95298 239828
rect 96418 239816 96424 239828
rect 95292 239788 96424 239816
rect 95292 239776 95298 239788
rect 96418 239776 96424 239788
rect 96476 239776 96482 239828
rect 102134 239776 102140 239828
rect 102192 239816 102198 239828
rect 102858 239816 102864 239828
rect 102192 239788 102864 239816
rect 102192 239776 102198 239788
rect 102858 239776 102864 239788
rect 102916 239776 102922 239828
rect 107654 239776 107660 239828
rect 107712 239816 107718 239828
rect 108654 239816 108660 239828
rect 107712 239788 108660 239816
rect 107712 239776 107718 239788
rect 108654 239776 108660 239788
rect 108712 239776 108718 239828
rect 110414 239776 110420 239828
rect 110472 239816 110478 239828
rect 111230 239816 111236 239828
rect 110472 239788 111236 239816
rect 110472 239776 110478 239788
rect 111230 239776 111236 239788
rect 111288 239776 111294 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 219434 239776 219440 239828
rect 219492 239816 219498 239828
rect 220584 239816 220590 239828
rect 219492 239788 220590 239816
rect 219492 239776 219498 239788
rect 220584 239776 220590 239788
rect 220642 239776 220648 239828
rect 238754 239776 238760 239828
rect 238812 239816 238818 239828
rect 239904 239816 239910 239828
rect 238812 239788 239910 239816
rect 238812 239776 238818 239788
rect 239904 239776 239910 239788
rect 239962 239776 239968 239828
rect 247034 239776 247040 239828
rect 247092 239816 247098 239828
rect 248276 239816 248282 239828
rect 247092 239788 248282 239816
rect 247092 239776 247098 239788
rect 248276 239776 248282 239788
rect 248334 239776 248340 239828
rect 258074 239776 258080 239828
rect 258132 239816 258138 239828
rect 259224 239816 259230 239828
rect 258132 239788 259230 239816
rect 258132 239776 258138 239788
rect 259224 239776 259230 239788
rect 259282 239776 259288 239828
rect 266354 239776 266360 239828
rect 266412 239816 266418 239828
rect 267596 239816 267602 239828
rect 266412 239788 267602 239816
rect 266412 239776 266418 239788
rect 267596 239776 267602 239788
rect 267654 239776 267660 239828
rect 285674 239776 285680 239828
rect 285732 239816 285738 239828
rect 286916 239816 286922 239828
rect 285732 239788 286922 239816
rect 285732 239776 285738 239788
rect 286916 239776 286922 239788
rect 286974 239776 286980 239828
rect 63126 239572 63132 239624
rect 63184 239612 63190 239624
rect 73798 239612 73804 239624
rect 63184 239584 73804 239612
rect 63184 239572 63190 239584
rect 73798 239572 73804 239584
rect 73856 239572 73862 239624
rect 60366 239504 60372 239556
rect 60424 239544 60430 239556
rect 76374 239544 76380 239556
rect 60424 239516 76380 239544
rect 60424 239504 60430 239516
rect 76374 239504 76380 239516
rect 76432 239504 76438 239556
rect 65978 239436 65984 239488
rect 66036 239476 66042 239488
rect 195054 239476 195060 239488
rect 66036 239448 195060 239476
rect 66036 239436 66042 239448
rect 195054 239436 195060 239448
rect 195112 239436 195118 239488
rect 204162 239436 204168 239488
rect 204220 239476 204226 239488
rect 319530 239476 319536 239488
rect 204220 239448 319536 239476
rect 204220 239436 204226 239448
rect 319530 239436 319536 239448
rect 319588 239436 319594 239488
rect 69842 239368 69848 239420
rect 69900 239408 69906 239420
rect 83458 239408 83464 239420
rect 69900 239380 83464 239408
rect 69900 239368 69906 239380
rect 83458 239368 83464 239380
rect 83516 239368 83522 239420
rect 191650 239368 191656 239420
rect 191708 239408 191714 239420
rect 320082 239408 320088 239420
rect 191708 239380 320088 239408
rect 191708 239368 191714 239380
rect 320082 239368 320088 239380
rect 320140 239408 320146 239420
rect 321738 239408 321744 239420
rect 320140 239380 321744 239408
rect 320140 239368 320146 239380
rect 321738 239368 321744 239380
rect 321796 239368 321802 239420
rect 535454 239368 535460 239420
rect 535512 239408 535518 239420
rect 580166 239408 580172 239420
rect 535512 239380 580172 239408
rect 535512 239368 535518 239380
rect 580166 239368 580172 239380
rect 580224 239368 580230 239420
rect 200942 239164 200948 239216
rect 201000 239204 201006 239216
rect 204898 239204 204904 239216
rect 201000 239176 204904 239204
rect 201000 239164 201006 239176
rect 204898 239164 204904 239176
rect 204956 239164 204962 239216
rect 199838 239096 199844 239148
rect 199896 239136 199902 239148
rect 202230 239136 202236 239148
rect 199896 239108 202236 239136
rect 199896 239096 199902 239108
rect 202230 239096 202236 239108
rect 202288 239096 202294 239148
rect 77754 239028 77760 239080
rect 77812 239068 77818 239080
rect 200114 239068 200120 239080
rect 77812 239040 200120 239068
rect 77812 239028 77818 239040
rect 200114 239028 200120 239040
rect 200172 239028 200178 239080
rect 104158 238960 104164 239012
rect 104216 239000 104222 239012
rect 120810 239000 120816 239012
rect 104216 238972 120816 239000
rect 104216 238960 104222 238972
rect 120810 238960 120816 238972
rect 120868 238960 120874 239012
rect 121454 238960 121460 239012
rect 121512 239000 121518 239012
rect 155586 239000 155592 239012
rect 121512 238972 155592 239000
rect 121512 238960 121518 238972
rect 155586 238960 155592 238972
rect 155644 238960 155650 239012
rect 195974 238960 195980 239012
rect 196032 239000 196038 239012
rect 202138 239000 202144 239012
rect 196032 238972 202144 239000
rect 196032 238960 196038 238972
rect 202138 238960 202144 238972
rect 202196 238960 202202 239012
rect 85574 238892 85580 238944
rect 85632 238932 85638 238944
rect 86770 238932 86776 238944
rect 85632 238904 86776 238932
rect 85632 238892 85638 238904
rect 86770 238892 86776 238904
rect 86828 238932 86834 238944
rect 123570 238932 123576 238944
rect 86828 238904 123576 238932
rect 86828 238892 86834 238904
rect 123570 238892 123576 238904
rect 123628 238892 123634 238944
rect 37182 238824 37188 238876
rect 37240 238864 37246 238876
rect 111886 238864 111892 238876
rect 37240 238836 111892 238864
rect 37240 238824 37246 238836
rect 111886 238824 111892 238836
rect 111944 238864 111950 238876
rect 112530 238864 112536 238876
rect 111944 238836 112536 238864
rect 111944 238824 111950 238836
rect 112530 238824 112536 238836
rect 112588 238824 112594 238876
rect 114462 238824 114468 238876
rect 114520 238864 114526 238876
rect 124398 238864 124404 238876
rect 114520 238836 124404 238864
rect 114520 238824 114526 238836
rect 124398 238824 124404 238836
rect 124456 238824 124462 238876
rect 152734 238824 152740 238876
rect 152792 238864 152798 238876
rect 237374 238864 237380 238876
rect 152792 238836 237380 238864
rect 152792 238824 152798 238836
rect 237374 238824 237380 238836
rect 237432 238864 237438 238876
rect 238018 238864 238024 238876
rect 237432 238836 238024 238864
rect 237432 238824 237438 238836
rect 238018 238824 238024 238836
rect 238076 238824 238082 238876
rect 201586 238756 201592 238808
rect 201644 238796 201650 238808
rect 252830 238796 252836 238808
rect 201644 238768 252836 238796
rect 201644 238756 201650 238768
rect 252830 238756 252836 238768
rect 252888 238796 252894 238808
rect 535454 238796 535460 238808
rect 252888 238768 535460 238796
rect 252888 238756 252894 238768
rect 535454 238756 535460 238768
rect 535512 238756 535518 238808
rect 50982 238688 50988 238740
rect 51040 238728 51046 238740
rect 82262 238728 82268 238740
rect 51040 238700 82268 238728
rect 51040 238688 51046 238700
rect 82262 238688 82268 238700
rect 82320 238688 82326 238740
rect 118970 238688 118976 238740
rect 119028 238728 119034 238740
rect 130562 238728 130568 238740
rect 119028 238700 130568 238728
rect 119028 238688 119034 238700
rect 130562 238688 130568 238700
rect 130620 238688 130626 238740
rect 48130 238620 48136 238672
rect 48188 238660 48194 238672
rect 72602 238660 72608 238672
rect 48188 238632 72608 238660
rect 48188 238620 48194 238632
rect 72602 238620 72608 238632
rect 72660 238620 72666 238672
rect 83550 238620 83556 238672
rect 83608 238660 83614 238672
rect 149054 238660 149060 238672
rect 83608 238632 149060 238660
rect 83608 238620 83614 238632
rect 149054 238620 149060 238632
rect 149112 238660 149118 238672
rect 316586 238660 316592 238672
rect 149112 238632 316592 238660
rect 149112 238620 149118 238632
rect 316586 238620 316592 238632
rect 316644 238620 316650 238672
rect 88702 238552 88708 238604
rect 88760 238592 88766 238604
rect 241882 238592 241888 238604
rect 88760 238564 241888 238592
rect 88760 238552 88766 238564
rect 241882 238552 241888 238564
rect 241940 238552 241946 238604
rect 118326 238484 118332 238536
rect 118384 238524 118390 238536
rect 144914 238524 144920 238536
rect 118384 238496 144920 238524
rect 118384 238484 118390 238496
rect 144914 238484 144920 238496
rect 144972 238484 144978 238536
rect 195330 238484 195336 238536
rect 195388 238524 195394 238536
rect 331582 238524 331588 238536
rect 195388 238496 331588 238524
rect 195388 238484 195394 238496
rect 331582 238484 331588 238496
rect 331640 238484 331646 238536
rect 115106 238416 115112 238468
rect 115164 238456 115170 238468
rect 146294 238456 146300 238468
rect 115164 238428 146300 238456
rect 115164 238416 115170 238428
rect 146294 238416 146300 238428
rect 146352 238416 146358 238468
rect 200114 238416 200120 238468
rect 200172 238456 200178 238468
rect 216766 238456 216772 238468
rect 200172 238428 216772 238456
rect 200172 238416 200178 238428
rect 216766 238416 216772 238428
rect 216824 238416 216830 238468
rect 105446 238348 105452 238400
rect 105504 238388 105510 238400
rect 282178 238388 282184 238400
rect 105504 238360 282184 238388
rect 105504 238348 105510 238360
rect 282178 238348 282184 238360
rect 282236 238348 282242 238400
rect 69934 238280 69940 238332
rect 69992 238320 69998 238332
rect 119982 238320 119988 238332
rect 69992 238292 119988 238320
rect 69992 238280 69998 238292
rect 119982 238280 119988 238292
rect 120040 238280 120046 238332
rect 71958 238144 71964 238196
rect 72016 238184 72022 238196
rect 79226 238184 79232 238196
rect 72016 238156 79232 238184
rect 72016 238144 72022 238156
rect 79226 238144 79232 238156
rect 79284 238144 79290 238196
rect 80974 238144 80980 238196
rect 81032 238184 81038 238196
rect 88978 238184 88984 238196
rect 81032 238156 88984 238184
rect 81032 238144 81038 238156
rect 88978 238144 88984 238156
rect 89036 238144 89042 238196
rect 73246 238076 73252 238128
rect 73304 238116 73310 238128
rect 86218 238116 86224 238128
rect 73304 238088 86224 238116
rect 73304 238076 73310 238088
rect 86218 238076 86224 238088
rect 86276 238076 86282 238128
rect 196618 238076 196624 238128
rect 196676 238116 196682 238128
rect 204070 238116 204076 238128
rect 196676 238088 204076 238116
rect 196676 238076 196682 238088
rect 204070 238076 204076 238088
rect 204128 238076 204134 238128
rect 315942 238076 315948 238128
rect 316000 238116 316006 238128
rect 320174 238116 320180 238128
rect 316000 238088 320180 238116
rect 316000 238076 316006 238088
rect 320174 238076 320180 238088
rect 320232 238076 320238 238128
rect 67542 238008 67548 238060
rect 67600 238048 67606 238060
rect 105538 238048 105544 238060
rect 67600 238020 105544 238048
rect 67600 238008 67606 238020
rect 105538 238008 105544 238020
rect 105596 238008 105602 238060
rect 184290 238008 184296 238060
rect 184348 238048 184354 238060
rect 200666 238048 200672 238060
rect 184348 238020 200672 238048
rect 184348 238008 184354 238020
rect 200666 238008 200672 238020
rect 200724 238008 200730 238060
rect 316586 238008 316592 238060
rect 316644 238048 316650 238060
rect 438854 238048 438860 238060
rect 316644 238020 438860 238048
rect 316644 238008 316650 238020
rect 438854 238008 438860 238020
rect 438912 238008 438918 238060
rect 204070 237668 204076 237720
rect 204128 237708 204134 237720
rect 205818 237708 205824 237720
rect 204128 237680 205824 237708
rect 204128 237668 204134 237680
rect 205818 237668 205824 237680
rect 205876 237668 205882 237720
rect 244274 237464 244280 237516
rect 244332 237504 244338 237516
rect 246390 237504 246396 237516
rect 244332 237476 246396 237504
rect 244332 237464 244338 237476
rect 246390 237464 246396 237476
rect 246448 237464 246454 237516
rect 216766 237396 216772 237448
rect 216824 237436 216830 237448
rect 217318 237436 217324 237448
rect 216824 237408 217324 237436
rect 216824 237396 216830 237408
rect 217318 237396 217324 237408
rect 217376 237396 217382 237448
rect 221458 237396 221464 237448
rect 221516 237436 221522 237448
rect 223206 237436 223212 237448
rect 221516 237408 223212 237436
rect 221516 237396 221522 237408
rect 223206 237396 223212 237408
rect 223264 237396 223270 237448
rect 229738 237396 229744 237448
rect 229796 237436 229802 237448
rect 231578 237436 231584 237448
rect 229796 237408 231584 237436
rect 229796 237396 229802 237408
rect 231578 237396 231584 237408
rect 231636 237396 231642 237448
rect 235350 237396 235356 237448
rect 235408 237436 235414 237448
rect 236086 237436 236092 237448
rect 235408 237408 236092 237436
rect 235408 237396 235414 237408
rect 236086 237396 236092 237408
rect 236144 237396 236150 237448
rect 246298 237396 246304 237448
rect 246356 237436 246362 237448
rect 250898 237436 250904 237448
rect 246356 237408 250904 237436
rect 246356 237396 246362 237408
rect 250898 237396 250904 237408
rect 250956 237396 250962 237448
rect 251818 237396 251824 237448
rect 251876 237436 251882 237448
rect 254762 237436 254768 237448
rect 251876 237408 254768 237436
rect 251876 237396 251882 237408
rect 254762 237396 254768 237408
rect 254820 237396 254826 237448
rect 291838 237396 291844 237448
rect 291896 237436 291902 237448
rect 297266 237436 297272 237448
rect 291896 237408 297272 237436
rect 291896 237396 291902 237408
rect 297266 237396 297272 237408
rect 297324 237396 297330 237448
rect 300118 237396 300124 237448
rect 300176 237436 300182 237448
rect 301774 237436 301780 237448
rect 300176 237408 301780 237436
rect 300176 237396 300182 237408
rect 301774 237396 301780 237408
rect 301832 237396 301838 237448
rect 307110 237396 307116 237448
rect 307168 237436 307174 237448
rect 308214 237436 308220 237448
rect 307168 237408 308220 237436
rect 307168 237396 307174 237408
rect 308214 237396 308220 237408
rect 308272 237396 308278 237448
rect 312630 237396 312636 237448
rect 312688 237436 312694 237448
rect 314010 237436 314016 237448
rect 312688 237408 314016 237436
rect 312688 237396 312694 237408
rect 314010 237396 314016 237408
rect 314068 237396 314074 237448
rect 318058 237396 318064 237448
rect 318116 237436 318122 237448
rect 318518 237436 318524 237448
rect 318116 237408 318524 237436
rect 318116 237396 318122 237408
rect 318518 237396 318524 237408
rect 318576 237436 318582 237448
rect 498286 237436 498292 237448
rect 318576 237408 498292 237436
rect 318576 237396 318582 237408
rect 498286 237396 498292 237408
rect 498344 237396 498350 237448
rect 58710 237328 58716 237380
rect 58768 237368 58774 237380
rect 103514 237368 103520 237380
rect 58768 237340 103520 237368
rect 58768 237328 58774 237340
rect 103514 237328 103520 237340
rect 103572 237328 103578 237380
rect 113174 237328 113180 237380
rect 113232 237368 113238 237380
rect 114462 237368 114468 237380
rect 113232 237340 114468 237368
rect 113232 237328 113238 237340
rect 114462 237328 114468 237340
rect 114520 237368 114526 237380
rect 149790 237368 149796 237380
rect 114520 237340 149796 237368
rect 114520 237328 114526 237340
rect 149790 237328 149796 237340
rect 149848 237328 149854 237380
rect 197998 237328 198004 237380
rect 198056 237368 198062 237380
rect 204162 237368 204168 237380
rect 198056 237340 204168 237368
rect 198056 237328 198062 237340
rect 204162 237328 204168 237340
rect 204220 237328 204226 237380
rect 55122 237260 55128 237312
rect 55180 237300 55186 237312
rect 86126 237300 86132 237312
rect 55180 237272 86132 237300
rect 55180 237260 55186 237272
rect 86126 237260 86132 237272
rect 86184 237260 86190 237312
rect 95786 237260 95792 237312
rect 95844 237300 95850 237312
rect 126974 237300 126980 237312
rect 95844 237272 126980 237300
rect 95844 237260 95850 237272
rect 126974 237260 126980 237272
rect 127032 237260 127038 237312
rect 142890 237260 142896 237312
rect 142948 237300 142954 237312
rect 331306 237300 331312 237312
rect 142948 237272 331312 237300
rect 142948 237260 142954 237272
rect 331306 237260 331312 237272
rect 331364 237260 331370 237312
rect 49602 237192 49608 237244
rect 49660 237232 49666 237244
rect 76650 237232 76656 237244
rect 49660 237204 76656 237232
rect 49660 237192 49666 237204
rect 76650 237192 76656 237204
rect 76708 237192 76714 237244
rect 113818 237192 113824 237244
rect 113876 237232 113882 237244
rect 133874 237232 133880 237244
rect 113876 237204 133880 237232
rect 113876 237192 113882 237204
rect 133874 237192 133880 237204
rect 133932 237192 133938 237244
rect 151354 237192 151360 237244
rect 151412 237232 151418 237244
rect 328546 237232 328552 237244
rect 151412 237204 328552 237232
rect 151412 237192 151418 237204
rect 328546 237192 328552 237204
rect 328604 237192 328610 237244
rect 195882 237124 195888 237176
rect 195940 237164 195946 237176
rect 303706 237164 303712 237176
rect 195940 237136 303712 237164
rect 195940 237124 195946 237136
rect 303706 237124 303712 237136
rect 303764 237124 303770 237176
rect 148594 237056 148600 237108
rect 148652 237096 148658 237108
rect 195974 237096 195980 237108
rect 148652 237068 195980 237096
rect 148652 237056 148658 237068
rect 195974 237056 195980 237068
rect 196032 237056 196038 237108
rect 183370 236988 183376 237040
rect 183428 237028 183434 237040
rect 504358 237028 504364 237040
rect 183428 237000 504364 237028
rect 183428 236988 183434 237000
rect 504358 236988 504364 237000
rect 504416 236988 504422 237040
rect 160922 236716 160928 236768
rect 160980 236756 160986 236768
rect 195330 236756 195336 236768
rect 160980 236728 195336 236756
rect 160980 236716 160986 236728
rect 195330 236716 195336 236728
rect 195388 236716 195394 236768
rect 68646 236648 68652 236700
rect 68704 236688 68710 236700
rect 249794 236688 249800 236700
rect 68704 236660 249800 236688
rect 68704 236648 68710 236660
rect 249794 236648 249800 236660
rect 249852 236648 249858 236700
rect 316678 235968 316684 236020
rect 316736 236008 316742 236020
rect 320266 236008 320272 236020
rect 316736 235980 320272 236008
rect 316736 235968 316742 235980
rect 320266 235968 320272 235980
rect 320324 235968 320330 236020
rect 503714 235968 503720 236020
rect 503772 236008 503778 236020
rect 504358 236008 504364 236020
rect 503772 235980 504364 236008
rect 503772 235968 503778 235980
rect 504358 235968 504364 235980
rect 504416 235968 504422 236020
rect 89346 235900 89352 235952
rect 89404 235940 89410 235952
rect 142154 235940 142160 235952
rect 89404 235912 142160 235940
rect 89404 235900 89410 235912
rect 142154 235900 142160 235912
rect 142212 235900 142218 235952
rect 158162 235900 158168 235952
rect 158220 235940 158226 235952
rect 329926 235940 329932 235952
rect 158220 235912 329932 235940
rect 158220 235900 158226 235912
rect 329926 235900 329932 235912
rect 329984 235900 329990 235952
rect 91278 235832 91284 235884
rect 91336 235872 91342 235884
rect 129274 235872 129280 235884
rect 91336 235844 129280 235872
rect 91336 235832 91342 235844
rect 129274 235832 129280 235844
rect 129332 235832 129338 235884
rect 174630 235832 174636 235884
rect 174688 235872 174694 235884
rect 244274 235872 244280 235884
rect 174688 235844 244280 235872
rect 174688 235832 174694 235844
rect 244274 235832 244280 235844
rect 244332 235872 244338 235884
rect 244918 235872 244924 235884
rect 244332 235844 244924 235872
rect 244332 235832 244338 235844
rect 244918 235832 244924 235844
rect 244976 235832 244982 235884
rect 73890 235764 73896 235816
rect 73948 235804 73954 235816
rect 120626 235804 120632 235816
rect 73948 235776 120632 235804
rect 73948 235764 73954 235776
rect 120626 235764 120632 235776
rect 120684 235764 120690 235816
rect 39758 235696 39764 235748
rect 39816 235736 39822 235748
rect 91738 235736 91744 235748
rect 39816 235708 91744 235736
rect 39816 235696 39822 235708
rect 91738 235696 91744 235708
rect 91796 235696 91802 235748
rect 118602 235696 118608 235748
rect 118660 235736 118666 235748
rect 131114 235736 131120 235748
rect 118660 235708 131120 235736
rect 118660 235696 118666 235708
rect 131114 235696 131120 235708
rect 131172 235696 131178 235748
rect 194226 235492 194232 235544
rect 194284 235532 194290 235544
rect 213178 235532 213184 235544
rect 194284 235504 213184 235532
rect 194284 235492 194290 235504
rect 213178 235492 213184 235504
rect 213236 235492 213242 235544
rect 163590 235424 163596 235476
rect 163648 235464 163654 235476
rect 196618 235464 196624 235476
rect 163648 235436 196624 235464
rect 163648 235424 163654 235436
rect 196618 235424 196624 235436
rect 196676 235424 196682 235476
rect 187050 235356 187056 235408
rect 187108 235396 187114 235408
rect 222838 235396 222844 235408
rect 187108 235368 222844 235396
rect 187108 235356 187114 235368
rect 222838 235356 222844 235368
rect 222896 235356 222902 235408
rect 106090 235288 106096 235340
rect 106148 235328 106154 235340
rect 175090 235328 175096 235340
rect 106148 235300 175096 235328
rect 106148 235288 106154 235300
rect 175090 235288 175096 235300
rect 175148 235288 175154 235340
rect 198826 235288 198832 235340
rect 198884 235328 198890 235340
rect 324682 235328 324688 235340
rect 198884 235300 324688 235328
rect 198884 235288 198890 235300
rect 324682 235288 324688 235300
rect 324740 235288 324746 235340
rect 67358 235220 67364 235272
rect 67416 235260 67422 235272
rect 280246 235260 280252 235272
rect 67416 235232 280252 235260
rect 67416 235220 67422 235232
rect 280246 235220 280252 235232
rect 280304 235220 280310 235272
rect 303706 235220 303712 235272
rect 303764 235260 303770 235272
rect 498378 235260 498384 235272
rect 303764 235232 498384 235260
rect 303764 235220 303770 235232
rect 498378 235220 498384 235232
rect 498436 235220 498442 235272
rect 175090 235084 175096 235136
rect 175148 235124 175154 235136
rect 176010 235124 176016 235136
rect 175148 235096 176016 235124
rect 175148 235084 175154 235096
rect 176010 235084 176016 235096
rect 176068 235084 176074 235136
rect 117682 234948 117688 235000
rect 117740 234988 117746 235000
rect 118602 234988 118608 235000
rect 117740 234960 118608 234988
rect 117740 234948 117746 234960
rect 118602 234948 118608 234960
rect 118660 234948 118666 235000
rect 288894 234608 288900 234660
rect 288952 234648 288958 234660
rect 289446 234648 289452 234660
rect 288952 234620 289452 234648
rect 288952 234608 288958 234620
rect 289446 234608 289452 234620
rect 289504 234648 289510 234660
rect 432598 234648 432604 234660
rect 289504 234620 432604 234648
rect 289504 234608 289510 234620
rect 432598 234608 432604 234620
rect 432656 234608 432662 234660
rect 46566 234540 46572 234592
rect 46624 234580 46630 234592
rect 109034 234580 109040 234592
rect 46624 234552 109040 234580
rect 46624 234540 46630 234552
rect 109034 234540 109040 234552
rect 109092 234540 109098 234592
rect 134702 234540 134708 234592
rect 134760 234580 134766 234592
rect 327258 234580 327264 234592
rect 134760 234552 327264 234580
rect 134760 234540 134766 234552
rect 327258 234540 327264 234552
rect 327316 234580 327322 234592
rect 328362 234580 328368 234592
rect 327316 234552 328368 234580
rect 327316 234540 327322 234552
rect 328362 234540 328368 234552
rect 328420 234540 328426 234592
rect 48222 234472 48228 234524
rect 48280 234512 48286 234524
rect 195146 234512 195152 234524
rect 48280 234484 195152 234512
rect 48280 234472 48286 234484
rect 195146 234472 195152 234484
rect 195204 234472 195210 234524
rect 196526 234472 196532 234524
rect 196584 234512 196590 234524
rect 321462 234512 321468 234524
rect 196584 234484 321468 234512
rect 196584 234472 196590 234484
rect 321462 234472 321468 234484
rect 321520 234512 321526 234524
rect 322198 234512 322204 234524
rect 321520 234484 322204 234512
rect 321520 234472 321526 234484
rect 322198 234472 322204 234484
rect 322256 234472 322262 234524
rect 50338 234404 50344 234456
rect 50396 234444 50402 234456
rect 85574 234444 85580 234456
rect 50396 234416 85580 234444
rect 50396 234404 50402 234416
rect 85574 234404 85580 234416
rect 85632 234404 85638 234456
rect 200666 234404 200672 234456
rect 200724 234444 200730 234456
rect 321554 234444 321560 234456
rect 200724 234416 321560 234444
rect 200724 234404 200730 234416
rect 321554 234404 321560 234416
rect 321612 234444 321618 234456
rect 321830 234444 321836 234456
rect 321612 234416 321836 234444
rect 321612 234404 321618 234416
rect 321830 234404 321836 234416
rect 321888 234404 321894 234456
rect 159634 234336 159640 234388
rect 159692 234376 159698 234388
rect 218698 234376 218704 234388
rect 159692 234348 218704 234376
rect 159692 234336 159698 234348
rect 218698 234336 218704 234348
rect 218756 234336 218762 234388
rect 109034 234132 109040 234184
rect 109092 234172 109098 234184
rect 109954 234172 109960 234184
rect 109092 234144 109960 234172
rect 109092 234132 109098 234144
rect 109954 234132 109960 234144
rect 110012 234132 110018 234184
rect 47578 234064 47584 234116
rect 47636 234104 47642 234116
rect 48222 234104 48228 234116
rect 47636 234076 48228 234104
rect 47636 234064 47642 234076
rect 48222 234064 48228 234076
rect 48280 234064 48286 234116
rect 84166 234008 93854 234036
rect 74534 233860 74540 233912
rect 74592 233900 74598 233912
rect 75178 233900 75184 233912
rect 74592 233872 75184 233900
rect 74592 233860 74598 233872
rect 75178 233860 75184 233872
rect 75236 233860 75242 233912
rect 79226 233860 79232 233912
rect 79284 233900 79290 233912
rect 84166 233900 84194 234008
rect 84286 233928 84292 233980
rect 84344 233928 84350 233980
rect 79284 233872 84194 233900
rect 79284 233860 79290 233872
rect 84194 233724 84200 233776
rect 84252 233764 84258 233776
rect 84304 233764 84332 233928
rect 93826 233900 93854 234008
rect 171870 233928 171876 233980
rect 171928 233968 171934 233980
rect 270494 233968 270500 233980
rect 171928 233940 270500 233968
rect 171928 233928 171934 233940
rect 270494 233928 270500 233940
rect 270552 233928 270558 233980
rect 328362 233928 328368 233980
rect 328420 233968 328426 233980
rect 335354 233968 335360 233980
rect 328420 233940 335360 233968
rect 328420 233928 328426 233940
rect 335354 233928 335360 233940
rect 335412 233928 335418 233980
rect 202782 233900 202788 233912
rect 93826 233872 202788 233900
rect 202782 233860 202788 233872
rect 202840 233900 202846 233912
rect 203886 233900 203892 233912
rect 202840 233872 203892 233900
rect 202840 233860 202846 233872
rect 203886 233860 203892 233872
rect 203944 233860 203950 233912
rect 321554 233860 321560 233912
rect 321612 233900 321618 233912
rect 333974 233900 333980 233912
rect 321612 233872 333980 233900
rect 321612 233860 321618 233872
rect 333974 233860 333980 233872
rect 334032 233860 334038 233912
rect 84252 233736 84332 233764
rect 84252 233724 84258 233736
rect 60458 233180 60464 233232
rect 60516 233220 60522 233232
rect 327074 233220 327080 233232
rect 60516 233192 327080 233220
rect 60516 233180 60522 233192
rect 327074 233180 327080 233192
rect 327132 233220 327138 233232
rect 328362 233220 328368 233232
rect 327132 233192 328368 233220
rect 327132 233180 327138 233192
rect 328362 233180 328368 233192
rect 328420 233180 328426 233232
rect 56502 233112 56508 233164
rect 56560 233152 56566 233164
rect 178862 233152 178868 233164
rect 56560 233124 178868 233152
rect 56560 233112 56566 233124
rect 178862 233112 178868 233124
rect 178920 233112 178926 233164
rect 81618 233044 81624 233096
rect 81676 233084 81682 233096
rect 132586 233084 132592 233096
rect 81676 233056 132592 233084
rect 81676 233044 81682 233056
rect 132586 233044 132592 233056
rect 132644 233044 132650 233096
rect 156782 233044 156788 233096
rect 156840 233084 156846 233096
rect 265618 233084 265624 233096
rect 156840 233056 265624 233084
rect 156840 233044 156846 233056
rect 265618 233044 265624 233056
rect 265676 233044 265682 233096
rect 166534 232976 166540 233028
rect 166592 233016 166598 233028
rect 262950 233016 262956 233028
rect 166592 232988 262956 233016
rect 166592 232976 166598 232988
rect 262950 232976 262956 232988
rect 263008 232976 263014 233028
rect 189810 232568 189816 232620
rect 189868 232608 189874 232620
rect 222930 232608 222936 232620
rect 189868 232580 222936 232608
rect 189868 232568 189874 232580
rect 222930 232568 222936 232580
rect 222988 232568 222994 232620
rect 328362 232568 328368 232620
rect 328420 232608 328426 232620
rect 345106 232608 345112 232620
rect 328420 232580 345112 232608
rect 328420 232568 328426 232580
rect 345106 232568 345112 232580
rect 345164 232568 345170 232620
rect 169662 232500 169668 232552
rect 169720 232540 169726 232552
rect 418154 232540 418160 232552
rect 169720 232512 418160 232540
rect 169720 232500 169726 232512
rect 418154 232500 418160 232512
rect 418212 232500 418218 232552
rect 418154 231820 418160 231872
rect 418212 231860 418218 231872
rect 419442 231860 419448 231872
rect 418212 231832 419448 231860
rect 418212 231820 418218 231832
rect 419442 231820 419448 231832
rect 419500 231860 419506 231872
rect 580166 231860 580172 231872
rect 419500 231832 580172 231860
rect 419500 231820 419506 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 54846 231752 54852 231804
rect 54904 231792 54910 231804
rect 319254 231792 319260 231804
rect 54904 231764 319260 231792
rect 54904 231752 54910 231764
rect 319254 231752 319260 231764
rect 319312 231752 319318 231804
rect 82814 231684 82820 231736
rect 82872 231724 82878 231736
rect 136634 231724 136640 231736
rect 82872 231696 136640 231724
rect 82872 231684 82878 231696
rect 136634 231684 136640 231696
rect 136692 231684 136698 231736
rect 144362 231684 144368 231736
rect 144420 231724 144426 231736
rect 334066 231724 334072 231736
rect 144420 231696 334072 231724
rect 144420 231684 144426 231696
rect 334066 231684 334072 231696
rect 334124 231684 334130 231736
rect 87046 231616 87052 231668
rect 87104 231656 87110 231668
rect 235350 231656 235356 231668
rect 87104 231628 235356 231656
rect 87104 231616 87110 231628
rect 235350 231616 235356 231628
rect 235408 231616 235414 231668
rect 147122 231548 147128 231600
rect 147180 231588 147186 231600
rect 292574 231588 292580 231600
rect 147180 231560 292580 231588
rect 147180 231548 147186 231560
rect 292574 231548 292580 231560
rect 292632 231548 292638 231600
rect 193030 231140 193036 231192
rect 193088 231180 193094 231192
rect 209130 231180 209136 231192
rect 193088 231152 209136 231180
rect 193088 231140 193094 231152
rect 209130 231140 209136 231152
rect 209188 231140 209194 231192
rect 182082 231072 182088 231124
rect 182140 231112 182146 231124
rect 496814 231112 496820 231124
rect 182140 231084 496820 231112
rect 182140 231072 182146 231084
rect 496814 231072 496820 231084
rect 496872 231072 496878 231124
rect 292574 230936 292580 230988
rect 292632 230976 292638 230988
rect 293218 230976 293224 230988
rect 292632 230948 293224 230976
rect 292632 230936 292638 230948
rect 293218 230936 293224 230948
rect 293276 230936 293282 230988
rect 38562 230392 38568 230444
rect 38620 230432 38626 230444
rect 327350 230432 327356 230444
rect 38620 230404 327356 230432
rect 38620 230392 38626 230404
rect 327350 230392 327356 230404
rect 327408 230432 327414 230444
rect 328362 230432 328368 230444
rect 327408 230404 328368 230432
rect 327408 230392 327414 230404
rect 328362 230392 328368 230404
rect 328420 230392 328426 230444
rect 76650 230324 76656 230376
rect 76708 230364 76714 230376
rect 280154 230364 280160 230376
rect 76708 230336 280160 230364
rect 76708 230324 76714 230336
rect 280154 230324 280160 230336
rect 280212 230364 280218 230376
rect 281442 230364 281448 230376
rect 280212 230336 281448 230364
rect 280212 230324 280218 230336
rect 281442 230324 281448 230336
rect 281500 230324 281506 230376
rect 73798 230256 73804 230308
rect 73856 230296 73862 230308
rect 187694 230296 187700 230308
rect 73856 230268 187700 230296
rect 73856 230256 73862 230268
rect 187694 230256 187700 230268
rect 187752 230256 187758 230308
rect 195330 230256 195336 230308
rect 195388 230296 195394 230308
rect 325694 230296 325700 230308
rect 195388 230268 325700 230296
rect 195388 230256 195394 230268
rect 325694 230256 325700 230268
rect 325752 230256 325758 230308
rect 100202 229848 100208 229900
rect 100260 229888 100266 229900
rect 249058 229888 249064 229900
rect 100260 229860 249064 229888
rect 100260 229848 100266 229860
rect 249058 229848 249064 229860
rect 249116 229848 249122 229900
rect 255958 229848 255964 229900
rect 256016 229888 256022 229900
rect 315942 229888 315948 229900
rect 256016 229860 315948 229888
rect 256016 229848 256022 229860
rect 315942 229848 315948 229860
rect 316000 229848 316006 229900
rect 328362 229848 328368 229900
rect 328420 229888 328426 229900
rect 336734 229888 336740 229900
rect 328420 229860 336740 229888
rect 328420 229848 328426 229860
rect 336734 229848 336740 229860
rect 336792 229848 336798 229900
rect 111886 229780 111892 229832
rect 111944 229820 111950 229832
rect 262858 229820 262864 229832
rect 111944 229792 262864 229820
rect 111944 229780 111950 229792
rect 262858 229780 262864 229792
rect 262916 229780 262922 229832
rect 281442 229780 281448 229832
rect 281500 229820 281506 229832
rect 340230 229820 340236 229832
rect 281500 229792 340236 229820
rect 281500 229780 281506 229792
rect 340230 229780 340236 229792
rect 340288 229780 340294 229832
rect 17218 229712 17224 229764
rect 17276 229752 17282 229764
rect 83550 229752 83556 229764
rect 17276 229724 83556 229752
rect 17276 229712 17282 229724
rect 83550 229712 83556 229724
rect 83608 229712 83614 229764
rect 187694 229712 187700 229764
rect 187752 229752 187758 229764
rect 188798 229752 188804 229764
rect 187752 229724 188804 229752
rect 187752 229712 187758 229724
rect 188798 229712 188804 229724
rect 188856 229752 188862 229764
rect 350626 229752 350632 229764
rect 188856 229724 350632 229752
rect 188856 229712 188862 229724
rect 350626 229712 350632 229724
rect 350684 229712 350690 229764
rect 315942 229100 315948 229152
rect 316000 229140 316006 229152
rect 316770 229140 316776 229152
rect 316000 229112 316776 229140
rect 316000 229100 316006 229112
rect 316770 229100 316776 229112
rect 316828 229100 316834 229152
rect 56318 229032 56324 229084
rect 56376 229072 56382 229084
rect 318058 229072 318064 229084
rect 56376 229044 318064 229072
rect 56376 229032 56382 229044
rect 318058 229032 318064 229044
rect 318116 229032 318122 229084
rect 155586 228964 155592 229016
rect 155644 229004 155650 229016
rect 311894 229004 311900 229016
rect 155644 228976 311900 229004
rect 155644 228964 155650 228976
rect 311894 228964 311900 228976
rect 311952 228964 311958 229016
rect 97626 228896 97632 228948
rect 97684 228936 97690 228948
rect 251818 228936 251824 228948
rect 97684 228908 251824 228936
rect 97684 228896 97690 228908
rect 251818 228896 251824 228908
rect 251876 228896 251882 228948
rect 162302 228828 162308 228880
rect 162360 228868 162366 228880
rect 277394 228868 277400 228880
rect 162360 228840 277400 228868
rect 162360 228828 162366 228840
rect 277394 228828 277400 228840
rect 277452 228828 277458 228880
rect 59078 228352 59084 228404
rect 59136 228392 59142 228404
rect 145650 228392 145656 228404
rect 59136 228364 145656 228392
rect 59136 228352 59142 228364
rect 145650 228352 145656 228364
rect 145708 228352 145714 228404
rect 190270 228352 190276 228404
rect 190328 228392 190334 228404
rect 521654 228392 521660 228404
rect 190328 228364 521660 228392
rect 190328 228352 190334 228364
rect 521654 228352 521660 228364
rect 521712 228352 521718 228404
rect 277394 227740 277400 227792
rect 277452 227780 277458 227792
rect 278038 227780 278044 227792
rect 277452 227752 278044 227780
rect 277452 227740 277458 227752
rect 278038 227740 278044 227752
rect 278096 227740 278102 227792
rect 311894 227740 311900 227792
rect 311952 227780 311958 227792
rect 312538 227780 312544 227792
rect 311952 227752 312544 227780
rect 311952 227740 311958 227752
rect 312538 227740 312544 227752
rect 312596 227740 312602 227792
rect 91738 227672 91744 227724
rect 91796 227712 91802 227724
rect 298738 227712 298744 227724
rect 91796 227684 298744 227712
rect 91796 227672 91802 227684
rect 298738 227672 298744 227684
rect 298796 227672 298802 227724
rect 178954 227604 178960 227656
rect 179012 227644 179018 227656
rect 340138 227644 340144 227656
rect 179012 227616 340144 227644
rect 179012 227604 179018 227616
rect 340138 227604 340144 227616
rect 340196 227604 340202 227656
rect 84378 227536 84384 227588
rect 84436 227576 84442 227588
rect 229738 227576 229744 227588
rect 84436 227548 229744 227576
rect 84436 227536 84442 227548
rect 229738 227536 229744 227548
rect 229796 227536 229802 227588
rect 95050 227468 95056 227520
rect 95108 227508 95114 227520
rect 181530 227508 181536 227520
rect 95108 227480 181536 227508
rect 95108 227468 95114 227480
rect 181530 227468 181536 227480
rect 181588 227468 181594 227520
rect 187602 227060 187608 227112
rect 187660 227100 187666 227112
rect 307018 227100 307024 227112
rect 187660 227072 307024 227100
rect 187660 227060 187666 227072
rect 307018 227060 307024 227072
rect 307076 227060 307082 227112
rect 52086 226992 52092 227044
rect 52144 227032 52150 227044
rect 245010 227032 245016 227044
rect 52144 227004 245016 227032
rect 52144 226992 52150 227004
rect 245010 226992 245016 227004
rect 245068 226992 245074 227044
rect 305638 226992 305644 227044
rect 305696 227032 305702 227044
rect 342898 227032 342904 227044
rect 305696 227004 342904 227032
rect 305696 226992 305702 227004
rect 342898 226992 342904 227004
rect 342956 226992 342962 227044
rect 202690 226312 202696 226364
rect 202748 226352 202754 226364
rect 318058 226352 318064 226364
rect 202748 226324 318064 226352
rect 202748 226312 202754 226324
rect 318058 226312 318064 226324
rect 318116 226312 318122 226364
rect 123754 226244 123760 226296
rect 123812 226284 123818 226296
rect 309134 226284 309140 226296
rect 123812 226256 309140 226284
rect 123812 226244 123818 226256
rect 309134 226244 309140 226256
rect 309192 226244 309198 226296
rect 56226 226176 56232 226228
rect 56284 226216 56290 226228
rect 233234 226216 233240 226228
rect 56284 226188 233240 226216
rect 56284 226176 56290 226188
rect 233234 226176 233240 226188
rect 233292 226176 233298 226228
rect 193858 226108 193864 226160
rect 193916 226148 193922 226160
rect 330018 226148 330024 226160
rect 193916 226120 330024 226148
rect 193916 226108 193922 226120
rect 330018 226108 330024 226120
rect 330076 226108 330082 226160
rect 70486 226040 70492 226092
rect 70544 226080 70550 226092
rect 201494 226080 201500 226092
rect 70544 226052 201500 226080
rect 70544 226040 70550 226052
rect 201494 226040 201500 226052
rect 201552 226080 201558 226092
rect 202690 226080 202696 226092
rect 201552 226052 202696 226080
rect 201552 226040 201558 226052
rect 202690 226040 202696 226052
rect 202748 226040 202754 226092
rect 185670 225700 185676 225752
rect 185728 225740 185734 225752
rect 211798 225740 211804 225752
rect 185728 225712 211804 225740
rect 185728 225700 185734 225712
rect 211798 225700 211804 225712
rect 211856 225700 211862 225752
rect 42702 225632 42708 225684
rect 42760 225672 42766 225684
rect 266446 225672 266452 225684
rect 42760 225644 266452 225672
rect 42760 225632 42766 225644
rect 266446 225632 266452 225644
rect 266504 225632 266510 225684
rect 210234 225564 210240 225616
rect 210292 225604 210298 225616
rect 485130 225604 485136 225616
rect 210292 225576 485136 225604
rect 210292 225564 210298 225576
rect 485130 225564 485136 225576
rect 485188 225564 485194 225616
rect 233234 224952 233240 225004
rect 233292 224992 233298 225004
rect 233878 224992 233884 225004
rect 233292 224964 233884 224992
rect 233292 224952 233298 224964
rect 233878 224952 233884 224964
rect 233936 224952 233942 225004
rect 309134 224952 309140 225004
rect 309192 224992 309198 225004
rect 309870 224992 309876 225004
rect 309192 224964 309876 224992
rect 309192 224952 309198 224964
rect 309870 224952 309876 224964
rect 309928 224952 309934 225004
rect 95234 224884 95240 224936
rect 95292 224924 95298 224936
rect 260834 224924 260840 224936
rect 95292 224896 260840 224924
rect 95292 224884 95298 224896
rect 260834 224884 260840 224896
rect 260892 224924 260898 224936
rect 261478 224924 261484 224936
rect 260892 224896 261484 224924
rect 260892 224884 260898 224896
rect 261478 224884 261484 224896
rect 261536 224884 261542 224936
rect 76006 224816 76012 224868
rect 76064 224856 76070 224868
rect 213914 224856 213920 224868
rect 76064 224828 213920 224856
rect 76064 224816 76070 224828
rect 213914 224816 213920 224828
rect 213972 224816 213978 224868
rect 222930 224816 222936 224868
rect 222988 224856 222994 224868
rect 321646 224856 321652 224868
rect 222988 224828 321652 224856
rect 222988 224816 222994 224828
rect 321646 224816 321652 224828
rect 321704 224816 321710 224868
rect 159542 224748 159548 224800
rect 159600 224788 159606 224800
rect 289814 224788 289820 224800
rect 159600 224760 289820 224788
rect 159600 224748 159606 224760
rect 289814 224748 289820 224760
rect 289872 224788 289878 224800
rect 290458 224788 290464 224800
rect 289872 224760 290464 224788
rect 289872 224748 289878 224760
rect 290458 224748 290464 224760
rect 290516 224748 290522 224800
rect 154022 224680 154028 224732
rect 154080 224720 154086 224732
rect 276014 224720 276020 224732
rect 154080 224692 276020 224720
rect 154080 224680 154086 224692
rect 276014 224680 276020 224692
rect 276072 224720 276078 224732
rect 276658 224720 276664 224732
rect 276072 224692 276664 224720
rect 276072 224680 276078 224692
rect 276658 224680 276664 224692
rect 276716 224680 276722 224732
rect 213914 224408 213920 224460
rect 213972 224448 213978 224460
rect 214558 224448 214564 224460
rect 213972 224420 214564 224448
rect 213972 224408 213978 224420
rect 214558 224408 214564 224420
rect 214616 224408 214622 224460
rect 66070 224272 66076 224324
rect 66128 224312 66134 224324
rect 220078 224312 220084 224324
rect 66128 224284 220084 224312
rect 66128 224272 66134 224284
rect 220078 224272 220084 224284
rect 220136 224272 220142 224324
rect 67450 224204 67456 224256
rect 67508 224244 67514 224256
rect 251174 224244 251180 224256
rect 67508 224216 251180 224244
rect 67508 224204 67514 224216
rect 251174 224204 251180 224216
rect 251232 224204 251238 224256
rect 276658 224204 276664 224256
rect 276716 224244 276722 224256
rect 478874 224244 478880 224256
rect 276716 224216 478880 224244
rect 276716 224204 276722 224216
rect 478874 224204 478880 224216
rect 478932 224204 478938 224256
rect 247034 223592 247040 223644
rect 247092 223632 247098 223644
rect 318150 223632 318156 223644
rect 247092 223604 318156 223632
rect 247092 223592 247098 223604
rect 318150 223592 318156 223604
rect 318208 223592 318214 223644
rect 102226 223524 102232 223576
rect 102284 223564 102290 223576
rect 273254 223564 273260 223576
rect 102284 223536 273260 223564
rect 102284 223524 102290 223536
rect 273254 223524 273260 223536
rect 273312 223564 273318 223576
rect 273990 223564 273996 223576
rect 273312 223536 273996 223564
rect 273312 223524 273318 223536
rect 273990 223524 273996 223536
rect 274048 223524 274054 223576
rect 93946 223456 93952 223508
rect 94004 223496 94010 223508
rect 247034 223496 247040 223508
rect 94004 223468 247040 223496
rect 94004 223456 94010 223468
rect 247034 223456 247040 223468
rect 247092 223456 247098 223508
rect 170582 223388 170588 223440
rect 170640 223428 170646 223440
rect 238754 223428 238760 223440
rect 170640 223400 238760 223428
rect 170640 223388 170646 223400
rect 238754 223388 238760 223400
rect 238812 223428 238818 223440
rect 239490 223428 239496 223440
rect 238812 223400 239496 223428
rect 238812 223388 238818 223400
rect 239490 223388 239496 223400
rect 239548 223388 239554 223440
rect 68738 222912 68744 222964
rect 68796 222952 68802 222964
rect 253934 222952 253940 222964
rect 68796 222924 253940 222952
rect 68796 222912 68802 222924
rect 253934 222912 253940 222924
rect 253992 222912 253998 222964
rect 183462 222844 183468 222896
rect 183520 222884 183526 222896
rect 475470 222884 475476 222896
rect 183520 222856 475476 222884
rect 183520 222844 183526 222856
rect 475470 222844 475476 222856
rect 475528 222844 475534 222896
rect 195974 222164 195980 222216
rect 196032 222204 196038 222216
rect 196802 222204 196808 222216
rect 196032 222176 196808 222204
rect 196032 222164 196038 222176
rect 196802 222164 196808 222176
rect 196860 222204 196866 222216
rect 347866 222204 347872 222216
rect 196860 222176 347872 222204
rect 196860 222164 196866 222176
rect 347866 222164 347872 222176
rect 347924 222164 347930 222216
rect 69198 222096 69204 222148
rect 69256 222136 69262 222148
rect 256694 222136 256700 222148
rect 69256 222108 256700 222136
rect 69256 222096 69262 222108
rect 256694 222096 256700 222108
rect 256752 222096 256758 222148
rect 163682 222028 163688 222080
rect 163740 222068 163746 222080
rect 300118 222068 300124 222080
rect 163740 222040 300124 222068
rect 163740 222028 163746 222040
rect 300118 222028 300124 222040
rect 300176 222028 300182 222080
rect 74626 221960 74632 222012
rect 74684 222000 74690 222012
rect 195974 222000 195980 222012
rect 74684 221972 195980 222000
rect 74684 221960 74690 221972
rect 195974 221960 195980 221972
rect 196032 221960 196038 222012
rect 256694 221960 256700 222012
rect 256752 222000 256758 222012
rect 257338 222000 257344 222012
rect 256752 221972 257344 222000
rect 256752 221960 256758 221972
rect 257338 221960 257344 221972
rect 257396 221960 257402 222012
rect 195238 221552 195244 221604
rect 195296 221592 195302 221604
rect 278774 221592 278780 221604
rect 195296 221564 278780 221592
rect 195296 221552 195302 221564
rect 278774 221552 278780 221564
rect 278832 221552 278838 221604
rect 49418 221484 49424 221536
rect 49476 221524 49482 221536
rect 232590 221524 232596 221536
rect 49476 221496 232596 221524
rect 49476 221484 49482 221496
rect 232590 221484 232596 221496
rect 232648 221484 232654 221536
rect 175182 221416 175188 221468
rect 175240 221456 175246 221468
rect 510706 221456 510712 221468
rect 175240 221428 510712 221456
rect 175240 221416 175246 221428
rect 510706 221416 510712 221428
rect 510764 221416 510770 221468
rect 323578 220844 323584 220856
rect 322952 220816 323584 220844
rect 142982 220736 142988 220788
rect 143040 220776 143046 220788
rect 322952 220776 322980 220816
rect 323578 220804 323584 220816
rect 323636 220844 323642 220856
rect 347958 220844 347964 220856
rect 323636 220816 347964 220844
rect 323636 220804 323642 220816
rect 347958 220804 347964 220816
rect 348016 220804 348022 220856
rect 143040 220748 322980 220776
rect 143040 220736 143046 220748
rect 158070 220668 158076 220720
rect 158128 220708 158134 220720
rect 332686 220708 332692 220720
rect 158128 220680 332692 220708
rect 158128 220668 158134 220680
rect 332686 220668 332692 220680
rect 332744 220668 332750 220720
rect 177482 220260 177488 220312
rect 177540 220300 177546 220312
rect 232498 220300 232504 220312
rect 177540 220272 232504 220300
rect 177540 220260 177546 220272
rect 232498 220260 232504 220272
rect 232556 220260 232562 220312
rect 101490 220192 101496 220244
rect 101548 220232 101554 220244
rect 255314 220232 255320 220244
rect 101548 220204 255320 220232
rect 101548 220192 101554 220204
rect 255314 220192 255320 220204
rect 255372 220192 255378 220244
rect 57698 220124 57704 220176
rect 57756 220164 57762 220176
rect 277394 220164 277400 220176
rect 57756 220136 277400 220164
rect 57756 220124 57762 220136
rect 277394 220124 277400 220136
rect 277452 220124 277458 220176
rect 181622 220056 181628 220108
rect 181680 220096 181686 220108
rect 417418 220096 417424 220108
rect 181680 220068 417424 220096
rect 181680 220056 181686 220068
rect 417418 220056 417424 220068
rect 417476 220056 417482 220108
rect 148502 219376 148508 219428
rect 148560 219416 148566 219428
rect 335446 219416 335452 219428
rect 148560 219388 335452 219416
rect 148560 219376 148566 219388
rect 335446 219376 335452 219388
rect 335504 219376 335510 219428
rect 84286 219308 84292 219360
rect 84344 219348 84350 219360
rect 229094 219348 229100 219360
rect 84344 219320 229100 219348
rect 84344 219308 84350 219320
rect 229094 219308 229100 219320
rect 229152 219348 229158 219360
rect 230382 219348 230388 219360
rect 229152 219320 230388 219348
rect 229152 219308 229158 219320
rect 230382 219308 230388 219320
rect 230440 219308 230446 219360
rect 86218 219240 86224 219292
rect 86276 219280 86282 219292
rect 208394 219280 208400 219292
rect 86276 219252 208400 219280
rect 86276 219240 86282 219252
rect 208394 219240 208400 219252
rect 208452 219240 208458 219292
rect 475378 218900 475384 218952
rect 475436 218940 475442 218952
rect 480254 218940 480260 218952
rect 475436 218912 480260 218940
rect 475436 218900 475442 218912
rect 480254 218900 480260 218912
rect 480312 218900 480318 218952
rect 230382 218832 230388 218884
rect 230440 218872 230446 218884
rect 291930 218872 291936 218884
rect 230440 218844 291936 218872
rect 230440 218832 230446 218844
rect 291930 218832 291936 218844
rect 291988 218832 291994 218884
rect 156690 218764 156696 218816
rect 156748 218804 156754 218816
rect 238018 218804 238024 218816
rect 156748 218776 238024 218804
rect 156748 218764 156754 218776
rect 238018 218764 238024 218776
rect 238076 218764 238082 218816
rect 140130 218696 140136 218748
rect 140188 218736 140194 218748
rect 258166 218736 258172 218748
rect 140188 218708 258172 218736
rect 140188 218696 140194 218708
rect 258166 218696 258172 218708
rect 258224 218696 258230 218748
rect 483658 218696 483664 218748
rect 483716 218736 483722 218748
rect 514846 218736 514852 218748
rect 483716 218708 514852 218736
rect 483716 218696 483722 218708
rect 514846 218696 514852 218708
rect 514904 218696 514910 218748
rect 208394 218016 208400 218068
rect 208452 218056 208458 218068
rect 209222 218056 209228 218068
rect 208452 218028 209228 218056
rect 208452 218016 208458 218028
rect 209222 218016 209228 218028
rect 209280 218016 209286 218068
rect 220722 218016 220728 218068
rect 220780 218056 220786 218068
rect 346486 218056 346492 218068
rect 220780 218028 346492 218056
rect 220780 218016 220786 218028
rect 346486 218016 346492 218028
rect 346544 218016 346550 218068
rect 514846 218016 514852 218068
rect 514904 218056 514910 218068
rect 580166 218056 580172 218068
rect 514904 218028 580172 218056
rect 514904 218016 514910 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 110506 217948 110512 218000
rect 110564 217988 110570 218000
rect 140774 217988 140780 218000
rect 110564 217960 140780 217988
rect 110564 217948 110570 217960
rect 140774 217948 140780 217960
rect 140832 217988 140838 218000
rect 335998 217988 336004 218000
rect 140832 217960 336004 217988
rect 140832 217948 140838 217960
rect 335998 217948 336004 217960
rect 336056 217948 336062 218000
rect 78766 217880 78772 217932
rect 78824 217920 78830 217932
rect 219434 217920 219440 217932
rect 78824 217892 219440 217920
rect 78824 217880 78830 217892
rect 219434 217880 219440 217892
rect 219492 217920 219498 217932
rect 220722 217920 220728 217932
rect 219492 217892 220728 217920
rect 219492 217880 219498 217892
rect 220722 217880 220728 217892
rect 220780 217880 220786 217932
rect 198918 217404 198924 217456
rect 198976 217444 198982 217456
rect 324498 217444 324504 217456
rect 198976 217416 324504 217444
rect 198976 217404 198982 217416
rect 324498 217404 324504 217416
rect 324556 217404 324562 217456
rect 130470 217336 130476 217388
rect 130528 217376 130534 217388
rect 263594 217376 263600 217388
rect 130528 217348 263600 217376
rect 130528 217336 130534 217348
rect 263594 217336 263600 217348
rect 263652 217336 263658 217388
rect 170490 217268 170496 217320
rect 170548 217308 170554 217320
rect 367094 217308 367100 217320
rect 170548 217280 367100 217308
rect 170548 217268 170554 217280
rect 367094 217268 367100 217280
rect 367152 217268 367158 217320
rect 53558 216588 53564 216640
rect 53616 216628 53622 216640
rect 312630 216628 312636 216640
rect 53616 216600 312636 216628
rect 53616 216588 53622 216600
rect 312630 216588 312636 216600
rect 312688 216588 312694 216640
rect 92566 216520 92572 216572
rect 92624 216560 92630 216572
rect 246298 216560 246304 216572
rect 92624 216532 246304 216560
rect 92624 216520 92630 216532
rect 246298 216520 246304 216532
rect 246356 216520 246362 216572
rect 152550 216044 152556 216096
rect 152608 216084 152614 216096
rect 240778 216084 240784 216096
rect 152608 216056 240784 216084
rect 152608 216044 152614 216056
rect 240778 216044 240784 216056
rect 240836 216044 240842 216096
rect 145650 215976 145656 216028
rect 145708 216016 145714 216028
rect 274726 216016 274732 216028
rect 145708 215988 274732 216016
rect 145708 215976 145714 215988
rect 274726 215976 274732 215988
rect 274784 215976 274790 216028
rect 184750 215908 184756 215960
rect 184808 215948 184814 215960
rect 446490 215948 446496 215960
rect 184808 215920 446496 215948
rect 184808 215908 184814 215920
rect 446490 215908 446496 215920
rect 446548 215908 446554 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 21358 215268 21364 215280
rect 3384 215240 21364 215268
rect 3384 215228 3390 215240
rect 21358 215228 21364 215240
rect 21416 215228 21422 215280
rect 118694 215228 118700 215280
rect 118752 215268 118758 215280
rect 307110 215268 307116 215280
rect 118752 215240 307116 215268
rect 118752 215228 118758 215240
rect 307110 215228 307116 215240
rect 307168 215228 307174 215280
rect 186130 214820 186136 214872
rect 186188 214860 186194 214872
rect 240870 214860 240876 214872
rect 186188 214832 240876 214860
rect 186188 214820 186194 214832
rect 240870 214820 240876 214832
rect 240928 214820 240934 214872
rect 93854 214752 93860 214804
rect 93912 214792 93918 214804
rect 246390 214792 246396 214804
rect 93912 214764 246396 214792
rect 93912 214752 93918 214764
rect 246390 214752 246396 214764
rect 246448 214752 246454 214804
rect 53650 214684 53656 214736
rect 53708 214724 53714 214736
rect 235258 214724 235264 214736
rect 53708 214696 235264 214724
rect 53708 214684 53714 214696
rect 235258 214684 235264 214696
rect 235316 214684 235322 214736
rect 233878 214616 233884 214668
rect 233936 214656 233942 214668
rect 486418 214656 486424 214668
rect 233936 214628 486424 214656
rect 233936 214616 233942 214628
rect 486418 214616 486424 214628
rect 486476 214616 486482 214668
rect 176562 214548 176568 214600
rect 176620 214588 176626 214600
rect 502978 214588 502984 214600
rect 176620 214560 502984 214588
rect 176620 214548 176626 214560
rect 502978 214548 502984 214560
rect 503036 214548 503042 214600
rect 72418 213868 72424 213920
rect 72476 213908 72482 213920
rect 258074 213908 258080 213920
rect 72476 213880 258080 213908
rect 72476 213868 72482 213880
rect 258074 213868 258080 213880
rect 258132 213908 258138 213920
rect 259362 213908 259368 213920
rect 258132 213880 259368 213908
rect 258132 213868 258138 213880
rect 259362 213868 259368 213880
rect 259420 213868 259426 213920
rect 103698 213800 103704 213852
rect 103756 213840 103762 213852
rect 271874 213840 271880 213852
rect 103756 213812 271880 213840
rect 103756 213800 103762 213812
rect 271874 213800 271880 213812
rect 271932 213840 271938 213852
rect 272518 213840 272524 213852
rect 271932 213812 272524 213840
rect 271932 213800 271938 213812
rect 272518 213800 272524 213812
rect 272576 213800 272582 213852
rect 80054 213732 80060 213784
rect 80112 213772 80118 213784
rect 221458 213772 221464 213784
rect 80112 213744 221464 213772
rect 80112 213732 80118 213744
rect 221458 213732 221464 213744
rect 221516 213732 221522 213784
rect 182910 213324 182916 213376
rect 182968 213364 182974 213376
rect 267734 213364 267740 213376
rect 182968 213336 267740 213364
rect 182968 213324 182974 213336
rect 267734 213324 267740 213336
rect 267792 213324 267798 213376
rect 127618 213256 127624 213308
rect 127676 213296 127682 213308
rect 236638 213296 236644 213308
rect 127676 213268 236644 213296
rect 127676 213256 127682 213268
rect 236638 213256 236644 213268
rect 236696 213256 236702 213308
rect 187510 213188 187516 213240
rect 187568 213228 187574 213240
rect 407758 213228 407764 213240
rect 187568 213200 407764 213228
rect 187568 213188 187574 213200
rect 407758 213188 407764 213200
rect 407816 213188 407822 213240
rect 114554 212440 114560 212492
rect 114612 212480 114618 212492
rect 295334 212480 295340 212492
rect 114612 212452 295340 212480
rect 114612 212440 114618 212452
rect 295334 212440 295340 212452
rect 295392 212440 295398 212492
rect 88978 212372 88984 212424
rect 89036 212412 89042 212424
rect 224954 212412 224960 212424
rect 89036 212384 224960 212412
rect 89036 212372 89042 212384
rect 224954 212372 224960 212384
rect 225012 212412 225018 212424
rect 225598 212412 225604 212424
rect 225012 212384 225604 212412
rect 225012 212372 225018 212384
rect 225598 212372 225604 212384
rect 225656 212372 225662 212424
rect 295334 212032 295340 212084
rect 295392 212072 295398 212084
rect 295978 212072 295984 212084
rect 295392 212044 295984 212072
rect 295392 212032 295398 212044
rect 295978 212032 295984 212044
rect 296036 212032 296042 212084
rect 153838 211964 153844 212016
rect 153896 212004 153902 212016
rect 286318 212004 286324 212016
rect 153896 211976 286324 212004
rect 153896 211964 153902 211976
rect 286318 211964 286324 211976
rect 286376 211964 286382 212016
rect 102134 211896 102140 211948
rect 102192 211936 102198 211948
rect 249978 211936 249984 211948
rect 102192 211908 249984 211936
rect 102192 211896 102198 211908
rect 249978 211896 249984 211908
rect 250036 211896 250042 211948
rect 259362 211896 259368 211948
rect 259420 211936 259426 211948
rect 341518 211936 341524 211948
rect 259420 211908 341524 211936
rect 259420 211896 259426 211908
rect 341518 211896 341524 211908
rect 341576 211896 341582 211948
rect 126422 211828 126428 211880
rect 126480 211868 126486 211880
rect 277486 211868 277492 211880
rect 126480 211840 277492 211868
rect 126480 211828 126486 211840
rect 277486 211828 277492 211840
rect 277544 211828 277550 211880
rect 173342 211760 173348 211812
rect 173400 211800 173406 211812
rect 507854 211800 507860 211812
rect 173400 211772 507860 211800
rect 173400 211760 173406 211772
rect 507854 211760 507860 211772
rect 507912 211760 507918 211812
rect 319530 211188 319536 211200
rect 287026 211160 319536 211188
rect 107746 211080 107752 211132
rect 107804 211120 107810 211132
rect 285674 211120 285680 211132
rect 107804 211092 285680 211120
rect 107804 211080 107810 211092
rect 285674 211080 285680 211092
rect 285732 211120 285738 211132
rect 287026 211120 287054 211160
rect 319530 211148 319536 211160
rect 319588 211148 319594 211200
rect 285732 211092 287054 211120
rect 285732 211080 285738 211092
rect 432598 211080 432604 211132
rect 432656 211120 432662 211132
rect 446398 211120 446404 211132
rect 432656 211092 446404 211120
rect 432656 211080 432662 211092
rect 446398 211080 446404 211092
rect 446456 211080 446462 211132
rect 431954 210672 431960 210724
rect 432012 210712 432018 210724
rect 432598 210712 432604 210724
rect 432012 210684 432604 210712
rect 432012 210672 432018 210684
rect 432598 210672 432604 210684
rect 432656 210672 432662 210724
rect 136082 210536 136088 210588
rect 136140 210576 136146 210588
rect 262214 210576 262220 210588
rect 136140 210548 262220 210576
rect 136140 210536 136146 210548
rect 262214 210536 262220 210548
rect 262272 210536 262278 210588
rect 43806 210468 43812 210520
rect 43864 210508 43870 210520
rect 239398 210508 239404 210520
rect 43864 210480 239404 210508
rect 43864 210468 43870 210480
rect 239398 210468 239404 210480
rect 239456 210468 239462 210520
rect 7558 210400 7564 210452
rect 7616 210440 7622 210452
rect 110506 210440 110512 210452
rect 7616 210412 110512 210440
rect 7616 210400 7622 210412
rect 110506 210400 110512 210412
rect 110564 210400 110570 210452
rect 167638 210400 167644 210452
rect 167696 210440 167702 210452
rect 231118 210440 231124 210452
rect 167696 210412 231124 210440
rect 167696 210400 167702 210412
rect 231118 210400 231124 210412
rect 231176 210400 231182 210452
rect 237374 210400 237380 210452
rect 237432 210440 237438 210452
rect 483014 210440 483020 210452
rect 237432 210412 483020 210440
rect 237432 210400 237438 210412
rect 483014 210400 483020 210412
rect 483072 210400 483078 210452
rect 422294 209992 422300 210044
rect 422352 210032 422358 210044
rect 425698 210032 425704 210044
rect 422352 210004 425704 210032
rect 422352 209992 422358 210004
rect 425698 209992 425704 210004
rect 425756 209992 425762 210044
rect 105538 209720 105544 209772
rect 105596 209760 105602 209772
rect 266354 209760 266360 209772
rect 105596 209732 266360 209760
rect 105596 209720 105602 209732
rect 266354 209720 266360 209732
rect 266412 209720 266418 209772
rect 162210 209176 162216 209228
rect 162268 209216 162274 209228
rect 226978 209216 226984 209228
rect 162268 209188 226984 209216
rect 162268 209176 162274 209188
rect 226978 209176 226984 209188
rect 227036 209176 227042 209228
rect 159450 209108 159456 209160
rect 159508 209148 159514 209160
rect 273898 209148 273904 209160
rect 159508 209120 273904 209148
rect 159508 209108 159514 209120
rect 273898 209108 273904 209120
rect 273956 209108 273962 209160
rect 56134 209040 56140 209092
rect 56192 209080 56198 209092
rect 222930 209080 222936 209092
rect 56192 209052 222936 209080
rect 56192 209040 56198 209052
rect 222930 209040 222936 209052
rect 222988 209040 222994 209092
rect 239490 209040 239496 209092
rect 239548 209080 239554 209092
rect 513282 209080 513288 209092
rect 239548 209052 513288 209080
rect 239548 209040 239554 209052
rect 513282 209040 513288 209052
rect 513340 209040 513346 209092
rect 266354 208360 266360 208412
rect 266412 208400 266418 208412
rect 266998 208400 267004 208412
rect 266412 208372 267004 208400
rect 266412 208360 266418 208372
rect 266998 208360 267004 208372
rect 267056 208360 267062 208412
rect 99374 208292 99380 208344
rect 99432 208332 99438 208344
rect 269114 208332 269120 208344
rect 99432 208304 269120 208332
rect 99432 208292 99438 208304
rect 269114 208292 269120 208304
rect 269172 208292 269178 208344
rect 196618 207816 196624 207868
rect 196676 207856 196682 207868
rect 280154 207856 280160 207868
rect 196676 207828 280160 207856
rect 196676 207816 196682 207828
rect 280154 207816 280160 207828
rect 280212 207816 280218 207868
rect 77294 207748 77300 207800
rect 77352 207788 77358 207800
rect 252830 207788 252836 207800
rect 77352 207760 252836 207788
rect 77352 207748 77358 207760
rect 252830 207748 252836 207760
rect 252888 207748 252894 207800
rect 272518 207748 272524 207800
rect 272576 207788 272582 207800
rect 325694 207788 325700 207800
rect 272576 207760 325700 207788
rect 272576 207748 272582 207760
rect 325694 207748 325700 207760
rect 325752 207748 325758 207800
rect 46750 207680 46756 207732
rect 46808 207720 46814 207732
rect 276014 207720 276020 207732
rect 46808 207692 276020 207720
rect 46808 207680 46814 207692
rect 276014 207680 276020 207692
rect 276072 207680 276078 207732
rect 194410 207612 194416 207664
rect 194468 207652 194474 207664
rect 517606 207652 517612 207664
rect 194468 207624 517612 207652
rect 194468 207612 194474 207624
rect 517606 207612 517612 207624
rect 517664 207612 517670 207664
rect 269114 207000 269120 207052
rect 269172 207040 269178 207052
rect 269758 207040 269764 207052
rect 269172 207012 269764 207040
rect 269172 207000 269178 207012
rect 269758 207000 269764 207012
rect 269816 207000 269822 207052
rect 149698 206456 149704 206508
rect 149756 206496 149762 206508
rect 196618 206496 196624 206508
rect 149756 206468 196624 206496
rect 149756 206456 149762 206468
rect 196618 206456 196624 206468
rect 196676 206456 196682 206508
rect 122190 206388 122196 206440
rect 122248 206428 122254 206440
rect 252738 206428 252744 206440
rect 122248 206400 252744 206428
rect 122248 206388 122254 206400
rect 252738 206388 252744 206400
rect 252796 206388 252802 206440
rect 74534 206320 74540 206372
rect 74592 206360 74598 206372
rect 254026 206360 254032 206372
rect 74592 206332 254032 206360
rect 74592 206320 74598 206332
rect 254026 206320 254032 206332
rect 254084 206320 254090 206372
rect 262950 206320 262956 206372
rect 263008 206360 263014 206372
rect 505186 206360 505192 206372
rect 263008 206332 505192 206360
rect 263008 206320 263014 206332
rect 505186 206320 505192 206332
rect 505244 206320 505250 206372
rect 180702 206252 180708 206304
rect 180760 206292 180766 206304
rect 436094 206292 436100 206304
rect 180760 206264 436100 206292
rect 180760 206252 180766 206264
rect 436094 206252 436100 206264
rect 436152 206252 436158 206304
rect 512638 206252 512644 206304
rect 512696 206292 512702 206304
rect 513282 206292 513288 206304
rect 512696 206264 513288 206292
rect 512696 206252 512702 206264
rect 513282 206252 513288 206264
rect 513340 206292 513346 206304
rect 580166 206292 580172 206304
rect 513340 206264 580172 206292
rect 513340 206252 513346 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 107654 205572 107660 205624
rect 107712 205612 107718 205624
rect 284294 205612 284300 205624
rect 107712 205584 284300 205612
rect 107712 205572 107718 205584
rect 284294 205572 284300 205584
rect 284352 205572 284358 205624
rect 140038 205096 140044 205148
rect 140096 205136 140102 205148
rect 195238 205136 195244 205148
rect 140096 205108 195244 205136
rect 140096 205096 140102 205108
rect 195238 205096 195244 205108
rect 195296 205096 195302 205148
rect 284294 205096 284300 205148
rect 284352 205136 284358 205148
rect 284938 205136 284944 205148
rect 284352 205108 284944 205136
rect 284352 205096 284358 205108
rect 284938 205096 284944 205108
rect 284996 205096 285002 205148
rect 89806 205028 89812 205080
rect 89864 205068 89870 205080
rect 228358 205068 228364 205080
rect 89864 205040 228364 205068
rect 89864 205028 89870 205040
rect 228358 205028 228364 205040
rect 228416 205028 228422 205080
rect 76558 204960 76564 205012
rect 76616 205000 76622 205012
rect 263686 205000 263692 205012
rect 76616 204972 263692 205000
rect 76616 204960 76622 204972
rect 263686 204960 263692 204972
rect 263744 204960 263750 205012
rect 188890 204892 188896 204944
rect 188948 204932 188954 204944
rect 400858 204932 400864 204944
rect 188948 204904 400864 204932
rect 188948 204892 188954 204904
rect 400858 204892 400864 204904
rect 400916 204892 400922 204944
rect 97994 204212 98000 204264
rect 98052 204252 98058 204264
rect 147674 204252 147680 204264
rect 98052 204224 147680 204252
rect 98052 204212 98058 204224
rect 147674 204212 147680 204224
rect 147732 204252 147738 204264
rect 148318 204252 148324 204264
rect 147732 204224 148324 204252
rect 147732 204212 147738 204224
rect 148318 204212 148324 204224
rect 148376 204212 148382 204264
rect 429838 204212 429844 204264
rect 429896 204252 429902 204264
rect 431218 204252 431224 204264
rect 429896 204224 431224 204252
rect 429896 204212 429902 204224
rect 431218 204212 431224 204224
rect 431276 204212 431282 204264
rect 147030 203736 147036 203788
rect 147088 203776 147094 203788
rect 233878 203776 233884 203788
rect 147088 203748 233884 203776
rect 147088 203736 147094 203748
rect 233878 203736 233884 203748
rect 233936 203736 233942 203788
rect 96614 203668 96620 203720
rect 96672 203708 96678 203720
rect 259454 203708 259460 203720
rect 96672 203680 259460 203708
rect 96672 203668 96678 203680
rect 259454 203668 259460 203680
rect 259512 203668 259518 203720
rect 111794 203600 111800 203652
rect 111852 203640 111858 203652
rect 276106 203640 276112 203652
rect 111852 203612 276112 203640
rect 111852 203600 111858 203612
rect 276106 203600 276112 203612
rect 276164 203600 276170 203652
rect 293218 203600 293224 203652
rect 293276 203640 293282 203652
rect 429838 203640 429844 203652
rect 293276 203612 429844 203640
rect 293276 203600 293282 203612
rect 429838 203600 429844 203612
rect 429896 203600 429902 203652
rect 147674 203532 147680 203584
rect 147732 203572 147738 203584
rect 399478 203572 399484 203584
rect 147732 203544 399484 203572
rect 147732 203532 147738 203544
rect 399478 203532 399484 203544
rect 399536 203532 399542 203584
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 120166 202824 120172 202836
rect 3476 202796 120172 202824
rect 3476 202784 3482 202796
rect 120166 202784 120172 202796
rect 120224 202784 120230 202836
rect 198550 202376 198556 202428
rect 198608 202416 198614 202428
rect 321554 202416 321560 202428
rect 198608 202388 321560 202416
rect 198608 202376 198614 202388
rect 321554 202376 321560 202388
rect 321612 202376 321618 202428
rect 115934 202308 115940 202360
rect 115992 202348 115998 202360
rect 245102 202348 245108 202360
rect 115992 202320 245108 202348
rect 115992 202308 115998 202320
rect 245102 202308 245108 202320
rect 245160 202308 245166 202360
rect 137278 202240 137284 202292
rect 137336 202280 137342 202292
rect 349246 202280 349252 202292
rect 137336 202252 349252 202280
rect 137336 202240 137342 202252
rect 349246 202240 349252 202252
rect 349304 202240 349310 202292
rect 55030 202172 55036 202224
rect 55088 202212 55094 202224
rect 269114 202212 269120 202224
rect 55088 202184 269120 202212
rect 55088 202172 55094 202184
rect 269114 202172 269120 202184
rect 269172 202172 269178 202224
rect 144270 202104 144276 202156
rect 144328 202144 144334 202156
rect 396718 202144 396724 202156
rect 144328 202116 396724 202144
rect 144328 202104 144334 202116
rect 396718 202104 396724 202116
rect 396776 202104 396782 202156
rect 157978 201016 157984 201068
rect 158036 201056 158042 201068
rect 213270 201056 213276 201068
rect 158036 201028 213276 201056
rect 158036 201016 158042 201028
rect 213270 201016 213276 201028
rect 213328 201016 213334 201068
rect 211798 200948 211804 201000
rect 211856 200988 211862 201000
rect 313918 200988 313924 201000
rect 211856 200960 313924 200988
rect 211856 200948 211862 200960
rect 313918 200948 313924 200960
rect 313976 200948 313982 201000
rect 191742 200880 191748 200932
rect 191800 200920 191806 200932
rect 296070 200920 296076 200932
rect 191800 200892 296076 200920
rect 191800 200880 191806 200892
rect 296070 200880 296076 200892
rect 296128 200880 296134 200932
rect 141510 200812 141516 200864
rect 141568 200852 141574 200864
rect 273254 200852 273260 200864
rect 141568 200824 273260 200852
rect 141568 200812 141574 200824
rect 273254 200812 273260 200824
rect 273312 200812 273318 200864
rect 166258 200744 166264 200796
rect 166316 200784 166322 200796
rect 199470 200784 199476 200796
rect 166316 200756 199476 200784
rect 166316 200744 166322 200756
rect 199470 200744 199476 200756
rect 199528 200744 199534 200796
rect 204898 200744 204904 200796
rect 204956 200784 204962 200796
rect 513374 200784 513380 200796
rect 204956 200756 513380 200784
rect 204956 200744 204962 200756
rect 513374 200744 513380 200756
rect 513432 200744 513438 200796
rect 155494 199588 155500 199640
rect 155552 199628 155558 199640
rect 238110 199628 238116 199640
rect 155552 199600 238116 199628
rect 155552 199588 155558 199600
rect 238110 199588 238116 199600
rect 238168 199588 238174 199640
rect 133138 199520 133144 199572
rect 133196 199560 133202 199572
rect 216030 199560 216036 199572
rect 133196 199532 216036 199560
rect 133196 199520 133202 199532
rect 216030 199520 216036 199532
rect 216088 199520 216094 199572
rect 177942 199452 177948 199504
rect 178000 199492 178006 199504
rect 338114 199492 338120 199504
rect 178000 199464 338120 199492
rect 178000 199452 178006 199464
rect 338114 199452 338120 199464
rect 338172 199452 338178 199504
rect 86954 199384 86960 199436
rect 87012 199424 87018 199436
rect 267826 199424 267832 199436
rect 87012 199396 267832 199424
rect 87012 199384 87018 199396
rect 267826 199384 267832 199396
rect 267884 199384 267890 199436
rect 300118 199384 300124 199436
rect 300176 199424 300182 199436
rect 509326 199424 509332 199436
rect 300176 199396 509332 199424
rect 300176 199384 300182 199396
rect 509326 199384 509332 199396
rect 509384 199384 509390 199436
rect 144178 198092 144184 198144
rect 144236 198132 144242 198144
rect 289170 198132 289176 198144
rect 144236 198104 289176 198132
rect 144236 198092 144242 198104
rect 289170 198092 289176 198104
rect 289228 198092 289234 198144
rect 83458 198024 83464 198076
rect 83516 198064 83522 198076
rect 232682 198064 232688 198076
rect 83516 198036 232688 198064
rect 83516 198024 83522 198036
rect 232682 198024 232688 198036
rect 232740 198024 232746 198076
rect 172422 197956 172428 198008
rect 172480 197996 172486 198008
rect 200758 197996 200764 198008
rect 172480 197968 200764 197996
rect 172480 197956 172486 197968
rect 200758 197956 200764 197968
rect 200816 197956 200822 198008
rect 218698 197956 218704 198008
rect 218756 197996 218762 198008
rect 516134 197996 516140 198008
rect 218756 197968 516140 197996
rect 218756 197956 218762 197968
rect 516134 197956 516140 197968
rect 516192 197956 516198 198008
rect 189718 196800 189724 196852
rect 189776 196840 189782 196852
rect 281534 196840 281540 196852
rect 189776 196812 281540 196840
rect 189776 196800 189782 196812
rect 281534 196800 281540 196812
rect 281592 196800 281598 196852
rect 151078 196732 151084 196784
rect 151136 196772 151142 196784
rect 291838 196772 291844 196784
rect 151136 196744 291844 196772
rect 151136 196732 151142 196744
rect 291838 196732 291844 196744
rect 291896 196732 291902 196784
rect 295978 196732 295984 196784
rect 296036 196772 296042 196784
rect 327166 196772 327172 196784
rect 296036 196744 327172 196772
rect 296036 196732 296042 196744
rect 327166 196732 327172 196744
rect 327224 196732 327230 196784
rect 138658 196664 138664 196716
rect 138716 196704 138722 196716
rect 351178 196704 351184 196716
rect 138716 196676 351184 196704
rect 138716 196664 138722 196676
rect 351178 196664 351184 196676
rect 351236 196664 351242 196716
rect 124950 196596 124956 196648
rect 125008 196636 125014 196648
rect 265158 196636 265164 196648
rect 125008 196608 265164 196636
rect 125008 196596 125014 196608
rect 265158 196596 265164 196608
rect 265216 196596 265222 196648
rect 278038 196596 278044 196648
rect 278096 196636 278102 196648
rect 506566 196636 506572 196648
rect 278096 196608 506572 196636
rect 278096 196596 278102 196608
rect 506566 196596 506572 196608
rect 506624 196596 506630 196648
rect 235350 195440 235356 195492
rect 235408 195480 235414 195492
rect 309778 195480 309784 195492
rect 235408 195452 309784 195480
rect 235408 195440 235414 195452
rect 309778 195440 309784 195452
rect 309836 195440 309842 195492
rect 178862 195372 178868 195424
rect 178920 195412 178926 195424
rect 314010 195412 314016 195424
rect 178920 195384 314016 195412
rect 178920 195372 178926 195384
rect 314010 195372 314016 195384
rect 314068 195372 314074 195424
rect 89714 195304 89720 195356
rect 89772 195344 89778 195356
rect 254118 195344 254124 195356
rect 89772 195316 254124 195344
rect 89772 195304 89778 195316
rect 254118 195304 254124 195316
rect 254176 195304 254182 195356
rect 257338 195304 257344 195356
rect 257396 195344 257402 195356
rect 325970 195344 325976 195356
rect 257396 195316 325976 195344
rect 257396 195304 257402 195316
rect 325970 195304 325976 195316
rect 326028 195304 326034 195356
rect 145558 195236 145564 195288
rect 145616 195276 145622 195288
rect 199378 195276 199384 195288
rect 145616 195248 199384 195276
rect 145616 195236 145622 195248
rect 199378 195236 199384 195248
rect 199436 195236 199442 195288
rect 213178 195236 213184 195288
rect 213236 195276 213242 195288
rect 503806 195276 503812 195288
rect 213236 195248 503812 195276
rect 213236 195236 213242 195248
rect 503806 195236 503812 195248
rect 503864 195236 503870 195288
rect 217318 194080 217324 194132
rect 217376 194120 217382 194132
rect 321646 194120 321652 194132
rect 217376 194092 321652 194120
rect 217376 194080 217382 194092
rect 321646 194080 321652 194092
rect 321704 194080 321710 194132
rect 126238 194012 126244 194064
rect 126296 194052 126302 194064
rect 240962 194052 240968 194064
rect 126296 194024 240968 194052
rect 126296 194012 126302 194024
rect 240962 194012 240968 194024
rect 241020 194012 241026 194064
rect 100754 193944 100760 193996
rect 100812 193984 100818 193996
rect 252646 193984 252652 193996
rect 100812 193956 252652 193984
rect 100812 193944 100818 193956
rect 252646 193944 252652 193956
rect 252704 193944 252710 193996
rect 142798 193876 142804 193928
rect 142856 193916 142862 193928
rect 354766 193916 354772 193928
rect 142856 193888 354772 193916
rect 142856 193876 142862 193888
rect 354766 193876 354772 193888
rect 354824 193876 354830 193928
rect 152642 193808 152648 193860
rect 152700 193848 152706 193860
rect 410610 193848 410616 193860
rect 152700 193820 410616 193848
rect 152700 193808 152706 193820
rect 410610 193808 410616 193820
rect 410668 193808 410674 193860
rect 151262 192788 151268 192840
rect 151320 192828 151326 192840
rect 242250 192828 242256 192840
rect 151320 192800 242256 192828
rect 151320 192788 151326 192800
rect 242250 192788 242256 192800
rect 242308 192788 242314 192840
rect 141418 192720 141424 192772
rect 141476 192760 141482 192772
rect 211798 192760 211804 192772
rect 141476 192732 211804 192760
rect 141476 192720 141482 192732
rect 211798 192720 211804 192732
rect 211856 192720 211862 192772
rect 225598 192720 225604 192772
rect 225656 192760 225662 192772
rect 328730 192760 328736 192772
rect 225656 192732 328736 192760
rect 225656 192720 225662 192732
rect 328730 192720 328736 192732
rect 328788 192720 328794 192772
rect 92474 192652 92480 192704
rect 92532 192692 92538 192704
rect 256970 192692 256976 192704
rect 92532 192664 256976 192692
rect 92532 192652 92538 192664
rect 256970 192652 256976 192664
rect 257028 192652 257034 192704
rect 175090 192584 175096 192636
rect 175148 192624 175154 192636
rect 343818 192624 343824 192636
rect 175148 192596 343824 192624
rect 175148 192584 175154 192596
rect 343818 192584 343824 192596
rect 343876 192584 343882 192636
rect 70394 192516 70400 192568
rect 70452 192556 70458 192568
rect 254210 192556 254216 192568
rect 70452 192528 254216 192556
rect 70452 192516 70458 192528
rect 254210 192516 254216 192528
rect 254268 192516 254274 192568
rect 165522 192448 165528 192500
rect 165580 192488 165586 192500
rect 411898 192488 411904 192500
rect 165580 192460 411904 192488
rect 165580 192448 165586 192460
rect 411898 192448 411904 192460
rect 411956 192448 411962 192500
rect 249058 191292 249064 191344
rect 249116 191332 249122 191344
rect 271874 191332 271880 191344
rect 249116 191304 271880 191332
rect 249116 191292 249122 191304
rect 271874 191292 271880 191304
rect 271932 191292 271938 191344
rect 202230 191224 202236 191276
rect 202288 191264 202294 191276
rect 335538 191264 335544 191276
rect 202288 191236 335544 191264
rect 202288 191224 202294 191236
rect 335538 191224 335544 191236
rect 335596 191224 335602 191276
rect 69106 191156 69112 191208
rect 69164 191196 69170 191208
rect 251266 191196 251272 191208
rect 69164 191168 251272 191196
rect 69164 191156 69170 191168
rect 251266 191156 251272 191168
rect 251324 191156 251330 191208
rect 273990 191156 273996 191208
rect 274048 191196 274054 191208
rect 331398 191196 331404 191208
rect 274048 191168 331404 191196
rect 274048 191156 274054 191168
rect 331398 191156 331404 191168
rect 331456 191156 331462 191208
rect 118602 191088 118608 191140
rect 118660 191128 118666 191140
rect 503898 191128 503904 191140
rect 118660 191100 503904 191128
rect 118660 191088 118666 191100
rect 503898 191088 503904 191100
rect 503956 191088 503962 191140
rect 153930 190068 153936 190120
rect 153988 190108 153994 190120
rect 195330 190108 195336 190120
rect 153988 190080 195336 190108
rect 153988 190068 153994 190080
rect 195330 190068 195336 190080
rect 195388 190068 195394 190120
rect 192570 190000 192576 190052
rect 192628 190040 192634 190052
rect 243538 190040 243544 190052
rect 192628 190012 243544 190040
rect 192628 190000 192634 190012
rect 243538 190000 243544 190012
rect 243596 190000 243602 190052
rect 169018 189932 169024 189984
rect 169076 189972 169082 189984
rect 264974 189972 264980 189984
rect 169076 189944 264980 189972
rect 169076 189932 169082 189944
rect 264974 189932 264980 189944
rect 265032 189932 265038 189984
rect 135990 189864 135996 189916
rect 136048 189904 136054 189916
rect 197998 189904 198004 189916
rect 136048 189876 198004 189904
rect 136048 189864 136054 189876
rect 197998 189864 198004 189876
rect 198056 189864 198062 189916
rect 221458 189864 221464 189916
rect 221516 189904 221522 189916
rect 335630 189904 335636 189916
rect 221516 189876 335636 189904
rect 221516 189864 221522 189876
rect 335630 189864 335636 189876
rect 335688 189864 335694 189916
rect 138750 189796 138756 189848
rect 138808 189836 138814 189848
rect 256786 189836 256792 189848
rect 138808 189808 256792 189836
rect 138808 189796 138814 189808
rect 256786 189796 256792 189808
rect 256844 189796 256850 189848
rect 181530 189728 181536 189780
rect 181588 189768 181594 189780
rect 345198 189768 345204 189780
rect 181588 189740 345204 189768
rect 181588 189728 181594 189740
rect 345198 189728 345204 189740
rect 345256 189728 345262 189780
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 53098 189020 53104 189032
rect 3476 188992 53104 189020
rect 3476 188980 3482 188992
rect 53098 188980 53104 188992
rect 53156 188980 53162 189032
rect 155218 188572 155224 188624
rect 155276 188612 155282 188624
rect 204990 188612 204996 188624
rect 155276 188584 204996 188612
rect 155276 188572 155282 188584
rect 204990 188572 204996 188584
rect 205048 188572 205054 188624
rect 220078 188572 220084 188624
rect 220136 188612 220142 188624
rect 273346 188612 273352 188624
rect 220136 188584 273352 188612
rect 220136 188572 220142 188584
rect 273346 188572 273352 188584
rect 273404 188572 273410 188624
rect 124858 188504 124864 188556
rect 124916 188544 124922 188556
rect 271966 188544 271972 188556
rect 124916 188516 271972 188544
rect 124916 188504 124922 188516
rect 271966 188504 271972 188516
rect 272024 188504 272030 188556
rect 84194 188436 84200 188488
rect 84252 188476 84258 188488
rect 250070 188476 250076 188488
rect 84252 188448 250076 188476
rect 84252 188436 84258 188448
rect 250070 188436 250076 188448
rect 250128 188436 250134 188488
rect 114462 188368 114468 188420
rect 114520 188408 114526 188420
rect 334066 188408 334072 188420
rect 114520 188380 334072 188408
rect 114520 188368 114526 188380
rect 334066 188368 334072 188380
rect 334124 188368 334130 188420
rect 57790 188300 57796 188352
rect 57848 188340 57854 188352
rect 259546 188340 259552 188352
rect 57848 188312 259552 188340
rect 57848 188300 57854 188312
rect 259546 188300 259552 188312
rect 259604 188300 259610 188352
rect 265618 188300 265624 188352
rect 265676 188340 265682 188352
rect 494330 188340 494336 188352
rect 265676 188312 494336 188340
rect 265676 188300 265682 188312
rect 494330 188300 494336 188312
rect 494388 188300 494394 188352
rect 137370 187144 137376 187196
rect 137428 187184 137434 187196
rect 255406 187184 255412 187196
rect 137428 187156 255412 187184
rect 137428 187144 137434 187156
rect 255406 187144 255412 187156
rect 255464 187144 255470 187196
rect 110414 187076 110420 187128
rect 110472 187116 110478 187128
rect 249886 187116 249892 187128
rect 110472 187088 249892 187116
rect 110472 187076 110478 187088
rect 249886 187076 249892 187088
rect 249944 187076 249950 187128
rect 146938 187008 146944 187060
rect 146996 187048 147002 187060
rect 352098 187048 352104 187060
rect 146996 187020 352104 187048
rect 146996 187008 147002 187020
rect 352098 187008 352104 187020
rect 352156 187008 352162 187060
rect 50890 186940 50896 186992
rect 50948 186980 50954 186992
rect 266354 186980 266360 186992
rect 50948 186952 266360 186980
rect 50948 186940 50954 186952
rect 266354 186940 266360 186952
rect 266412 186940 266418 186992
rect 228358 185920 228364 185972
rect 228416 185960 228422 185972
rect 262398 185960 262404 185972
rect 228416 185932 262404 185960
rect 228416 185920 228422 185932
rect 262398 185920 262404 185932
rect 262456 185920 262462 185972
rect 134518 185852 134524 185904
rect 134576 185892 134582 185904
rect 213178 185892 213184 185904
rect 134576 185864 213184 185892
rect 134576 185852 134582 185864
rect 213178 185852 213184 185864
rect 213236 185852 213242 185904
rect 229738 185852 229744 185904
rect 229796 185892 229802 185904
rect 342438 185892 342444 185904
rect 229796 185864 342444 185892
rect 229796 185852 229802 185864
rect 342438 185852 342444 185864
rect 342496 185852 342502 185904
rect 122098 185784 122104 185836
rect 122156 185824 122162 185836
rect 249058 185824 249064 185836
rect 122156 185796 249064 185824
rect 122156 185784 122162 185796
rect 249058 185784 249064 185796
rect 249116 185784 249122 185836
rect 131758 185716 131764 185768
rect 131816 185756 131822 185768
rect 263778 185756 263784 185768
rect 131816 185728 263784 185756
rect 131816 185716 131822 185728
rect 263778 185716 263784 185728
rect 263836 185716 263842 185768
rect 191190 185648 191196 185700
rect 191248 185688 191254 185700
rect 339586 185688 339592 185700
rect 191248 185660 339592 185688
rect 191248 185648 191254 185660
rect 339586 185648 339592 185660
rect 339644 185648 339650 185700
rect 393958 185648 393964 185700
rect 394016 185688 394022 185700
rect 425330 185688 425336 185700
rect 394016 185660 425336 185688
rect 394016 185648 394022 185660
rect 425330 185648 425336 185660
rect 425388 185648 425394 185700
rect 125042 185580 125048 185632
rect 125100 185620 125106 185632
rect 258350 185620 258356 185632
rect 125100 185592 258356 185620
rect 125100 185580 125106 185592
rect 258350 185580 258356 185592
rect 258408 185580 258414 185632
rect 290458 185580 290464 185632
rect 290516 185620 290522 185632
rect 498470 185620 498476 185632
rect 290516 185592 498476 185620
rect 290516 185580 290522 185592
rect 498470 185580 498476 185592
rect 498528 185580 498534 185632
rect 102042 184900 102048 184952
rect 102100 184940 102106 184952
rect 205082 184940 205088 184952
rect 102100 184912 205088 184940
rect 102100 184900 102106 184912
rect 205082 184900 205088 184912
rect 205140 184900 205146 184952
rect 244918 184356 244924 184408
rect 244976 184396 244982 184408
rect 290458 184396 290464 184408
rect 244976 184368 290464 184396
rect 244976 184356 244982 184368
rect 290458 184356 290464 184368
rect 290516 184356 290522 184408
rect 485038 184356 485044 184408
rect 485096 184396 485102 184408
rect 501138 184396 501144 184408
rect 485096 184368 501144 184396
rect 485096 184356 485102 184368
rect 501138 184356 501144 184368
rect 501196 184356 501202 184408
rect 173250 184288 173256 184340
rect 173308 184328 173314 184340
rect 251358 184328 251364 184340
rect 173308 184300 251364 184328
rect 173308 184288 173314 184300
rect 251358 184288 251364 184300
rect 251416 184288 251422 184340
rect 251818 184288 251824 184340
rect 251876 184328 251882 184340
rect 340966 184328 340972 184340
rect 251876 184300 340972 184328
rect 251876 184288 251882 184300
rect 340966 184288 340972 184300
rect 341024 184288 341030 184340
rect 471238 184288 471244 184340
rect 471296 184328 471302 184340
rect 488626 184328 488632 184340
rect 471296 184300 488632 184328
rect 471296 184288 471302 184300
rect 488626 184288 488632 184300
rect 488684 184288 488690 184340
rect 152458 184220 152464 184272
rect 152516 184260 152522 184272
rect 202230 184260 202236 184272
rect 152516 184232 202236 184260
rect 152516 184220 152522 184232
rect 202230 184220 202236 184232
rect 202288 184220 202294 184272
rect 214558 184220 214564 184272
rect 214616 184260 214622 184272
rect 330110 184260 330116 184272
rect 214616 184232 330116 184260
rect 214616 184220 214622 184232
rect 330110 184220 330116 184232
rect 330168 184220 330174 184272
rect 457438 184220 457444 184272
rect 457496 184260 457502 184272
rect 510798 184260 510804 184272
rect 457496 184232 510804 184260
rect 457496 184220 457502 184232
rect 510798 184220 510804 184232
rect 510856 184220 510862 184272
rect 160830 184152 160836 184204
rect 160888 184192 160894 184204
rect 506658 184192 506664 184204
rect 160888 184164 506664 184192
rect 160888 184152 160894 184164
rect 506658 184152 506664 184164
rect 506716 184152 506722 184204
rect 107562 183608 107568 183660
rect 107620 183648 107626 183660
rect 173158 183648 173164 183660
rect 107620 183620 173164 183648
rect 107620 183608 107626 183620
rect 173158 183608 173164 183620
rect 173216 183608 173222 183660
rect 125502 183540 125508 183592
rect 125560 183580 125566 183592
rect 214650 183580 214656 183592
rect 125560 183552 214656 183580
rect 125560 183540 125566 183552
rect 214650 183540 214656 183552
rect 214708 183540 214714 183592
rect 169110 183132 169116 183184
rect 169168 183172 169174 183184
rect 260926 183172 260932 183184
rect 169168 183144 260932 183172
rect 169168 183132 169174 183144
rect 260926 183132 260932 183144
rect 260984 183132 260990 183184
rect 160738 183064 160744 183116
rect 160796 183104 160802 183116
rect 215938 183104 215944 183116
rect 160796 183076 215944 183104
rect 160796 183064 160802 183076
rect 215938 183064 215944 183076
rect 215996 183064 216002 183116
rect 242158 183064 242164 183116
rect 242216 183104 242222 183116
rect 341058 183104 341064 183116
rect 242216 183076 341064 183104
rect 242216 183064 242222 183076
rect 341058 183064 341064 183076
rect 341116 183064 341122 183116
rect 133322 182996 133328 183048
rect 133380 183036 133386 183048
rect 248046 183036 248052 183048
rect 133380 183008 248052 183036
rect 133380 182996 133386 183008
rect 248046 182996 248052 183008
rect 248104 182996 248110 183048
rect 202782 182928 202788 182980
rect 202840 182968 202846 182980
rect 352190 182968 352196 182980
rect 202840 182940 352196 182968
rect 202840 182928 202846 182940
rect 352190 182928 352196 182940
rect 352248 182928 352254 182980
rect 184842 182860 184848 182912
rect 184900 182900 184906 182912
rect 345290 182900 345296 182912
rect 184900 182872 345296 182900
rect 184900 182860 184906 182872
rect 345290 182860 345296 182872
rect 345348 182860 345354 182912
rect 414658 182860 414664 182912
rect 414716 182900 414722 182912
rect 505094 182900 505100 182912
rect 414716 182872 505100 182900
rect 414716 182860 414722 182872
rect 505094 182860 505100 182872
rect 505152 182860 505158 182912
rect 22738 182792 22744 182844
rect 22796 182832 22802 182844
rect 109034 182832 109040 182844
rect 22796 182804 109040 182832
rect 22796 182792 22802 182804
rect 109034 182792 109040 182804
rect 109092 182792 109098 182844
rect 178770 182792 178776 182844
rect 178828 182832 178834 182844
rect 343910 182832 343916 182844
rect 178828 182804 343916 182832
rect 178828 182792 178834 182804
rect 343910 182792 343916 182804
rect 343968 182792 343974 182844
rect 419258 182792 419264 182844
rect 419316 182832 419322 182844
rect 580258 182832 580264 182844
rect 419316 182804 580264 182832
rect 419316 182792 419322 182804
rect 580258 182792 580264 182804
rect 580316 182792 580322 182844
rect 132402 182384 132408 182436
rect 132460 182424 132466 182436
rect 164878 182424 164884 182436
rect 132460 182396 164884 182424
rect 132460 182384 132466 182396
rect 164878 182384 164884 182396
rect 164936 182384 164942 182436
rect 110690 182316 110696 182368
rect 110748 182356 110754 182368
rect 170490 182356 170496 182368
rect 110748 182328 170496 182356
rect 110748 182316 110754 182328
rect 170490 182316 170496 182328
rect 170548 182316 170554 182368
rect 112438 182248 112444 182300
rect 112496 182288 112502 182300
rect 171962 182288 171968 182300
rect 112496 182260 171968 182288
rect 112496 182248 112502 182260
rect 171962 182248 171968 182260
rect 172020 182248 172026 182300
rect 119522 182180 119528 182232
rect 119580 182220 119586 182232
rect 196802 182220 196808 182232
rect 119580 182192 196808 182220
rect 119580 182180 119586 182192
rect 196802 182180 196808 182192
rect 196860 182180 196866 182232
rect 489178 182180 489184 182232
rect 489236 182220 489242 182232
rect 490558 182220 490564 182232
rect 489236 182192 490564 182220
rect 489236 182180 489242 182192
rect 490558 182180 490564 182192
rect 490616 182180 490622 182232
rect 454678 182112 454684 182164
rect 454736 182152 454742 182164
rect 455598 182152 455604 182164
rect 454736 182124 455604 182152
rect 454736 182112 454742 182124
rect 455598 182112 455604 182124
rect 455656 182112 455662 182164
rect 461578 182112 461584 182164
rect 461636 182152 461642 182164
rect 462590 182152 462596 182164
rect 461636 182124 462596 182152
rect 461636 182112 461642 182124
rect 462590 182112 462596 182124
rect 462648 182112 462654 182164
rect 475470 182112 475476 182164
rect 475528 182152 475534 182164
rect 476574 182152 476580 182164
rect 475528 182124 476580 182152
rect 475528 182112 475534 182124
rect 476574 182112 476580 182124
rect 476632 182112 476638 182164
rect 485130 182112 485136 182164
rect 485188 182152 485194 182164
rect 485774 182152 485780 182164
rect 485188 182124 485780 182152
rect 485188 182112 485194 182124
rect 485774 182112 485780 182124
rect 485832 182112 485838 182164
rect 242250 181704 242256 181756
rect 242308 181744 242314 181756
rect 260834 181744 260840 181756
rect 242308 181716 260840 181744
rect 242308 181704 242314 181716
rect 260834 181704 260840 181716
rect 260892 181704 260898 181756
rect 486418 181704 486424 181756
rect 486476 181744 486482 181756
rect 492858 181744 492864 181756
rect 486476 181716 492864 181744
rect 486476 181704 486482 181716
rect 492858 181704 492864 181716
rect 492916 181704 492922 181756
rect 240962 181636 240968 181688
rect 241020 181676 241026 181688
rect 262306 181676 262312 181688
rect 241020 181648 262312 181676
rect 241020 181636 241026 181648
rect 262306 181636 262312 181648
rect 262364 181636 262370 181688
rect 410518 181636 410524 181688
rect 410576 181676 410582 181688
rect 444006 181676 444012 181688
rect 410576 181648 444012 181676
rect 410576 181636 410582 181648
rect 444006 181636 444012 181648
rect 444064 181636 444070 181688
rect 446490 181636 446496 181688
rect 446548 181676 446554 181688
rect 460198 181676 460204 181688
rect 446548 181648 460204 181676
rect 446548 181636 446554 181648
rect 460198 181636 460204 181648
rect 460256 181636 460262 181688
rect 464338 181636 464344 181688
rect 464396 181676 464402 181688
rect 474182 181676 474188 181688
rect 464396 181648 474188 181676
rect 464396 181636 464402 181648
rect 474182 181636 474188 181648
rect 474240 181636 474246 181688
rect 482278 181636 482284 181688
rect 482336 181676 482342 181688
rect 502518 181676 502524 181688
rect 482336 181648 502524 181676
rect 482336 181636 482342 181648
rect 502518 181636 502524 181648
rect 502576 181636 502582 181688
rect 159358 181568 159364 181620
rect 159416 181608 159422 181620
rect 198090 181608 198096 181620
rect 159416 181580 198096 181608
rect 159416 181568 159422 181580
rect 198090 181568 198096 181580
rect 198148 181568 198154 181620
rect 222838 181568 222844 181620
rect 222896 181608 222902 181620
rect 269206 181608 269212 181620
rect 222896 181580 269212 181608
rect 222896 181568 222902 181580
rect 269206 181568 269212 181580
rect 269264 181568 269270 181620
rect 284938 181568 284944 181620
rect 284996 181608 285002 181620
rect 338206 181608 338212 181620
rect 284996 181580 338212 181608
rect 284996 181568 285002 181580
rect 338206 181568 338212 181580
rect 338264 181568 338270 181620
rect 403618 181568 403624 181620
rect 403676 181608 403682 181620
rect 441614 181608 441620 181620
rect 403676 181580 441620 181608
rect 403676 181568 403682 181580
rect 441614 181568 441620 181580
rect 441672 181568 441678 181620
rect 443638 181568 443644 181620
rect 443696 181608 443702 181620
rect 505278 181608 505284 181620
rect 443696 181580 505284 181608
rect 443696 181568 443702 181580
rect 505278 181568 505284 181580
rect 505336 181568 505342 181620
rect 166350 181500 166356 181552
rect 166408 181540 166414 181552
rect 209038 181540 209044 181552
rect 166408 181512 209044 181540
rect 166408 181500 166414 181512
rect 209038 181500 209044 181512
rect 209096 181500 209102 181552
rect 232682 181500 232688 181552
rect 232740 181540 232746 181552
rect 259638 181540 259644 181552
rect 232740 181512 259644 181540
rect 232740 181500 232746 181512
rect 259638 181500 259644 181512
rect 259696 181500 259702 181552
rect 262858 181500 262864 181552
rect 262916 181540 262922 181552
rect 446398 181540 446404 181552
rect 262916 181512 446404 181540
rect 262916 181500 262922 181512
rect 446398 181500 446404 181512
rect 446456 181500 446462 181552
rect 447778 181500 447784 181552
rect 447836 181540 447842 181552
rect 507946 181540 507952 181552
rect 447836 181512 507952 181540
rect 447836 181500 447842 181512
rect 507946 181500 507952 181512
rect 508004 181500 508010 181552
rect 196710 181432 196716 181484
rect 196768 181472 196774 181484
rect 451366 181472 451372 181484
rect 196768 181444 451372 181472
rect 196768 181432 196774 181444
rect 451366 181432 451372 181444
rect 451424 181432 451430 181484
rect 468478 181432 468484 181484
rect 468536 181472 468542 181484
rect 501230 181472 501236 181484
rect 468536 181444 501236 181472
rect 468536 181432 468542 181444
rect 501230 181432 501236 181444
rect 501288 181432 501294 181484
rect 129458 180956 129464 181008
rect 129516 180996 129522 181008
rect 166534 180996 166540 181008
rect 129516 180968 166540 180996
rect 129516 180956 129522 180968
rect 166534 180956 166540 180968
rect 166592 180956 166598 181008
rect 124030 180888 124036 180940
rect 124088 180928 124094 180940
rect 167914 180928 167920 180940
rect 124088 180900 167920 180928
rect 124088 180888 124094 180900
rect 167914 180888 167920 180900
rect 167972 180888 167978 180940
rect 118418 180820 118424 180872
rect 118476 180860 118482 180872
rect 169202 180860 169208 180872
rect 118476 180832 169208 180860
rect 118476 180820 118482 180832
rect 169202 180820 169208 180832
rect 169260 180820 169266 180872
rect 238110 180344 238116 180396
rect 238168 180384 238174 180396
rect 261018 180384 261024 180396
rect 238168 180356 261024 180384
rect 238168 180344 238174 180356
rect 261018 180344 261024 180356
rect 261076 180344 261082 180396
rect 222930 180276 222936 180328
rect 222988 180316 222994 180328
rect 249334 180316 249340 180328
rect 222988 180288 249340 180316
rect 222988 180276 222994 180288
rect 249334 180276 249340 180288
rect 249392 180276 249398 180328
rect 165430 180208 165436 180260
rect 165488 180248 165494 180260
rect 239030 180248 239036 180260
rect 165488 180220 239036 180248
rect 165488 180208 165494 180220
rect 239030 180208 239036 180220
rect 239088 180208 239094 180260
rect 309870 180208 309876 180260
rect 309928 180248 309934 180260
rect 325878 180248 325884 180260
rect 309928 180220 325884 180248
rect 309928 180208 309934 180220
rect 325878 180208 325884 180220
rect 325936 180208 325942 180260
rect 167822 180140 167828 180192
rect 167880 180180 167886 180192
rect 335446 180180 335452 180192
rect 167880 180152 335452 180180
rect 167880 180140 167886 180152
rect 335446 180140 335452 180152
rect 335504 180140 335510 180192
rect 493318 180140 493324 180192
rect 493376 180180 493382 180192
rect 512086 180180 512092 180192
rect 493376 180152 512092 180180
rect 493376 180140 493382 180152
rect 512086 180140 512092 180152
rect 512144 180140 512150 180192
rect 156598 180072 156604 180124
rect 156656 180112 156662 180124
rect 210418 180112 210424 180124
rect 156656 180084 210424 180112
rect 156656 180072 156662 180084
rect 210418 180072 210424 180084
rect 210476 180072 210482 180124
rect 216122 180072 216128 180124
rect 216180 180112 216186 180124
rect 509234 180112 509240 180124
rect 216180 180084 509240 180112
rect 216180 180072 216186 180084
rect 509234 180072 509240 180084
rect 509292 180072 509298 180124
rect 385678 180004 385684 180056
rect 385736 180044 385742 180056
rect 386322 180044 386328 180056
rect 385736 180016 386328 180044
rect 385736 180004 385742 180016
rect 386322 180004 386328 180016
rect 386380 180004 386386 180056
rect 490650 179868 490656 179920
rect 490708 179908 490714 179920
rect 495526 179908 495532 179920
rect 490708 179880 495532 179908
rect 490708 179868 490714 179880
rect 495526 179868 495532 179880
rect 495584 179868 495590 179920
rect 134702 179596 134708 179648
rect 134760 179636 134766 179648
rect 165430 179636 165436 179648
rect 134760 179608 165436 179636
rect 134760 179596 134766 179608
rect 165430 179596 165436 179608
rect 165488 179596 165494 179648
rect 126606 179528 126612 179580
rect 126664 179568 126670 179580
rect 170674 179568 170680 179580
rect 126664 179540 170680 179568
rect 126664 179528 126670 179540
rect 170674 179528 170680 179540
rect 170732 179528 170738 179580
rect 115842 179460 115848 179512
rect 115900 179500 115906 179512
rect 166258 179500 166264 179512
rect 115900 179472 166264 179500
rect 115900 179460 115906 179472
rect 166258 179460 166264 179472
rect 166316 179460 166322 179512
rect 414658 179460 414664 179512
rect 414716 179500 414722 179512
rect 492582 179500 492588 179512
rect 414716 179472 492588 179500
rect 414716 179460 414722 179472
rect 492582 179460 492588 179472
rect 492640 179460 492646 179512
rect 97810 179392 97816 179444
rect 97868 179432 97874 179444
rect 171870 179432 171876 179444
rect 97868 179404 171876 179432
rect 97868 179392 97874 179404
rect 171870 179392 171876 179404
rect 171928 179392 171934 179444
rect 386322 179392 386328 179444
rect 386380 179432 386386 179444
rect 580258 179432 580264 179444
rect 386380 179404 580264 179432
rect 386380 179392 386386 179404
rect 580258 179392 580264 179404
rect 580316 179392 580322 179444
rect 236638 178984 236644 179036
rect 236696 179024 236702 179036
rect 255498 179024 255504 179036
rect 236696 178996 255504 179024
rect 236696 178984 236702 178996
rect 255498 178984 255504 178996
rect 255556 178984 255562 179036
rect 240778 178916 240784 178968
rect 240836 178956 240842 178968
rect 265066 178956 265072 178968
rect 240836 178928 265072 178956
rect 240836 178916 240842 178928
rect 265066 178916 265072 178928
rect 265124 178916 265130 178968
rect 231118 178848 231124 178900
rect 231176 178888 231182 178900
rect 274634 178888 274640 178900
rect 231176 178860 274640 178888
rect 231176 178848 231182 178860
rect 274634 178848 274640 178860
rect 274692 178848 274698 178900
rect 312538 178848 312544 178900
rect 312596 178888 312602 178900
rect 327258 178888 327264 178900
rect 312596 178860 327264 178888
rect 312596 178848 312602 178860
rect 327258 178848 327264 178860
rect 327316 178848 327322 178900
rect 180242 178780 180248 178832
rect 180300 178820 180306 178832
rect 247954 178820 247960 178832
rect 180300 178792 247960 178820
rect 180300 178780 180306 178792
rect 247954 178780 247960 178792
rect 248012 178780 248018 178832
rect 261478 178780 261484 178832
rect 261536 178820 261542 178832
rect 321278 178820 321284 178832
rect 261536 178792 321284 178820
rect 261536 178780 261542 178792
rect 321278 178780 321284 178792
rect 321336 178780 321342 178832
rect 246298 178712 246304 178764
rect 246356 178752 246362 178764
rect 349338 178752 349344 178764
rect 246356 178724 349344 178752
rect 246356 178712 246362 178724
rect 349338 178712 349344 178724
rect 349396 178712 349402 178764
rect 195882 178644 195888 178696
rect 195940 178684 195946 178696
rect 417510 178684 417516 178696
rect 195940 178656 417516 178684
rect 195940 178644 195946 178656
rect 417510 178644 417516 178656
rect 417568 178644 417574 178696
rect 502978 178644 502984 178696
rect 503036 178684 503042 178696
rect 580166 178684 580172 178696
rect 503036 178656 580172 178684
rect 503036 178644 503042 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 98730 178372 98736 178424
rect 98788 178412 98794 178424
rect 196710 178412 196716 178424
rect 98788 178384 196716 178412
rect 98788 178372 98794 178384
rect 196710 178372 196716 178384
rect 196768 178372 196774 178424
rect 148226 178304 148232 178356
rect 148284 178344 148290 178356
rect 170398 178344 170404 178356
rect 148284 178316 170404 178344
rect 148284 178304 148290 178316
rect 170398 178304 170404 178316
rect 170456 178304 170462 178356
rect 110322 178236 110328 178288
rect 110380 178276 110386 178288
rect 178770 178276 178776 178288
rect 110380 178248 178776 178276
rect 110380 178236 110386 178248
rect 178770 178236 178776 178248
rect 178828 178236 178834 178288
rect 113726 178168 113732 178220
rect 113784 178208 113790 178220
rect 196894 178208 196900 178220
rect 113784 178180 196900 178208
rect 113784 178168 113790 178180
rect 196894 178168 196900 178180
rect 196952 178168 196958 178220
rect 127066 178100 127072 178152
rect 127124 178140 127130 178152
rect 214558 178140 214564 178152
rect 127124 178112 214564 178140
rect 127124 178100 127130 178112
rect 214558 178100 214564 178112
rect 214616 178100 214622 178152
rect 159910 178032 159916 178084
rect 159968 178072 159974 178084
rect 169018 178072 169024 178084
rect 159968 178044 169024 178072
rect 159968 178032 159974 178044
rect 169018 178032 169024 178044
rect 169076 178032 169082 178084
rect 308398 178032 308404 178084
rect 308456 178072 308462 178084
rect 316034 178072 316040 178084
rect 308456 178044 316040 178072
rect 308456 178032 308462 178044
rect 316034 178032 316040 178044
rect 316092 178072 316098 178084
rect 316402 178072 316408 178084
rect 316092 178044 316408 178072
rect 316092 178032 316098 178044
rect 316402 178032 316408 178044
rect 316460 178032 316466 178084
rect 246390 177624 246396 177676
rect 246448 177664 246454 177676
rect 255590 177664 255596 177676
rect 246448 177636 255596 177664
rect 246448 177624 246454 177636
rect 255590 177624 255596 177636
rect 255648 177624 255654 177676
rect 314010 177624 314016 177676
rect 314068 177664 314074 177676
rect 332778 177664 332784 177676
rect 314068 177636 332784 177664
rect 314068 177624 314074 177636
rect 332778 177624 332784 177636
rect 332836 177624 332842 177676
rect 238018 177556 238024 177608
rect 238076 177596 238082 177608
rect 258258 177596 258264 177608
rect 238076 177568 258264 177596
rect 238076 177556 238082 177568
rect 258258 177556 258264 177568
rect 258316 177556 258322 177608
rect 312630 177556 312636 177608
rect 312688 177596 312694 177608
rect 339494 177596 339500 177608
rect 312688 177568 339500 177596
rect 312688 177556 312694 177568
rect 339494 177556 339500 177568
rect 339552 177556 339558 177608
rect 174538 177488 174544 177540
rect 174596 177528 174602 177540
rect 258074 177528 258080 177540
rect 174596 177500 258080 177528
rect 174596 177488 174602 177500
rect 258074 177488 258080 177500
rect 258132 177488 258138 177540
rect 307110 177488 307116 177540
rect 307168 177528 307174 177540
rect 334158 177528 334164 177540
rect 307168 177500 334164 177528
rect 307168 177488 307174 177500
rect 334158 177488 334164 177500
rect 334216 177488 334222 177540
rect 239030 177420 239036 177472
rect 239088 177460 239094 177472
rect 334250 177460 334256 177472
rect 239088 177432 334256 177460
rect 239088 177420 239094 177432
rect 334250 177420 334256 177432
rect 334308 177420 334314 177472
rect 209130 177352 209136 177404
rect 209188 177392 209194 177404
rect 332594 177392 332600 177404
rect 209188 177364 332600 177392
rect 209188 177352 209194 177364
rect 332594 177352 332600 177364
rect 332652 177352 332658 177404
rect 198642 177284 198648 177336
rect 198700 177324 198706 177336
rect 323118 177324 323124 177336
rect 198700 177296 323124 177324
rect 198700 177284 198706 177296
rect 323118 177284 323124 177296
rect 323176 177284 323182 177336
rect 133138 177012 133144 177064
rect 133196 177052 133202 177064
rect 165522 177052 165528 177064
rect 133196 177024 165528 177052
rect 133196 177012 133202 177024
rect 165522 177012 165528 177024
rect 165580 177012 165586 177064
rect 108114 176944 108120 176996
rect 108172 176984 108178 176996
rect 169110 176984 169116 176996
rect 108172 176956 169116 176984
rect 108172 176944 108178 176956
rect 169110 176944 169116 176956
rect 169168 176944 169174 176996
rect 103330 176876 103336 176928
rect 103388 176916 103394 176928
rect 167546 176916 167552 176928
rect 103388 176888 167552 176916
rect 103388 176876 103394 176888
rect 167546 176876 167552 176888
rect 167604 176876 167610 176928
rect 136082 176808 136088 176860
rect 136140 176848 136146 176860
rect 202782 176848 202788 176860
rect 136140 176820 202788 176848
rect 136140 176808 136146 176820
rect 202782 176808 202788 176820
rect 202840 176808 202846 176860
rect 104618 176740 104624 176792
rect 104676 176780 104682 176792
rect 174630 176780 174636 176792
rect 104676 176752 174636 176780
rect 104676 176740 104682 176752
rect 174630 176740 174636 176752
rect 174688 176740 174694 176792
rect 128170 176672 128176 176724
rect 128228 176712 128234 176724
rect 214190 176712 214196 176724
rect 128228 176684 214196 176712
rect 128228 176672 128234 176684
rect 214190 176672 214196 176684
rect 214248 176672 214254 176724
rect 340138 176672 340144 176724
rect 340196 176712 340202 176724
rect 416774 176712 416780 176724
rect 340196 176684 416780 176712
rect 340196 176672 340202 176684
rect 416774 176672 416780 176684
rect 416832 176672 416838 176724
rect 202782 176604 202788 176656
rect 202840 176644 202846 176656
rect 213914 176644 213920 176656
rect 202840 176616 213920 176644
rect 202840 176604 202846 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 243538 176604 243544 176656
rect 243596 176644 243602 176656
rect 249242 176644 249248 176656
rect 243596 176616 249248 176644
rect 243596 176604 243602 176616
rect 249242 176604 249248 176616
rect 249300 176604 249306 176656
rect 319530 176604 319536 176656
rect 319588 176644 319594 176656
rect 327074 176644 327080 176656
rect 319588 176616 327080 176644
rect 319588 176604 319594 176616
rect 327074 176604 327080 176616
rect 327132 176604 327138 176656
rect 163498 176264 163504 176316
rect 163556 176304 163562 176316
rect 206370 176304 206376 176316
rect 163556 176276 206376 176304
rect 163556 176264 163562 176276
rect 206370 176264 206376 176276
rect 206428 176264 206434 176316
rect 120810 176196 120816 176248
rect 120868 176236 120874 176248
rect 166626 176236 166632 176248
rect 120868 176208 166632 176236
rect 120868 176196 120874 176208
rect 166626 176196 166632 176208
rect 166684 176196 166690 176248
rect 121914 176128 121920 176180
rect 121972 176168 121978 176180
rect 173250 176168 173256 176180
rect 121972 176140 173256 176168
rect 121972 176128 121978 176140
rect 173250 176128 173256 176140
rect 173308 176128 173314 176180
rect 102042 176060 102048 176112
rect 102100 176100 102106 176112
rect 167822 176100 167828 176112
rect 102100 176072 167828 176100
rect 102100 176060 102106 176072
rect 167822 176060 167828 176072
rect 167880 176060 167886 176112
rect 318150 176060 318156 176112
rect 318208 176100 318214 176112
rect 328638 176100 328644 176112
rect 318208 176072 328644 176100
rect 318208 176060 318214 176072
rect 328638 176060 328644 176072
rect 328696 176060 328702 176112
rect 130746 175992 130752 176044
rect 130804 176032 130810 176044
rect 214098 176032 214104 176044
rect 130804 176004 214104 176032
rect 130804 175992 130810 176004
rect 214098 175992 214104 176004
rect 214156 175992 214162 176044
rect 245102 175992 245108 176044
rect 245160 176032 245166 176044
rect 261110 176032 261116 176044
rect 245160 176004 261116 176032
rect 245160 175992 245166 176004
rect 261110 175992 261116 176004
rect 261168 175992 261174 176044
rect 318058 175992 318064 176044
rect 318116 176032 318122 176044
rect 331490 176032 331496 176044
rect 318116 176004 331496 176032
rect 318116 175992 318122 176004
rect 331490 175992 331496 176004
rect 331548 175992 331554 176044
rect 116946 175924 116952 175976
rect 117004 175964 117010 175976
rect 166350 175964 166356 175976
rect 117004 175936 166356 175964
rect 117004 175924 117010 175936
rect 166350 175924 166356 175936
rect 166408 175924 166414 175976
rect 166442 175924 166448 175976
rect 166500 175964 166506 175976
rect 251450 175964 251456 175976
rect 166500 175936 251456 175964
rect 166500 175924 166506 175936
rect 251450 175924 251456 175936
rect 251508 175924 251514 175976
rect 269758 175924 269764 175976
rect 269816 175964 269822 175976
rect 324406 175964 324412 175976
rect 269816 175936 324412 175964
rect 269816 175924 269822 175936
rect 324406 175924 324412 175936
rect 324464 175924 324470 175976
rect 495526 175924 495532 175976
rect 495584 175964 495590 175976
rect 502426 175964 502432 175976
rect 495584 175936 502432 175964
rect 495584 175924 495590 175936
rect 502426 175924 502432 175936
rect 502484 175924 502490 175976
rect 248046 175788 248052 175840
rect 248104 175828 248110 175840
rect 249150 175828 249156 175840
rect 248104 175800 249156 175828
rect 248104 175788 248110 175800
rect 249150 175788 249156 175800
rect 249208 175788 249214 175840
rect 165430 175176 165436 175228
rect 165488 175216 165494 175228
rect 213914 175216 213920 175228
rect 165488 175188 213920 175216
rect 165488 175176 165494 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165522 175108 165528 175160
rect 165580 175148 165586 175160
rect 214006 175148 214012 175160
rect 165580 175120 214012 175148
rect 165580 175108 165586 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 338758 174496 338764 174548
rect 338816 174536 338822 174548
rect 348418 174536 348424 174548
rect 338816 174508 348424 174536
rect 338816 174496 338822 174508
rect 348418 174496 348424 174508
rect 348476 174496 348482 174548
rect 296254 174020 296260 174072
rect 296312 174060 296318 174072
rect 307662 174060 307668 174072
rect 296312 174032 307668 174060
rect 296312 174020 296318 174032
rect 307662 174020 307668 174032
rect 307720 174020 307726 174072
rect 285214 173952 285220 174004
rect 285272 173992 285278 174004
rect 307570 173992 307576 174004
rect 285272 173964 307576 173992
rect 285272 173952 285278 173964
rect 307570 173952 307576 173964
rect 307628 173952 307634 174004
rect 265802 173884 265808 173936
rect 265860 173924 265866 173936
rect 307110 173924 307116 173936
rect 265860 173896 307116 173924
rect 265860 173884 265866 173896
rect 307110 173884 307116 173896
rect 307168 173884 307174 173936
rect 358078 173884 358084 173936
rect 358136 173924 358142 173936
rect 416774 173924 416780 173936
rect 358136 173896 416780 173924
rect 358136 173884 358142 173896
rect 416774 173884 416780 173896
rect 416832 173884 416838 173936
rect 164878 173816 164884 173868
rect 164936 173856 164942 173868
rect 213914 173856 213920 173868
rect 164936 173828 213920 173856
rect 164936 173816 164942 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 252462 173816 252468 173868
rect 252520 173856 252526 173868
rect 263594 173856 263600 173868
rect 252520 173828 263600 173856
rect 252520 173816 252526 173828
rect 263594 173816 263600 173828
rect 263652 173816 263658 173868
rect 280798 172660 280804 172712
rect 280856 172700 280862 172712
rect 307570 172700 307576 172712
rect 280856 172672 307576 172700
rect 280856 172660 280862 172672
rect 307570 172660 307576 172672
rect 307628 172660 307634 172712
rect 263042 172592 263048 172644
rect 263100 172632 263106 172644
rect 307110 172632 307116 172644
rect 263100 172604 307116 172632
rect 263100 172592 263106 172604
rect 307110 172592 307116 172604
rect 307168 172592 307174 172644
rect 260374 172524 260380 172576
rect 260432 172564 260438 172576
rect 307662 172564 307668 172576
rect 260432 172536 307668 172564
rect 260432 172524 260438 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 496906 172524 496912 172576
rect 496964 172564 496970 172576
rect 501046 172564 501052 172576
rect 496964 172536 501052 172564
rect 496964 172524 496970 172536
rect 501046 172524 501052 172536
rect 501104 172524 501110 172576
rect 166534 172456 166540 172508
rect 166592 172496 166598 172508
rect 213914 172496 213920 172508
rect 166592 172468 213920 172496
rect 166592 172456 166598 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 252462 172456 252468 172508
rect 252520 172496 252526 172508
rect 260926 172496 260932 172508
rect 252520 172468 260932 172496
rect 252520 172456 252526 172468
rect 260926 172456 260932 172468
rect 260984 172456 260990 172508
rect 324314 172456 324320 172508
rect 324372 172496 324378 172508
rect 358814 172496 358820 172508
rect 324372 172468 358820 172496
rect 324372 172456 324378 172468
rect 358814 172456 358820 172468
rect 358872 172456 358878 172508
rect 252094 172388 252100 172440
rect 252152 172428 252158 172440
rect 255406 172428 255412 172440
rect 252152 172400 255412 172428
rect 252152 172388 252158 172400
rect 255406 172388 255412 172400
rect 255464 172388 255470 172440
rect 261662 171776 261668 171828
rect 261720 171816 261726 171828
rect 307294 171816 307300 171828
rect 261720 171788 307300 171816
rect 261720 171776 261726 171788
rect 307294 171776 307300 171788
rect 307352 171776 307358 171828
rect 252462 171504 252468 171556
rect 252520 171544 252526 171556
rect 258074 171544 258080 171556
rect 252520 171516 258080 171544
rect 252520 171504 252526 171516
rect 258074 171504 258080 171516
rect 258132 171504 258138 171556
rect 167638 171300 167644 171352
rect 167696 171340 167702 171352
rect 170582 171340 170588 171352
rect 167696 171312 170588 171340
rect 167696 171300 167702 171312
rect 170582 171300 170588 171312
rect 170640 171300 170646 171352
rect 283650 171164 283656 171216
rect 283708 171204 283714 171216
rect 306926 171204 306932 171216
rect 283708 171176 306932 171204
rect 283708 171164 283714 171176
rect 306926 171164 306932 171176
rect 306984 171164 306990 171216
rect 267182 171096 267188 171148
rect 267240 171136 267246 171148
rect 307662 171136 307668 171148
rect 267240 171108 307668 171136
rect 267240 171096 267246 171108
rect 307662 171096 307668 171108
rect 307720 171096 307726 171148
rect 170674 171028 170680 171080
rect 170732 171068 170738 171080
rect 213914 171068 213920 171080
rect 170732 171040 213920 171068
rect 170732 171028 170738 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 354674 171068 354680 171080
rect 324372 171040 354680 171068
rect 324372 171028 324378 171040
rect 354674 171028 354680 171040
rect 354732 171028 354738 171080
rect 252370 170552 252376 170604
rect 252428 170592 252434 170604
rect 256878 170592 256884 170604
rect 252428 170564 256884 170592
rect 252428 170552 252434 170564
rect 256878 170552 256884 170564
rect 256936 170552 256942 170604
rect 252462 170144 252468 170196
rect 252520 170184 252526 170196
rect 259638 170184 259644 170196
rect 252520 170156 259644 170184
rect 252520 170144 252526 170156
rect 259638 170144 259644 170156
rect 259696 170144 259702 170196
rect 285122 169872 285128 169924
rect 285180 169912 285186 169924
rect 307294 169912 307300 169924
rect 285180 169884 307300 169912
rect 285180 169872 285186 169884
rect 307294 169872 307300 169884
rect 307352 169872 307358 169924
rect 268470 169804 268476 169856
rect 268528 169844 268534 169856
rect 307662 169844 307668 169856
rect 268528 169816 307668 169844
rect 268528 169804 268534 169816
rect 307662 169804 307668 169816
rect 307720 169804 307726 169856
rect 260282 169736 260288 169788
rect 260340 169776 260346 169788
rect 307478 169776 307484 169788
rect 260340 169748 307484 169776
rect 260340 169736 260346 169748
rect 307478 169736 307484 169748
rect 307536 169736 307542 169788
rect 324958 169736 324964 169788
rect 325016 169776 325022 169788
rect 327074 169776 327080 169788
rect 325016 169748 327080 169776
rect 325016 169736 325022 169748
rect 327074 169736 327080 169748
rect 327132 169736 327138 169788
rect 167914 169668 167920 169720
rect 167972 169708 167978 169720
rect 213914 169708 213920 169720
rect 167972 169680 213920 169708
rect 167972 169668 167978 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 335630 169708 335636 169720
rect 324372 169680 335636 169708
rect 324372 169668 324378 169680
rect 335630 169668 335636 169680
rect 335688 169668 335694 169720
rect 324498 169600 324504 169652
rect 324556 169640 324562 169652
rect 332594 169640 332600 169652
rect 324556 169612 332600 169640
rect 324556 169600 324562 169612
rect 332594 169600 332600 169612
rect 332652 169600 332658 169652
rect 252370 169464 252376 169516
rect 252428 169504 252434 169516
rect 258166 169504 258172 169516
rect 252428 169476 258172 169504
rect 252428 169464 252434 169476
rect 258166 169464 258172 169476
rect 258224 169464 258230 169516
rect 252462 169124 252468 169176
rect 252520 169164 252526 169176
rect 259454 169164 259460 169176
rect 252520 169136 259460 169164
rect 252520 169124 252526 169136
rect 259454 169124 259460 169136
rect 259512 169124 259518 169176
rect 174630 168988 174636 169040
rect 174688 169028 174694 169040
rect 214466 169028 214472 169040
rect 174688 169000 214472 169028
rect 174688 168988 174694 169000
rect 214466 168988 214472 169000
rect 214524 168988 214530 169040
rect 297358 168988 297364 169040
rect 297416 169028 297422 169040
rect 306558 169028 306564 169040
rect 297416 169000 306564 169028
rect 297416 168988 297422 169000
rect 306558 168988 306564 169000
rect 306616 168988 306622 169040
rect 264422 168444 264428 168496
rect 264480 168484 264486 168496
rect 307110 168484 307116 168496
rect 264480 168456 307116 168484
rect 264480 168444 264486 168456
rect 307110 168444 307116 168456
rect 307168 168444 307174 168496
rect 264238 168376 264244 168428
rect 264296 168416 264302 168428
rect 307662 168416 307668 168428
rect 264296 168388 307668 168416
rect 264296 168376 264302 168388
rect 307662 168376 307668 168388
rect 307720 168376 307726 168428
rect 338758 168376 338764 168428
rect 338816 168416 338822 168428
rect 416774 168416 416780 168428
rect 338816 168388 416780 168416
rect 338816 168376 338822 168388
rect 416774 168376 416780 168388
rect 416832 168376 416838 168428
rect 166626 168308 166632 168360
rect 166684 168348 166690 168360
rect 214006 168348 214012 168360
rect 166684 168320 214012 168348
rect 166684 168308 166690 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 252462 168308 252468 168360
rect 252520 168348 252526 168360
rect 262214 168348 262220 168360
rect 252520 168320 262220 168348
rect 252520 168308 252526 168320
rect 262214 168308 262220 168320
rect 262272 168308 262278 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 347774 168348 347780 168360
rect 324372 168320 347780 168348
rect 324372 168308 324378 168320
rect 347774 168308 347780 168320
rect 347832 168308 347838 168360
rect 496906 168308 496912 168360
rect 496964 168348 496970 168360
rect 502334 168348 502340 168360
rect 496964 168320 502340 168348
rect 496964 168308 496970 168320
rect 502334 168308 502340 168320
rect 502392 168348 502398 168360
rect 503622 168348 503628 168360
rect 502392 168320 503628 168348
rect 502392 168308 502398 168320
rect 503622 168308 503628 168320
rect 503680 168308 503686 168360
rect 173250 168240 173256 168292
rect 173308 168280 173314 168292
rect 213914 168280 213920 168292
rect 173308 168252 213920 168280
rect 173308 168240 173314 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 324498 168240 324504 168292
rect 324556 168280 324562 168292
rect 345014 168280 345020 168292
rect 324556 168252 345020 168280
rect 324556 168240 324562 168252
rect 345014 168240 345020 168252
rect 345072 168240 345078 168292
rect 300210 167696 300216 167748
rect 300268 167736 300274 167748
rect 306742 167736 306748 167748
rect 300268 167708 306748 167736
rect 300268 167696 300274 167708
rect 306742 167696 306748 167708
rect 306800 167696 306806 167748
rect 259362 167628 259368 167680
rect 259420 167668 259426 167680
rect 307018 167668 307024 167680
rect 259420 167640 307024 167668
rect 259420 167628 259426 167640
rect 307018 167628 307024 167640
rect 307076 167628 307082 167680
rect 503622 167628 503628 167680
rect 503680 167668 503686 167680
rect 542998 167668 543004 167680
rect 503680 167640 543004 167668
rect 503680 167628 503686 167640
rect 542998 167628 543004 167640
rect 543056 167628 543062 167680
rect 252462 167560 252468 167612
rect 252520 167600 252526 167612
rect 258258 167600 258264 167612
rect 252520 167572 258264 167600
rect 252520 167560 252526 167572
rect 258258 167560 258264 167572
rect 258316 167560 258322 167612
rect 269850 167016 269856 167068
rect 269908 167056 269914 167068
rect 307478 167056 307484 167068
rect 269908 167028 307484 167056
rect 269908 167016 269914 167028
rect 307478 167016 307484 167028
rect 307536 167016 307542 167068
rect 166350 166948 166356 167000
rect 166408 166988 166414 167000
rect 214098 166988 214104 167000
rect 166408 166960 214104 166988
rect 166408 166948 166414 166960
rect 214098 166948 214104 166960
rect 214156 166948 214162 167000
rect 252370 166948 252376 167000
rect 252428 166988 252434 167000
rect 263686 166988 263692 167000
rect 252428 166960 263692 166988
rect 252428 166948 252434 166960
rect 263686 166948 263692 166960
rect 263744 166948 263750 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 334250 166988 334256 167000
rect 324372 166960 334256 166988
rect 324372 166948 324378 166960
rect 334250 166948 334256 166960
rect 334308 166948 334314 167000
rect 496906 166948 496912 167000
rect 496964 166988 496970 167000
rect 503898 166988 503904 167000
rect 496964 166960 503904 166988
rect 496964 166948 496970 166960
rect 503898 166948 503904 166960
rect 503956 166988 503962 167000
rect 504174 166988 504180 167000
rect 503956 166960 504180 166988
rect 503956 166948 503962 166960
rect 504174 166948 504180 166960
rect 504232 166948 504238 167000
rect 169202 166880 169208 166932
rect 169260 166920 169266 166932
rect 214006 166920 214012 166932
rect 169260 166892 214012 166920
rect 169260 166880 169266 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 252462 166880 252468 166932
rect 252520 166920 252526 166932
rect 261018 166920 261024 166932
rect 252520 166892 261024 166920
rect 252520 166880 252526 166892
rect 261018 166880 261024 166892
rect 261076 166880 261082 166932
rect 196802 166812 196808 166864
rect 196860 166852 196866 166864
rect 213914 166852 213920 166864
rect 196860 166824 213920 166852
rect 196860 166812 196866 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 252278 166812 252284 166864
rect 252336 166852 252342 166864
rect 256970 166852 256976 166864
rect 252336 166824 256976 166852
rect 252336 166812 252342 166824
rect 256970 166812 256976 166824
rect 257028 166812 257034 166864
rect 287790 166268 287796 166320
rect 287848 166308 287854 166320
rect 307294 166308 307300 166320
rect 287848 166280 307300 166308
rect 287848 166268 287854 166280
rect 307294 166268 307300 166280
rect 307352 166268 307358 166320
rect 504174 166268 504180 166320
rect 504232 166308 504238 166320
rect 555418 166308 555424 166320
rect 504232 166280 555424 166308
rect 504232 166268 504238 166280
rect 555418 166268 555424 166280
rect 555476 166268 555482 166320
rect 271322 165656 271328 165708
rect 271380 165696 271386 165708
rect 307662 165696 307668 165708
rect 271380 165668 307668 165696
rect 271380 165656 271386 165668
rect 307662 165656 307668 165668
rect 307720 165656 307726 165708
rect 257430 165588 257436 165640
rect 257488 165628 257494 165640
rect 306742 165628 306748 165640
rect 257488 165600 306748 165628
rect 257488 165588 257494 165600
rect 306742 165588 306748 165600
rect 306800 165588 306806 165640
rect 353938 165588 353944 165640
rect 353996 165628 354002 165640
rect 416774 165628 416780 165640
rect 353996 165600 416780 165628
rect 353996 165588 354002 165600
rect 416774 165588 416780 165600
rect 416832 165588 416838 165640
rect 556154 165588 556160 165640
rect 556212 165628 556218 165640
rect 580166 165628 580172 165640
rect 556212 165600 580172 165628
rect 556212 165588 556218 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 166258 165520 166264 165572
rect 166316 165560 166322 165572
rect 213914 165560 213920 165572
rect 166316 165532 213920 165560
rect 166316 165520 166322 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252462 165520 252468 165572
rect 252520 165560 252526 165572
rect 270494 165560 270500 165572
rect 252520 165532 270500 165560
rect 252520 165520 252526 165532
rect 270494 165520 270500 165532
rect 270552 165520 270558 165572
rect 324314 165520 324320 165572
rect 324372 165560 324378 165572
rect 335538 165560 335544 165572
rect 324372 165532 335544 165560
rect 324372 165520 324378 165532
rect 335538 165520 335544 165532
rect 335596 165520 335602 165572
rect 496998 165520 497004 165572
rect 497056 165560 497062 165572
rect 509326 165560 509332 165572
rect 497056 165532 509332 165560
rect 497056 165520 497062 165532
rect 509326 165520 509332 165532
rect 509384 165560 509390 165572
rect 510522 165560 510528 165572
rect 509384 165532 510528 165560
rect 509384 165520 509390 165532
rect 510522 165520 510528 165532
rect 510580 165520 510586 165572
rect 252278 165452 252284 165504
rect 252336 165492 252342 165504
rect 262398 165492 262404 165504
rect 252336 165464 262404 165492
rect 252336 165452 252342 165464
rect 262398 165452 262404 165464
rect 262456 165452 262462 165504
rect 324498 165452 324504 165504
rect 324556 165492 324562 165504
rect 331398 165492 331404 165504
rect 324556 165464 331404 165492
rect 324556 165452 324562 165464
rect 331398 165452 331404 165464
rect 331456 165452 331462 165504
rect 257522 164840 257528 164892
rect 257580 164880 257586 164892
rect 306558 164880 306564 164892
rect 257580 164852 306564 164880
rect 257580 164840 257586 164852
rect 306558 164840 306564 164852
rect 306616 164840 306622 164892
rect 496906 164840 496912 164892
rect 496964 164880 496970 164892
rect 501230 164880 501236 164892
rect 496964 164852 501236 164880
rect 496964 164840 496970 164852
rect 501230 164840 501236 164852
rect 501288 164880 501294 164892
rect 504358 164880 504364 164892
rect 501288 164852 504364 164880
rect 501288 164840 501294 164852
rect 504358 164840 504364 164852
rect 504416 164840 504422 164892
rect 510522 164840 510528 164892
rect 510580 164880 510586 164892
rect 525058 164880 525064 164892
rect 510580 164852 525064 164880
rect 510580 164840 510586 164852
rect 525058 164840 525064 164852
rect 525116 164840 525122 164892
rect 276658 164296 276664 164348
rect 276716 164336 276722 164348
rect 307110 164336 307116 164348
rect 276716 164308 307116 164336
rect 276716 164296 276722 164308
rect 307110 164296 307116 164308
rect 307168 164296 307174 164348
rect 252370 164228 252376 164280
rect 252428 164268 252434 164280
rect 259546 164268 259552 164280
rect 252428 164240 259552 164268
rect 252428 164228 252434 164240
rect 259546 164228 259552 164240
rect 259604 164228 259610 164280
rect 269758 164228 269764 164280
rect 269816 164268 269822 164280
rect 307662 164268 307668 164280
rect 269816 164240 307668 164268
rect 269816 164228 269822 164240
rect 307662 164228 307668 164240
rect 307720 164228 307726 164280
rect 334618 164228 334624 164280
rect 334676 164268 334682 164280
rect 416774 164268 416780 164280
rect 334676 164240 416780 164268
rect 334676 164228 334682 164240
rect 416774 164228 416780 164240
rect 416832 164228 416838 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 33778 164200 33784 164212
rect 3292 164172 33784 164200
rect 3292 164160 3298 164172
rect 33778 164160 33784 164172
rect 33836 164160 33842 164212
rect 171962 164160 171968 164212
rect 172020 164200 172026 164212
rect 214006 164200 214012 164212
rect 172020 164172 214012 164200
rect 172020 164160 172026 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 252462 164160 252468 164212
rect 252520 164200 252526 164212
rect 269114 164200 269120 164212
rect 252520 164172 269120 164200
rect 252520 164160 252526 164172
rect 269114 164160 269120 164172
rect 269172 164160 269178 164212
rect 324314 164160 324320 164212
rect 324372 164200 324378 164212
rect 332778 164200 332784 164212
rect 324372 164172 332784 164200
rect 324372 164160 324378 164172
rect 332778 164160 332784 164172
rect 332836 164160 332842 164212
rect 496906 164160 496912 164212
rect 496964 164200 496970 164212
rect 506658 164200 506664 164212
rect 496964 164172 506664 164200
rect 496964 164160 496970 164172
rect 506658 164160 506664 164172
rect 506716 164200 506722 164212
rect 556154 164200 556160 164212
rect 506716 164172 556160 164200
rect 506716 164160 506722 164172
rect 556154 164160 556160 164172
rect 556212 164160 556218 164212
rect 196894 164092 196900 164144
rect 196952 164132 196958 164144
rect 213914 164132 213920 164144
rect 196952 164104 213920 164132
rect 196952 164092 196958 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 252370 164092 252376 164144
rect 252428 164132 252434 164144
rect 256786 164132 256792 164144
rect 252428 164104 256792 164132
rect 252428 164092 252434 164104
rect 256786 164092 256792 164104
rect 256844 164092 256850 164144
rect 268562 163548 268568 163600
rect 268620 163588 268626 163600
rect 307478 163588 307484 163600
rect 268620 163560 307484 163588
rect 268620 163548 268626 163560
rect 307478 163548 307484 163560
rect 307536 163548 307542 163600
rect 261478 163480 261484 163532
rect 261536 163520 261542 163532
rect 307386 163520 307392 163532
rect 261536 163492 307392 163520
rect 261536 163480 261542 163492
rect 307386 163480 307392 163492
rect 307444 163480 307450 163532
rect 286410 162868 286416 162920
rect 286468 162908 286474 162920
rect 307662 162908 307668 162920
rect 286468 162880 307668 162908
rect 286468 162868 286474 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 170490 162800 170496 162852
rect 170548 162840 170554 162852
rect 213914 162840 213920 162852
rect 170548 162812 213920 162840
rect 170548 162800 170554 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252370 162800 252376 162852
rect 252428 162840 252434 162852
rect 266354 162840 266360 162852
rect 252428 162812 266360 162840
rect 252428 162800 252434 162812
rect 266354 162800 266360 162812
rect 266412 162800 266418 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 342346 162840 342352 162852
rect 324372 162812 342352 162840
rect 324372 162800 324378 162812
rect 342346 162800 342352 162812
rect 342404 162800 342410 162852
rect 496906 162800 496912 162852
rect 496964 162840 496970 162852
rect 512638 162840 512644 162852
rect 496964 162812 512644 162840
rect 496964 162800 496970 162812
rect 512638 162800 512644 162812
rect 512696 162800 512702 162852
rect 178770 162732 178776 162784
rect 178828 162772 178834 162784
rect 214006 162772 214012 162784
rect 178828 162744 214012 162772
rect 178828 162732 178834 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 252462 162732 252468 162784
rect 252520 162772 252526 162784
rect 265158 162772 265164 162784
rect 252520 162744 265164 162772
rect 252520 162732 252526 162744
rect 265158 162732 265164 162744
rect 265216 162732 265222 162784
rect 274082 162120 274088 162172
rect 274140 162160 274146 162172
rect 306742 162160 306748 162172
rect 274140 162132 306748 162160
rect 274140 162120 274146 162132
rect 306742 162120 306748 162132
rect 306800 162120 306806 162172
rect 304258 161576 304264 161628
rect 304316 161616 304322 161628
rect 307478 161616 307484 161628
rect 304316 161588 307484 161616
rect 304316 161576 304322 161588
rect 307478 161576 307484 161588
rect 307536 161576 307542 161628
rect 278130 161508 278136 161560
rect 278188 161548 278194 161560
rect 307570 161548 307576 161560
rect 278188 161520 307576 161548
rect 278188 161508 278194 161520
rect 307570 161508 307576 161520
rect 307628 161508 307634 161560
rect 262950 161440 262956 161492
rect 263008 161480 263014 161492
rect 307662 161480 307668 161492
rect 263008 161452 307668 161480
rect 263008 161440 263014 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 345658 161440 345664 161492
rect 345716 161480 345722 161492
rect 416774 161480 416780 161492
rect 345716 161452 416780 161480
rect 345716 161440 345722 161452
rect 416774 161440 416780 161452
rect 416832 161440 416838 161492
rect 169110 161372 169116 161424
rect 169168 161412 169174 161424
rect 213914 161412 213920 161424
rect 169168 161384 213920 161412
rect 169168 161372 169174 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252462 161372 252468 161424
rect 252520 161412 252526 161424
rect 261110 161412 261116 161424
rect 252520 161384 261116 161412
rect 252520 161372 252526 161384
rect 261110 161372 261116 161384
rect 261168 161372 261174 161424
rect 496906 161372 496912 161424
rect 496964 161412 496970 161424
rect 535454 161412 535460 161424
rect 496964 161384 535460 161412
rect 496964 161372 496970 161384
rect 535454 161372 535460 161384
rect 535512 161372 535518 161424
rect 173158 161304 173164 161356
rect 173216 161344 173222 161356
rect 214006 161344 214012 161356
rect 173216 161316 214012 161344
rect 173216 161304 173222 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 301498 160216 301504 160268
rect 301556 160256 301562 160268
rect 307570 160256 307576 160268
rect 301556 160228 307576 160256
rect 301556 160216 301562 160228
rect 307570 160216 307576 160228
rect 307628 160216 307634 160268
rect 324314 160216 324320 160268
rect 324372 160256 324378 160268
rect 327442 160256 327448 160268
rect 324372 160228 327448 160256
rect 324372 160216 324378 160228
rect 327442 160216 327448 160228
rect 327500 160216 327506 160268
rect 264330 160148 264336 160200
rect 264388 160188 264394 160200
rect 307662 160188 307668 160200
rect 264388 160160 307668 160188
rect 264388 160148 264394 160160
rect 307662 160148 307668 160160
rect 307720 160148 307726 160200
rect 253474 160080 253480 160132
rect 253532 160120 253538 160132
rect 307478 160120 307484 160132
rect 253532 160092 307484 160120
rect 253532 160080 253538 160092
rect 307478 160080 307484 160092
rect 307536 160080 307542 160132
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 331490 160052 331496 160064
rect 324372 160024 331496 160052
rect 324372 160012 324378 160024
rect 331490 160012 331496 160024
rect 331548 160012 331554 160064
rect 496906 160012 496912 160064
rect 496964 160052 496970 160064
rect 529934 160052 529940 160064
rect 496964 160024 529940 160052
rect 496964 160012 496970 160024
rect 529934 160012 529940 160024
rect 529992 160012 529998 160064
rect 496998 159944 497004 159996
rect 497056 159984 497062 159996
rect 503714 159984 503720 159996
rect 497056 159956 503720 159984
rect 497056 159944 497062 159956
rect 503714 159944 503720 159956
rect 503772 159944 503778 159996
rect 167638 159332 167644 159384
rect 167696 159372 167702 159384
rect 214006 159372 214012 159384
rect 167696 159344 214012 159372
rect 167696 159332 167702 159344
rect 214006 159332 214012 159344
rect 214064 159332 214070 159384
rect 293402 158856 293408 158908
rect 293460 158896 293466 158908
rect 306558 158896 306564 158908
rect 293460 158868 306564 158896
rect 293460 158856 293466 158868
rect 306558 158856 306564 158868
rect 306616 158856 306622 158908
rect 260466 158788 260472 158840
rect 260524 158828 260530 158840
rect 307662 158828 307668 158840
rect 260524 158800 307668 158828
rect 260524 158788 260530 158800
rect 307662 158788 307668 158800
rect 307720 158788 307726 158840
rect 258810 158720 258816 158772
rect 258868 158760 258874 158772
rect 307570 158760 307576 158772
rect 258868 158732 307576 158760
rect 258868 158720 258874 158732
rect 307570 158720 307576 158732
rect 307628 158720 307634 158772
rect 167822 158652 167828 158704
rect 167880 158692 167886 158704
rect 213914 158692 213920 158704
rect 167880 158664 213920 158692
rect 167880 158652 167886 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 251358 158652 251364 158704
rect 251416 158692 251422 158704
rect 253934 158692 253940 158704
rect 251416 158664 253940 158692
rect 251416 158652 251422 158664
rect 253934 158652 253940 158664
rect 253992 158652 253998 158704
rect 324314 158652 324320 158704
rect 324372 158692 324378 158704
rect 336918 158692 336924 158704
rect 324372 158664 336924 158692
rect 324372 158652 324378 158664
rect 336918 158652 336924 158664
rect 336976 158652 336982 158704
rect 496906 158652 496912 158704
rect 496964 158692 496970 158704
rect 517606 158692 517612 158704
rect 496964 158664 517612 158692
rect 496964 158652 496970 158664
rect 517606 158652 517612 158664
rect 517664 158692 517670 158704
rect 544378 158692 544384 158704
rect 517664 158664 544384 158692
rect 517664 158652 517670 158664
rect 544378 158652 544384 158664
rect 544436 158652 544442 158704
rect 252186 158584 252192 158636
rect 252244 158624 252250 158636
rect 255498 158624 255504 158636
rect 252244 158596 255504 158624
rect 252244 158584 252250 158596
rect 255498 158584 255504 158596
rect 255556 158584 255562 158636
rect 251910 157972 251916 158024
rect 251968 158012 251974 158024
rect 264238 158012 264244 158024
rect 251968 157984 264244 158012
rect 251968 157972 251974 157984
rect 264238 157972 264244 157984
rect 264296 157972 264302 158024
rect 287882 157496 287888 157548
rect 287940 157536 287946 157548
rect 306558 157536 306564 157548
rect 287940 157508 306564 157536
rect 287940 157496 287946 157508
rect 306558 157496 306564 157508
rect 306616 157496 306622 157548
rect 266998 157428 267004 157480
rect 267056 157468 267062 157480
rect 307662 157468 307668 157480
rect 267056 157440 307668 157468
rect 267056 157428 267062 157440
rect 307662 157428 307668 157440
rect 307720 157428 307726 157480
rect 263594 157360 263600 157412
rect 263652 157400 263658 157412
rect 307478 157400 307484 157412
rect 263652 157372 307484 157400
rect 263652 157360 263658 157372
rect 307478 157360 307484 157372
rect 307536 157360 307542 157412
rect 331858 157360 331864 157412
rect 331916 157400 331922 157412
rect 416774 157400 416780 157412
rect 331916 157372 416780 157400
rect 331916 157360 331922 157372
rect 416774 157360 416780 157372
rect 416832 157360 416838 157412
rect 205082 157292 205088 157344
rect 205140 157332 205146 157344
rect 213914 157332 213920 157344
rect 205140 157304 213920 157332
rect 205140 157292 205146 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 273254 157332 273260 157344
rect 252520 157304 273260 157332
rect 252520 157292 252526 157304
rect 273254 157292 273260 157304
rect 273312 157292 273318 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 338298 157332 338304 157344
rect 324372 157304 338304 157332
rect 324372 157292 324378 157304
rect 338298 157292 338304 157304
rect 338356 157292 338362 157344
rect 496906 157292 496912 157344
rect 496964 157332 496970 157344
rect 582374 157332 582380 157344
rect 496964 157304 582380 157332
rect 496964 157292 496970 157304
rect 582374 157292 582380 157304
rect 582432 157292 582438 157344
rect 252370 157224 252376 157276
rect 252428 157264 252434 157276
rect 263778 157264 263784 157276
rect 252428 157236 263784 157264
rect 252428 157224 252434 157236
rect 263778 157224 263784 157236
rect 263836 157224 263842 157276
rect 285030 156068 285036 156120
rect 285088 156108 285094 156120
rect 307662 156108 307668 156120
rect 285088 156080 307668 156108
rect 285088 156068 285094 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 272702 156000 272708 156052
rect 272760 156040 272766 156052
rect 306558 156040 306564 156052
rect 272760 156012 306564 156040
rect 272760 156000 272766 156012
rect 306558 156000 306564 156012
rect 306616 156000 306622 156052
rect 260190 155932 260196 155984
rect 260248 155972 260254 155984
rect 307570 155972 307576 155984
rect 260248 155944 307576 155972
rect 260248 155932 260254 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 335998 155932 336004 155984
rect 336056 155972 336062 155984
rect 416774 155972 416780 155984
rect 336056 155944 416780 155972
rect 336056 155932 336062 155944
rect 416774 155932 416780 155944
rect 416832 155932 416838 155984
rect 171870 155864 171876 155916
rect 171928 155904 171934 155916
rect 214006 155904 214012 155916
rect 171928 155876 214012 155904
rect 171928 155864 171934 155876
rect 214006 155864 214012 155876
rect 214064 155864 214070 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 331306 155904 331312 155916
rect 324372 155876 331312 155904
rect 324372 155864 324378 155876
rect 331306 155864 331312 155876
rect 331364 155864 331370 155916
rect 496906 155864 496912 155916
rect 496964 155904 496970 155916
rect 519538 155904 519544 155916
rect 496964 155876 519544 155904
rect 496964 155864 496970 155876
rect 519538 155864 519544 155876
rect 519596 155864 519602 155916
rect 196710 155796 196716 155848
rect 196768 155836 196774 155848
rect 213914 155836 213920 155848
rect 196768 155808 213920 155836
rect 196768 155796 196774 155808
rect 213914 155796 213920 155808
rect 213972 155796 213978 155848
rect 170582 155184 170588 155236
rect 170640 155224 170646 155236
rect 214558 155224 214564 155236
rect 170640 155196 214564 155224
rect 170640 155184 170646 155196
rect 214558 155184 214564 155196
rect 214616 155184 214622 155236
rect 272794 155184 272800 155236
rect 272852 155224 272858 155236
rect 307386 155224 307392 155236
rect 272852 155196 307392 155224
rect 272852 155184 272858 155196
rect 307386 155184 307392 155196
rect 307444 155184 307450 155236
rect 262858 154640 262864 154692
rect 262916 154680 262922 154692
rect 307570 154680 307576 154692
rect 262916 154652 307576 154680
rect 262916 154640 262922 154652
rect 307570 154640 307576 154652
rect 307628 154640 307634 154692
rect 261754 154572 261760 154624
rect 261812 154612 261818 154624
rect 307662 154612 307668 154624
rect 261812 154584 307668 154612
rect 261812 154572 261818 154584
rect 307662 154572 307668 154584
rect 307720 154572 307726 154624
rect 356790 154572 356796 154624
rect 356848 154612 356854 154624
rect 416774 154612 416780 154624
rect 356848 154584 416780 154612
rect 356848 154572 356854 154584
rect 416774 154572 416780 154584
rect 416832 154572 416838 154624
rect 251542 154504 251548 154556
rect 251600 154544 251606 154556
rect 254210 154544 254216 154556
rect 251600 154516 254216 154544
rect 251600 154504 251606 154516
rect 254210 154504 254216 154516
rect 254268 154504 254274 154556
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 341058 154544 341064 154556
rect 324372 154516 341064 154544
rect 324372 154504 324378 154516
rect 341058 154504 341064 154516
rect 341116 154504 341122 154556
rect 496998 154504 497004 154556
rect 497056 154544 497062 154556
rect 505278 154544 505284 154556
rect 497056 154516 505284 154544
rect 497056 154504 497062 154516
rect 505278 154504 505284 154516
rect 505336 154504 505342 154556
rect 252462 154436 252468 154488
rect 252520 154476 252526 154488
rect 267826 154476 267832 154488
rect 252520 154448 267832 154476
rect 252520 154436 252526 154448
rect 267826 154436 267832 154448
rect 267884 154436 267890 154488
rect 324406 154436 324412 154488
rect 324464 154476 324470 154488
rect 328730 154476 328736 154488
rect 324464 154448 328736 154476
rect 324464 154436 324470 154448
rect 328730 154436 328736 154448
rect 328788 154436 328794 154488
rect 496906 154436 496912 154488
rect 496964 154476 496970 154488
rect 502518 154476 502524 154488
rect 496964 154448 502524 154476
rect 496964 154436 496970 154448
rect 502518 154436 502524 154448
rect 502576 154436 502582 154488
rect 252370 154368 252376 154420
rect 252428 154408 252434 154420
rect 274726 154408 274732 154420
rect 252428 154380 274732 154408
rect 252428 154368 252434 154380
rect 274726 154368 274732 154380
rect 274784 154368 274790 154420
rect 251818 153824 251824 153876
rect 251876 153864 251882 153876
rect 263594 153864 263600 153876
rect 251876 153836 263600 153864
rect 251876 153824 251882 153836
rect 263594 153824 263600 153836
rect 263652 153824 263658 153876
rect 267090 153824 267096 153876
rect 267148 153864 267154 153876
rect 307478 153864 307484 153876
rect 267148 153836 307484 153864
rect 267148 153824 267154 153836
rect 307478 153824 307484 153836
rect 307536 153824 307542 153876
rect 174538 153280 174544 153332
rect 174596 153320 174602 153332
rect 214006 153320 214012 153332
rect 174596 153292 214012 153320
rect 174596 153280 174602 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 302970 153280 302976 153332
rect 303028 153320 303034 153332
rect 307662 153320 307668 153332
rect 303028 153292 307668 153320
rect 303028 153280 303034 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 166258 153212 166264 153264
rect 166316 153252 166322 153264
rect 213914 153252 213920 153264
rect 166316 153224 213920 153252
rect 166316 153212 166322 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 298738 153212 298744 153264
rect 298796 153252 298802 153264
rect 306558 153252 306564 153264
rect 298796 153224 306564 153252
rect 298796 153212 298802 153224
rect 306558 153212 306564 153224
rect 306616 153212 306622 153264
rect 360838 153212 360844 153264
rect 360896 153252 360902 153264
rect 416774 153252 416780 153264
rect 360896 153224 416780 153252
rect 360896 153212 360902 153224
rect 416774 153212 416780 153224
rect 416832 153212 416838 153264
rect 252370 153144 252376 153196
rect 252428 153184 252434 153196
rect 271966 153184 271972 153196
rect 252428 153156 271972 153184
rect 252428 153144 252434 153156
rect 271966 153144 271972 153156
rect 272024 153144 272030 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 330018 153184 330024 153196
rect 324372 153156 330024 153184
rect 324372 153144 324378 153156
rect 330018 153144 330024 153156
rect 330076 153144 330082 153196
rect 252278 153076 252284 153128
rect 252336 153116 252342 153128
rect 269206 153116 269212 153128
rect 252336 153088 269212 153116
rect 252336 153076 252342 153088
rect 269206 153076 269212 153088
rect 269264 153076 269270 153128
rect 252462 153008 252468 153060
rect 252520 153048 252526 153060
rect 266446 153048 266452 153060
rect 252520 153020 266452 153048
rect 252520 153008 252526 153020
rect 266446 153008 266452 153020
rect 266504 153008 266510 153060
rect 496906 152600 496912 152652
rect 496964 152640 496970 152652
rect 498470 152640 498476 152652
rect 496964 152612 498476 152640
rect 496964 152600 496970 152612
rect 498470 152600 498476 152612
rect 498528 152600 498534 152652
rect 276842 152464 276848 152516
rect 276900 152504 276906 152516
rect 307662 152504 307668 152516
rect 276900 152476 307668 152504
rect 276900 152464 276906 152476
rect 307662 152464 307668 152476
rect 307720 152464 307726 152516
rect 189718 151784 189724 151836
rect 189776 151824 189782 151836
rect 213914 151824 213920 151836
rect 189776 151796 213920 151824
rect 189776 151784 189782 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 258718 151784 258724 151836
rect 258776 151824 258782 151836
rect 307662 151824 307668 151836
rect 258776 151796 307668 151824
rect 258776 151784 258782 151796
rect 307662 151784 307668 151796
rect 307720 151784 307726 151836
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 339586 151756 339592 151768
rect 324372 151728 339592 151756
rect 324372 151716 324378 151728
rect 339586 151716 339592 151728
rect 339644 151716 339650 151768
rect 252370 151648 252376 151700
rect 252428 151688 252434 151700
rect 271874 151688 271880 151700
rect 252428 151660 271880 151688
rect 252428 151648 252434 151660
rect 271874 151648 271880 151660
rect 271932 151648 271938 151700
rect 252462 151580 252468 151632
rect 252520 151620 252526 151632
rect 276106 151620 276112 151632
rect 252520 151592 276112 151620
rect 252520 151580 252526 151592
rect 276106 151580 276112 151592
rect 276164 151580 276170 151632
rect 252278 151444 252284 151496
rect 252336 151484 252342 151496
rect 254118 151484 254124 151496
rect 252336 151456 254124 151484
rect 252336 151444 252342 151456
rect 254118 151444 254124 151456
rect 254176 151444 254182 151496
rect 256142 151036 256148 151088
rect 256200 151076 256206 151088
rect 306650 151076 306656 151088
rect 256200 151048 306656 151076
rect 256200 151036 256206 151048
rect 306650 151036 306656 151048
rect 306708 151036 306714 151088
rect 303062 150560 303068 150612
rect 303120 150600 303126 150612
rect 307662 150600 307668 150612
rect 303120 150572 307668 150600
rect 303120 150560 303126 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 209130 150492 209136 150544
rect 209188 150532 209194 150544
rect 214006 150532 214012 150544
rect 209188 150504 214012 150532
rect 209188 150492 209194 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 289262 150492 289268 150544
rect 289320 150532 289326 150544
rect 307294 150532 307300 150544
rect 289320 150504 307300 150532
rect 289320 150492 289326 150504
rect 307294 150492 307300 150504
rect 307352 150492 307358 150544
rect 196710 150424 196716 150476
rect 196768 150464 196774 150476
rect 213914 150464 213920 150476
rect 196768 150436 213920 150464
rect 196768 150424 196774 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 264238 150424 264244 150476
rect 264296 150464 264302 150476
rect 306926 150464 306932 150476
rect 264296 150436 306932 150464
rect 264296 150424 264302 150436
rect 306926 150424 306932 150436
rect 306984 150424 306990 150476
rect 359550 150424 359556 150476
rect 359608 150464 359614 150476
rect 416774 150464 416780 150476
rect 359608 150436 416780 150464
rect 359608 150424 359614 150436
rect 416774 150424 416780 150436
rect 416832 150424 416838 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 15838 150396 15844 150408
rect 3476 150368 15844 150396
rect 3476 150356 3482 150368
rect 15838 150356 15844 150368
rect 15896 150356 15902 150408
rect 170398 150356 170404 150408
rect 170456 150396 170462 150408
rect 214006 150396 214012 150408
rect 170456 150368 214012 150396
rect 170456 150356 170462 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 252462 150356 252468 150408
rect 252520 150396 252526 150408
rect 264974 150396 264980 150408
rect 252520 150368 264980 150396
rect 252520 150356 252526 150368
rect 264974 150356 264980 150368
rect 265032 150356 265038 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 335446 150396 335452 150408
rect 324372 150368 335452 150396
rect 324372 150356 324378 150368
rect 335446 150356 335452 150368
rect 335504 150356 335510 150408
rect 496814 150356 496820 150408
rect 496872 150396 496878 150408
rect 506566 150396 506572 150408
rect 496872 150368 506572 150396
rect 496872 150356 496878 150368
rect 506566 150356 506572 150368
rect 506624 150356 506630 150408
rect 252278 150288 252284 150340
rect 252336 150328 252342 150340
rect 255590 150328 255596 150340
rect 252336 150300 255596 150328
rect 252336 150288 252342 150300
rect 255590 150288 255596 150300
rect 255648 150288 255654 150340
rect 324406 150288 324412 150340
rect 324464 150328 324470 150340
rect 333974 150328 333980 150340
rect 324464 150300 333980 150328
rect 324464 150288 324470 150300
rect 333974 150288 333980 150300
rect 334032 150288 334038 150340
rect 287974 149200 287980 149252
rect 288032 149240 288038 149252
rect 306926 149240 306932 149252
rect 288032 149212 306932 149240
rect 288032 149200 288038 149212
rect 306926 149200 306932 149212
rect 306984 149200 306990 149252
rect 279510 149132 279516 149184
rect 279568 149172 279574 149184
rect 306558 149172 306564 149184
rect 279568 149144 306564 149172
rect 279568 149132 279574 149144
rect 306558 149132 306564 149144
rect 306616 149132 306622 149184
rect 265710 149064 265716 149116
rect 265768 149104 265774 149116
rect 307294 149104 307300 149116
rect 265768 149076 307300 149104
rect 265768 149064 265774 149076
rect 307294 149064 307300 149076
rect 307352 149064 307358 149116
rect 363598 149064 363604 149116
rect 363656 149104 363662 149116
rect 416774 149104 416780 149116
rect 363656 149076 416780 149104
rect 363656 149064 363662 149076
rect 416774 149064 416780 149076
rect 416832 149064 416838 149116
rect 169018 148996 169024 149048
rect 169076 149036 169082 149048
rect 213914 149036 213920 149048
rect 169076 149008 213920 149036
rect 169076 148996 169082 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 278774 149036 278780 149048
rect 252520 149008 278780 149036
rect 252520 148996 252526 149008
rect 278774 148996 278780 149008
rect 278832 148996 278838 149048
rect 324406 148996 324412 149048
rect 324464 149036 324470 149048
rect 342438 149036 342444 149048
rect 324464 149008 342444 149036
rect 324464 148996 324470 149008
rect 342438 148996 342444 149008
rect 342496 148996 342502 149048
rect 496814 148996 496820 149048
rect 496872 149036 496878 149048
rect 505186 149036 505192 149048
rect 496872 149008 505192 149036
rect 496872 148996 496878 149008
rect 505186 148996 505192 149008
rect 505244 148996 505250 149048
rect 252370 148928 252376 148980
rect 252428 148968 252434 148980
rect 254026 148968 254032 148980
rect 252428 148940 254032 148968
rect 252428 148928 252434 148940
rect 254026 148928 254032 148940
rect 254084 148928 254090 148980
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 329926 148968 329932 148980
rect 324372 148940 329932 148968
rect 324372 148928 324378 148940
rect 329926 148928 329932 148940
rect 329984 148928 329990 148980
rect 286594 147772 286600 147824
rect 286652 147812 286658 147824
rect 307478 147812 307484 147824
rect 286652 147784 307484 147812
rect 286652 147772 286658 147784
rect 307478 147772 307484 147784
rect 307536 147772 307542 147824
rect 257338 147704 257344 147756
rect 257396 147744 257402 147756
rect 307570 147744 307576 147756
rect 257396 147716 307576 147744
rect 257396 147704 257402 147716
rect 307570 147704 307576 147716
rect 307628 147704 307634 147756
rect 256234 147636 256240 147688
rect 256292 147676 256298 147688
rect 307662 147676 307668 147688
rect 256292 147648 307668 147676
rect 256292 147636 256298 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 369854 147636 369860 147688
rect 369912 147676 369918 147688
rect 416774 147676 416780 147688
rect 369912 147648 416780 147676
rect 369912 147636 369918 147648
rect 416774 147636 416780 147648
rect 416832 147636 416838 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 280154 147608 280160 147620
rect 252520 147580 280160 147608
rect 252520 147568 252526 147580
rect 280154 147568 280160 147580
rect 280212 147568 280218 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 352006 147608 352012 147620
rect 324372 147580 352012 147608
rect 324372 147568 324378 147580
rect 352006 147568 352012 147580
rect 352064 147568 352070 147620
rect 496814 147568 496820 147620
rect 496872 147608 496878 147620
rect 510798 147608 510804 147620
rect 496872 147580 510804 147608
rect 496872 147568 496878 147580
rect 510798 147568 510804 147580
rect 510856 147568 510862 147620
rect 252094 147500 252100 147552
rect 252152 147540 252158 147552
rect 255314 147540 255320 147552
rect 252152 147512 255320 147540
rect 252152 147500 252158 147512
rect 255314 147500 255320 147512
rect 255372 147500 255378 147552
rect 249886 147296 249892 147348
rect 249944 147296 249950 147348
rect 249794 147092 249800 147144
rect 249852 147132 249858 147144
rect 249904 147132 249932 147296
rect 249852 147104 249932 147132
rect 249852 147092 249858 147104
rect 300302 146412 300308 146464
rect 300360 146452 300366 146464
rect 307570 146452 307576 146464
rect 300360 146424 307576 146452
rect 300360 146412 300366 146424
rect 307570 146412 307576 146424
rect 307628 146412 307634 146464
rect 209222 146344 209228 146396
rect 209280 146384 209286 146396
rect 214006 146384 214012 146396
rect 209280 146356 214012 146384
rect 209280 146344 209286 146356
rect 214006 146344 214012 146356
rect 214064 146344 214070 146396
rect 269942 146344 269948 146396
rect 270000 146384 270006 146396
rect 307662 146384 307668 146396
rect 270000 146356 307668 146384
rect 270000 146344 270006 146356
rect 307662 146344 307668 146356
rect 307720 146344 307726 146396
rect 176010 146276 176016 146328
rect 176068 146316 176074 146328
rect 213914 146316 213920 146328
rect 176068 146288 213920 146316
rect 176068 146276 176074 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 254762 146276 254768 146328
rect 254820 146316 254826 146328
rect 307478 146316 307484 146328
rect 254820 146288 307484 146316
rect 254820 146276 254826 146288
rect 307478 146276 307484 146288
rect 307536 146276 307542 146328
rect 356698 146276 356704 146328
rect 356756 146316 356762 146328
rect 416774 146316 416780 146328
rect 356756 146288 416780 146316
rect 356756 146276 356762 146288
rect 416774 146276 416780 146288
rect 416832 146276 416838 146328
rect 252462 146208 252468 146260
rect 252520 146248 252526 146260
rect 273346 146248 273352 146260
rect 252520 146220 273352 146248
rect 252520 146208 252526 146220
rect 273346 146208 273352 146220
rect 273404 146208 273410 146260
rect 324406 146208 324412 146260
rect 324464 146248 324470 146260
rect 350626 146248 350632 146260
rect 324464 146220 350632 146248
rect 324464 146208 324470 146220
rect 350626 146208 350632 146220
rect 350684 146208 350690 146260
rect 252370 146140 252376 146192
rect 252428 146180 252434 146192
rect 270586 146180 270592 146192
rect 252428 146152 270592 146180
rect 252428 146140 252434 146152
rect 270586 146140 270592 146152
rect 270644 146140 270650 146192
rect 324314 146140 324320 146192
rect 324372 146180 324378 146192
rect 328454 146180 328460 146192
rect 324372 146152 328460 146180
rect 324372 146140 324378 146152
rect 328454 146140 328460 146152
rect 328512 146140 328518 146192
rect 496814 145664 496820 145716
rect 496872 145704 496878 145716
rect 499666 145704 499672 145716
rect 496872 145676 499672 145704
rect 496872 145664 496878 145676
rect 499666 145664 499672 145676
rect 499724 145664 499730 145716
rect 255958 145596 255964 145648
rect 256016 145636 256022 145648
rect 306926 145636 306932 145648
rect 256016 145608 306932 145636
rect 256016 145596 256022 145608
rect 306926 145596 306932 145608
rect 306984 145596 306990 145648
rect 254946 145528 254952 145580
rect 255004 145568 255010 145580
rect 307202 145568 307208 145580
rect 255004 145540 307208 145568
rect 255004 145528 255010 145540
rect 307202 145528 307208 145540
rect 307260 145528 307266 145580
rect 171870 144916 171876 144968
rect 171928 144956 171934 144968
rect 213914 144956 213920 144968
rect 171928 144928 213920 144956
rect 171928 144916 171934 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 296162 144916 296168 144968
rect 296220 144956 296226 144968
rect 306926 144956 306932 144968
rect 296220 144928 306932 144956
rect 296220 144916 296226 144928
rect 306926 144916 306932 144928
rect 306984 144916 306990 144968
rect 252370 144848 252376 144900
rect 252428 144888 252434 144900
rect 262306 144888 262312 144900
rect 252428 144860 262312 144888
rect 252428 144848 252434 144860
rect 262306 144848 262312 144860
rect 262364 144848 262370 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 260834 144820 260840 144832
rect 252520 144792 260840 144820
rect 252520 144780 252526 144792
rect 260834 144780 260840 144792
rect 260892 144780 260898 144832
rect 169018 144168 169024 144220
rect 169076 144208 169082 144220
rect 214650 144208 214656 144220
rect 169076 144180 214656 144208
rect 169076 144168 169082 144180
rect 214650 144168 214656 144180
rect 214708 144168 214714 144220
rect 264514 144168 264520 144220
rect 264572 144208 264578 144220
rect 307478 144208 307484 144220
rect 264572 144180 307484 144208
rect 264572 144168 264578 144180
rect 307478 144168 307484 144180
rect 307536 144168 307542 144220
rect 507762 144168 507768 144220
rect 507820 144208 507826 144220
rect 511994 144208 512000 144220
rect 507820 144180 512000 144208
rect 507820 144168 507826 144180
rect 511994 144168 512000 144180
rect 512052 144168 512058 144220
rect 280890 143624 280896 143676
rect 280948 143664 280954 143676
rect 306558 143664 306564 143676
rect 280948 143636 306564 143664
rect 280948 143624 280954 143636
rect 306558 143624 306564 143636
rect 306616 143624 306622 143676
rect 187142 143556 187148 143608
rect 187200 143596 187206 143608
rect 213914 143596 213920 143608
rect 187200 143568 213920 143596
rect 187200 143556 187206 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 253382 143556 253388 143608
rect 253440 143596 253446 143608
rect 307662 143596 307668 143608
rect 253440 143568 307668 143596
rect 253440 143556 253446 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 342346 143556 342352 143608
rect 342404 143596 342410 143608
rect 416866 143596 416872 143608
rect 342404 143568 416872 143596
rect 342404 143556 342410 143568
rect 416866 143556 416872 143568
rect 416924 143556 416930 143608
rect 496814 143556 496820 143608
rect 496872 143596 496878 143608
rect 507762 143596 507768 143608
rect 496872 143568 507768 143596
rect 496872 143556 496878 143568
rect 507762 143556 507768 143568
rect 507820 143556 507826 143608
rect 252462 143488 252468 143540
rect 252520 143528 252526 143540
rect 265066 143528 265072 143540
rect 252520 143500 265072 143528
rect 252520 143488 252526 143500
rect 265066 143488 265072 143500
rect 265124 143488 265130 143540
rect 324314 143488 324320 143540
rect 324372 143528 324378 143540
rect 332686 143528 332692 143540
rect 324372 143500 332692 143528
rect 324372 143488 324378 143500
rect 332686 143488 332692 143500
rect 332744 143488 332750 143540
rect 342254 143488 342260 143540
rect 342312 143528 342318 143540
rect 416774 143528 416780 143540
rect 342312 143500 416780 143528
rect 342312 143488 342318 143500
rect 416774 143488 416780 143500
rect 416832 143488 416838 143540
rect 252370 143420 252376 143472
rect 252428 143460 252434 143472
rect 258350 143460 258356 143472
rect 252428 143432 258356 143460
rect 252428 143420 252434 143432
rect 258350 143420 258356 143432
rect 258408 143420 258414 143472
rect 257614 142808 257620 142860
rect 257672 142848 257678 142860
rect 307110 142848 307116 142860
rect 257672 142820 307116 142848
rect 257672 142808 257678 142820
rect 307110 142808 307116 142820
rect 307168 142808 307174 142860
rect 333238 142808 333244 142860
rect 333296 142848 333302 142860
rect 342254 142848 342260 142860
rect 333296 142820 342260 142848
rect 333296 142808 333302 142820
rect 342254 142808 342260 142820
rect 342312 142808 342318 142860
rect 211890 142264 211896 142316
rect 211948 142304 211954 142316
rect 214466 142304 214472 142316
rect 211948 142276 214472 142304
rect 211948 142264 211954 142276
rect 214466 142264 214472 142276
rect 214524 142264 214530 142316
rect 283742 142196 283748 142248
rect 283800 142236 283806 142248
rect 307662 142236 307668 142248
rect 283800 142208 307668 142236
rect 283800 142196 283806 142208
rect 307662 142196 307668 142208
rect 307720 142196 307726 142248
rect 181530 142128 181536 142180
rect 181588 142168 181594 142180
rect 213914 142168 213920 142180
rect 181588 142140 213920 142168
rect 181588 142128 181594 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 253198 142128 253204 142180
rect 253256 142168 253262 142180
rect 307570 142168 307576 142180
rect 253256 142140 307576 142168
rect 253256 142128 253262 142140
rect 307570 142128 307576 142140
rect 307628 142128 307634 142180
rect 496906 142128 496912 142180
rect 496964 142168 496970 142180
rect 513282 142168 513288 142180
rect 496964 142140 513288 142168
rect 496964 142128 496970 142140
rect 513282 142128 513288 142140
rect 513340 142128 513346 142180
rect 324406 142060 324412 142112
rect 324464 142100 324470 142112
rect 349154 142100 349160 142112
rect 324464 142072 349160 142100
rect 324464 142060 324470 142072
rect 349154 142060 349160 142072
rect 349212 142060 349218 142112
rect 353294 142060 353300 142112
rect 353352 142100 353358 142112
rect 416774 142100 416780 142112
rect 353352 142072 416780 142100
rect 353352 142060 353358 142072
rect 416774 142060 416780 142072
rect 416832 142060 416838 142112
rect 496814 142060 496820 142112
rect 496872 142100 496878 142112
rect 512086 142100 512092 142112
rect 496872 142072 512092 142100
rect 496872 142060 496878 142072
rect 512086 142060 512092 142072
rect 512144 142100 512150 142112
rect 519538 142100 519544 142112
rect 512144 142072 519544 142100
rect 512144 142060 512150 142072
rect 519538 142060 519544 142072
rect 519596 142060 519602 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 328546 142032 328552 142044
rect 324372 142004 328552 142032
rect 324372 141992 324378 142004
rect 328546 141992 328552 142004
rect 328604 141992 328610 142044
rect 253658 141380 253664 141432
rect 253716 141420 253722 141432
rect 307018 141420 307024 141432
rect 253716 141392 307024 141420
rect 253716 141380 253722 141392
rect 307018 141380 307024 141392
rect 307076 141380 307082 141432
rect 496814 141380 496820 141432
rect 496872 141420 496878 141432
rect 516134 141420 516140 141432
rect 496872 141392 516140 141420
rect 496872 141380 496878 141392
rect 516134 141380 516140 141392
rect 516192 141380 516198 141432
rect 174630 140836 174636 140888
rect 174688 140876 174694 140888
rect 214006 140876 214012 140888
rect 174688 140848 214012 140876
rect 174688 140836 174694 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 290642 140836 290648 140888
rect 290700 140876 290706 140888
rect 307570 140876 307576 140888
rect 290700 140848 307576 140876
rect 290700 140836 290706 140848
rect 307570 140836 307576 140848
rect 307628 140836 307634 140888
rect 170398 140768 170404 140820
rect 170456 140808 170462 140820
rect 213914 140808 213920 140820
rect 170456 140780 213920 140808
rect 170456 140768 170462 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 254854 140768 254860 140820
rect 254912 140808 254918 140820
rect 307662 140808 307668 140820
rect 254912 140780 307668 140808
rect 254912 140768 254918 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 352650 140768 352656 140820
rect 352708 140808 352714 140820
rect 353294 140808 353300 140820
rect 352708 140780 353300 140808
rect 352708 140768 352714 140780
rect 353294 140768 353300 140780
rect 353352 140768 353358 140820
rect 252370 140700 252376 140752
rect 252428 140740 252434 140752
rect 277486 140740 277492 140752
rect 252428 140712 277492 140740
rect 252428 140700 252434 140712
rect 277486 140700 277492 140712
rect 277544 140700 277550 140752
rect 496814 140700 496820 140752
rect 496872 140740 496878 140752
rect 502978 140740 502984 140752
rect 496872 140712 502984 140740
rect 496872 140700 496878 140712
rect 502978 140700 502984 140712
rect 503036 140700 503042 140752
rect 252462 140632 252468 140684
rect 252520 140672 252526 140684
rect 276014 140672 276020 140684
rect 252520 140644 276020 140672
rect 252520 140632 252526 140644
rect 276014 140632 276020 140644
rect 276072 140632 276078 140684
rect 167914 140020 167920 140072
rect 167972 140060 167978 140072
rect 209130 140060 209136 140072
rect 167972 140032 209136 140060
rect 167972 140020 167978 140032
rect 209130 140020 209136 140032
rect 209188 140020 209194 140072
rect 516134 140020 516140 140072
rect 516192 140060 516198 140072
rect 580166 140060 580172 140072
rect 516192 140032 580172 140060
rect 516192 140020 516198 140032
rect 580166 140020 580172 140032
rect 580224 140020 580230 140072
rect 252002 139748 252008 139800
rect 252060 139788 252066 139800
rect 260466 139788 260472 139800
rect 252060 139760 260472 139788
rect 252060 139748 252066 139760
rect 260466 139748 260472 139760
rect 260524 139748 260530 139800
rect 294782 139544 294788 139596
rect 294840 139584 294846 139596
rect 307570 139584 307576 139596
rect 294840 139556 307576 139584
rect 294840 139544 294846 139556
rect 307570 139544 307576 139556
rect 307628 139544 307634 139596
rect 210510 139476 210516 139528
rect 210568 139516 210574 139528
rect 214006 139516 214012 139528
rect 210568 139488 214012 139516
rect 210568 139476 210574 139488
rect 214006 139476 214012 139488
rect 214064 139476 214070 139528
rect 260098 139476 260104 139528
rect 260156 139516 260162 139528
rect 307662 139516 307668 139528
rect 260156 139488 307668 139516
rect 260156 139476 260162 139488
rect 307662 139476 307668 139488
rect 307720 139476 307726 139528
rect 206462 139408 206468 139460
rect 206520 139448 206526 139460
rect 213914 139448 213920 139460
rect 206520 139420 213920 139448
rect 206520 139408 206526 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 256050 139408 256056 139460
rect 256108 139448 256114 139460
rect 307478 139448 307484 139460
rect 256108 139420 307484 139448
rect 256108 139408 256114 139420
rect 307478 139408 307484 139420
rect 307536 139408 307542 139460
rect 367738 139408 367744 139460
rect 367796 139448 367802 139460
rect 416774 139448 416780 139460
rect 367796 139420 416780 139448
rect 367796 139408 367802 139420
rect 416774 139408 416780 139420
rect 416832 139408 416838 139460
rect 252462 139340 252468 139392
rect 252520 139380 252526 139392
rect 280246 139380 280252 139392
rect 252520 139352 280252 139380
rect 252520 139340 252526 139352
rect 280246 139340 280252 139352
rect 280304 139340 280310 139392
rect 496814 139340 496820 139392
rect 496872 139380 496878 139392
rect 514846 139380 514852 139392
rect 496872 139352 514852 139380
rect 496872 139340 496878 139352
rect 514846 139340 514852 139352
rect 514904 139340 514910 139392
rect 324314 139068 324320 139120
rect 324372 139108 324378 139120
rect 325970 139108 325976 139120
rect 324372 139080 325976 139108
rect 324372 139068 324378 139080
rect 325970 139068 325976 139080
rect 326028 139068 326034 139120
rect 202322 138048 202328 138100
rect 202380 138088 202386 138100
rect 214006 138088 214012 138100
rect 202380 138060 214012 138088
rect 202380 138048 202386 138060
rect 214006 138048 214012 138060
rect 214064 138048 214070 138100
rect 286502 138048 286508 138100
rect 286560 138088 286566 138100
rect 307662 138088 307668 138100
rect 286560 138060 307668 138088
rect 286560 138048 286566 138060
rect 307662 138048 307668 138060
rect 307720 138048 307726 138100
rect 170490 137980 170496 138032
rect 170548 138020 170554 138032
rect 213914 138020 213920 138032
rect 170548 137992 213920 138020
rect 170548 137980 170554 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 250622 137980 250628 138032
rect 250680 138020 250686 138032
rect 307570 138020 307576 138032
rect 250680 137992 307576 138020
rect 250680 137980 250686 137992
rect 307570 137980 307576 137992
rect 307628 137980 307634 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 14458 137952 14464 137964
rect 3292 137924 14464 137952
rect 3292 137912 3298 137924
rect 14458 137912 14464 137924
rect 14516 137912 14522 137964
rect 252370 137912 252376 137964
rect 252428 137952 252434 137964
rect 281534 137952 281540 137964
rect 252428 137924 281540 137952
rect 252428 137912 252434 137924
rect 281534 137912 281540 137924
rect 281592 137912 281598 137964
rect 324406 137912 324412 137964
rect 324464 137952 324470 137964
rect 346486 137952 346492 137964
rect 324464 137924 346492 137952
rect 324464 137912 324470 137924
rect 346486 137912 346492 137924
rect 346544 137912 346550 137964
rect 496814 137912 496820 137964
rect 496872 137952 496878 137964
rect 520918 137952 520924 137964
rect 496872 137924 520924 137952
rect 496872 137912 496878 137924
rect 520918 137912 520924 137924
rect 520976 137912 520982 137964
rect 252462 137844 252468 137896
rect 252520 137884 252526 137896
rect 267734 137884 267740 137896
rect 252520 137856 267740 137884
rect 252520 137844 252526 137856
rect 267734 137844 267740 137856
rect 267792 137844 267798 137896
rect 324314 137844 324320 137896
rect 324372 137884 324378 137896
rect 338114 137884 338120 137896
rect 324372 137856 338120 137884
rect 324372 137844 324378 137856
rect 338114 137844 338120 137856
rect 338172 137844 338178 137896
rect 252094 137232 252100 137284
rect 252152 137272 252158 137284
rect 267182 137272 267188 137284
rect 252152 137244 267188 137272
rect 252152 137232 252158 137244
rect 267182 137232 267188 137244
rect 267240 137232 267246 137284
rect 275278 137232 275284 137284
rect 275336 137272 275342 137284
rect 307386 137272 307392 137284
rect 275336 137244 307392 137272
rect 275336 137232 275342 137244
rect 307386 137232 307392 137244
rect 307444 137232 307450 137284
rect 253290 136892 253296 136944
rect 253348 136932 253354 136944
rect 253658 136932 253664 136944
rect 253348 136904 253664 136932
rect 253348 136892 253354 136904
rect 253658 136892 253664 136904
rect 253716 136892 253722 136944
rect 268378 136688 268384 136740
rect 268436 136728 268442 136740
rect 307662 136728 307668 136740
rect 268436 136700 307668 136728
rect 268436 136688 268442 136700
rect 307662 136688 307668 136700
rect 307720 136688 307726 136740
rect 198182 136620 198188 136672
rect 198240 136660 198246 136672
rect 213914 136660 213920 136672
rect 198240 136632 213920 136660
rect 198240 136620 198246 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 250530 136620 250536 136672
rect 250588 136660 250594 136672
rect 307110 136660 307116 136672
rect 250588 136632 307116 136660
rect 250588 136620 250594 136632
rect 307110 136620 307116 136632
rect 307168 136620 307174 136672
rect 370498 136620 370504 136672
rect 370556 136660 370562 136672
rect 416774 136660 416780 136672
rect 370556 136632 416780 136660
rect 370556 136620 370562 136632
rect 416774 136620 416780 136632
rect 416832 136620 416838 136672
rect 252186 136552 252192 136604
rect 252244 136592 252250 136604
rect 296254 136592 296260 136604
rect 252244 136564 296260 136592
rect 252244 136552 252250 136564
rect 296254 136552 296260 136564
rect 296312 136552 296318 136604
rect 324314 136552 324320 136604
rect 324372 136592 324378 136604
rect 352190 136592 352196 136604
rect 324372 136564 352196 136592
rect 324372 136552 324378 136564
rect 352190 136552 352196 136564
rect 352248 136552 352254 136604
rect 496906 136552 496912 136604
rect 496964 136592 496970 136604
rect 508498 136592 508504 136604
rect 496964 136564 508504 136592
rect 496964 136552 496970 136564
rect 508498 136552 508504 136564
rect 508556 136552 508562 136604
rect 252370 136484 252376 136536
rect 252428 136524 252434 136536
rect 285214 136524 285220 136536
rect 252428 136496 285220 136524
rect 252428 136484 252434 136496
rect 285214 136484 285220 136496
rect 285272 136484 285278 136536
rect 496814 136484 496820 136536
rect 496872 136524 496878 136536
rect 502426 136524 502432 136536
rect 496872 136496 502432 136524
rect 496872 136484 496878 136496
rect 502426 136484 502432 136496
rect 502484 136484 502490 136536
rect 252462 136416 252468 136468
rect 252520 136456 252526 136468
rect 277394 136456 277400 136468
rect 252520 136428 277400 136456
rect 252520 136416 252526 136428
rect 277394 136416 277400 136428
rect 277452 136416 277458 136468
rect 252278 136348 252284 136400
rect 252336 136388 252342 136400
rect 265802 136388 265808 136400
rect 252336 136360 265808 136388
rect 252336 136348 252342 136360
rect 265802 136348 265808 136360
rect 265860 136348 265866 136400
rect 295978 135464 295984 135516
rect 296036 135504 296042 135516
rect 307110 135504 307116 135516
rect 296036 135476 307116 135504
rect 296036 135464 296042 135476
rect 307110 135464 307116 135476
rect 307168 135464 307174 135516
rect 284938 135396 284944 135448
rect 284996 135436 285002 135448
rect 307662 135436 307668 135448
rect 284996 135408 307668 135436
rect 284996 135396 285002 135408
rect 307662 135396 307668 135408
rect 307720 135396 307726 135448
rect 207750 135328 207756 135380
rect 207808 135368 207814 135380
rect 214006 135368 214012 135380
rect 207808 135340 214012 135368
rect 207808 135328 207814 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 283558 135328 283564 135380
rect 283616 135368 283622 135380
rect 307570 135368 307576 135380
rect 283616 135340 307576 135368
rect 283616 135328 283622 135340
rect 307570 135328 307576 135340
rect 307628 135328 307634 135380
rect 178770 135260 178776 135312
rect 178828 135300 178834 135312
rect 213914 135300 213920 135312
rect 178828 135272 213920 135300
rect 178828 135260 178834 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 265618 135260 265624 135312
rect 265676 135300 265682 135312
rect 307478 135300 307484 135312
rect 265676 135272 307484 135300
rect 265676 135260 265682 135272
rect 307478 135260 307484 135272
rect 307536 135260 307542 135312
rect 376018 135260 376024 135312
rect 376076 135300 376082 135312
rect 416774 135300 416780 135312
rect 376076 135272 416780 135300
rect 376076 135260 376082 135272
rect 416774 135260 416780 135272
rect 416832 135260 416838 135312
rect 252462 135192 252468 135244
rect 252520 135232 252526 135244
rect 280798 135232 280804 135244
rect 252520 135204 280804 135232
rect 252520 135192 252526 135204
rect 280798 135192 280804 135204
rect 280856 135192 280862 135244
rect 340230 135192 340236 135244
rect 340288 135232 340294 135244
rect 417326 135232 417332 135244
rect 340288 135204 417332 135232
rect 340288 135192 340294 135204
rect 417326 135192 417332 135204
rect 417384 135192 417390 135244
rect 252370 135124 252376 135176
rect 252428 135164 252434 135176
rect 263042 135164 263048 135176
rect 252428 135136 263048 135164
rect 252428 135124 252434 135136
rect 263042 135124 263048 135136
rect 263100 135124 263106 135176
rect 324314 135124 324320 135176
rect 324372 135164 324378 135176
rect 350534 135164 350540 135176
rect 324372 135136 350540 135164
rect 324372 135124 324378 135136
rect 350534 135124 350540 135136
rect 350592 135124 350598 135176
rect 324406 135056 324412 135108
rect 324464 135096 324470 135108
rect 346578 135096 346584 135108
rect 324464 135068 346584 135096
rect 324464 135056 324470 135068
rect 346578 135056 346584 135068
rect 346636 135056 346642 135108
rect 276934 134512 276940 134564
rect 276992 134552 276998 134564
rect 307294 134552 307300 134564
rect 276992 134524 307300 134552
rect 276992 134512 276998 134524
rect 307294 134512 307300 134524
rect 307352 134512 307358 134564
rect 300118 133968 300124 134020
rect 300176 134008 300182 134020
rect 307570 134008 307576 134020
rect 300176 133980 307576 134008
rect 300176 133968 300182 133980
rect 307570 133968 307576 133980
rect 307628 133968 307634 134020
rect 177482 133900 177488 133952
rect 177540 133940 177546 133952
rect 213914 133940 213920 133952
rect 177540 133912 213920 133940
rect 177540 133900 177546 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 282270 133900 282276 133952
rect 282328 133940 282334 133952
rect 307662 133940 307668 133952
rect 282328 133912 307668 133940
rect 282328 133900 282334 133912
rect 307662 133900 307668 133912
rect 307720 133900 307726 133952
rect 252370 133832 252376 133884
rect 252428 133872 252434 133884
rect 283650 133872 283656 133884
rect 252428 133844 283656 133872
rect 252428 133832 252434 133844
rect 283650 133832 283656 133844
rect 283708 133832 283714 133884
rect 374638 133832 374644 133884
rect 374696 133872 374702 133884
rect 419350 133872 419356 133884
rect 374696 133844 419356 133872
rect 374696 133832 374702 133844
rect 419350 133832 419356 133844
rect 419408 133832 419414 133884
rect 496814 133832 496820 133884
rect 496872 133872 496878 133884
rect 503806 133872 503812 133884
rect 496872 133844 503812 133872
rect 496872 133832 496878 133844
rect 503806 133832 503812 133844
rect 503864 133832 503870 133884
rect 252462 133764 252468 133816
rect 252520 133804 252526 133816
rect 260374 133804 260380 133816
rect 252520 133776 260380 133804
rect 252520 133764 252526 133776
rect 260374 133764 260380 133776
rect 260432 133764 260438 133816
rect 324314 133560 324320 133612
rect 324372 133600 324378 133612
rect 327258 133600 327264 133612
rect 324372 133572 327264 133600
rect 324372 133560 324378 133572
rect 327258 133560 327264 133572
rect 327316 133560 327322 133612
rect 260466 133152 260472 133204
rect 260524 133192 260530 133204
rect 306834 133192 306840 133204
rect 260524 133164 306840 133192
rect 260524 133152 260530 133164
rect 306834 133152 306840 133164
rect 306892 133152 306898 133204
rect 386322 133152 386328 133204
rect 386380 133192 386386 133204
rect 419626 133192 419632 133204
rect 386380 133164 419632 133192
rect 386380 133152 386386 133164
rect 419626 133152 419632 133164
rect 419684 133152 419690 133204
rect 304350 132608 304356 132660
rect 304408 132648 304414 132660
rect 306926 132648 306932 132660
rect 304408 132620 306932 132648
rect 304408 132608 304414 132620
rect 306926 132608 306932 132620
rect 306984 132608 306990 132660
rect 297450 132540 297456 132592
rect 297508 132580 297514 132592
rect 307662 132580 307668 132592
rect 297508 132552 307668 132580
rect 297508 132540 297514 132552
rect 307662 132540 307668 132552
rect 307720 132540 307726 132592
rect 254670 132472 254676 132524
rect 254728 132512 254734 132524
rect 307570 132512 307576 132524
rect 254728 132484 307576 132512
rect 254728 132472 254734 132484
rect 307570 132472 307576 132484
rect 307628 132472 307634 132524
rect 252462 132404 252468 132456
rect 252520 132444 252526 132456
rect 300210 132444 300216 132456
rect 252520 132416 300216 132444
rect 252520 132404 252526 132416
rect 300210 132404 300216 132416
rect 300268 132404 300274 132456
rect 411898 132404 411904 132456
rect 411956 132444 411962 132456
rect 417326 132444 417332 132456
rect 411956 132416 417332 132444
rect 411956 132404 411962 132416
rect 417326 132404 417332 132416
rect 417384 132404 417390 132456
rect 252370 132336 252376 132388
rect 252428 132376 252434 132388
rect 285122 132376 285128 132388
rect 252428 132348 285128 132376
rect 252428 132336 252434 132348
rect 285122 132336 285128 132348
rect 285180 132336 285186 132388
rect 252462 132268 252468 132320
rect 252520 132308 252526 132320
rect 268470 132308 268476 132320
rect 252520 132280 268476 132308
rect 252520 132268 252526 132280
rect 268470 132268 268476 132280
rect 268528 132268 268534 132320
rect 301590 131248 301596 131300
rect 301648 131288 301654 131300
rect 307662 131288 307668 131300
rect 301648 131260 307668 131288
rect 301648 131248 301654 131260
rect 307662 131248 307668 131260
rect 307720 131248 307726 131300
rect 180242 131180 180248 131232
rect 180300 131220 180306 131232
rect 214006 131220 214012 131232
rect 180300 131192 214012 131220
rect 180300 131180 180306 131192
rect 214006 131180 214012 131192
rect 214064 131180 214070 131232
rect 289078 131180 289084 131232
rect 289136 131220 289142 131232
rect 306558 131220 306564 131232
rect 289136 131192 306564 131220
rect 289136 131180 289142 131192
rect 306558 131180 306564 131192
rect 306616 131180 306622 131232
rect 171962 131112 171968 131164
rect 172020 131152 172026 131164
rect 213914 131152 213920 131164
rect 172020 131124 213920 131152
rect 172020 131112 172026 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 278038 131112 278044 131164
rect 278096 131152 278102 131164
rect 307570 131152 307576 131164
rect 278096 131124 307576 131152
rect 278096 131112 278102 131124
rect 307570 131112 307576 131124
rect 307628 131112 307634 131164
rect 252462 131044 252468 131096
rect 252520 131084 252526 131096
rect 297358 131084 297364 131096
rect 252520 131056 297364 131084
rect 252520 131044 252526 131056
rect 297358 131044 297364 131056
rect 297416 131044 297422 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 349338 131084 349344 131096
rect 324372 131056 349344 131084
rect 324372 131044 324378 131056
rect 349338 131044 349344 131056
rect 349396 131044 349402 131096
rect 496814 131044 496820 131096
rect 496872 131084 496878 131096
rect 509234 131084 509240 131096
rect 496872 131056 509240 131084
rect 496872 131044 496878 131056
rect 509234 131044 509240 131056
rect 509292 131044 509298 131096
rect 252370 130976 252376 131028
rect 252428 131016 252434 131028
rect 264422 131016 264428 131028
rect 252428 130988 264428 131016
rect 252428 130976 252434 130988
rect 264422 130976 264428 130988
rect 264480 130976 264486 131028
rect 252462 130432 252468 130484
rect 252520 130472 252526 130484
rect 260282 130472 260288 130484
rect 252520 130444 260288 130472
rect 252520 130432 252526 130444
rect 260282 130432 260288 130444
rect 260340 130432 260346 130484
rect 297542 129888 297548 129940
rect 297600 129928 297606 129940
rect 307662 129928 307668 129940
rect 297600 129900 307668 129928
rect 297600 129888 297606 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 205082 129820 205088 129872
rect 205140 129860 205146 129872
rect 214006 129860 214012 129872
rect 205140 129832 214012 129860
rect 205140 129820 205146 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 294598 129820 294604 129872
rect 294656 129860 294662 129872
rect 307570 129860 307576 129872
rect 294656 129832 307576 129860
rect 294656 129820 294662 129832
rect 307570 129820 307576 129832
rect 307628 129820 307634 129872
rect 173250 129752 173256 129804
rect 173308 129792 173314 129804
rect 213914 129792 213920 129804
rect 173308 129764 213920 129792
rect 173308 129752 173314 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 261570 129752 261576 129804
rect 261628 129792 261634 129804
rect 307294 129792 307300 129804
rect 261628 129764 307300 129792
rect 261628 129752 261634 129764
rect 307294 129752 307300 129764
rect 307352 129752 307358 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 269850 129724 269856 129736
rect 252520 129696 269856 129724
rect 252520 129684 252526 129696
rect 269850 129684 269856 129696
rect 269908 129684 269914 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 334158 129724 334164 129736
rect 324372 129696 334164 129724
rect 324372 129684 324378 129696
rect 334158 129684 334164 129696
rect 334216 129684 334222 129736
rect 496814 129684 496820 129736
rect 496872 129724 496878 129736
rect 514754 129724 514760 129736
rect 496872 129696 514760 129724
rect 496872 129684 496878 129696
rect 514754 129684 514760 129696
rect 514812 129684 514818 129736
rect 252370 129616 252376 129668
rect 252428 129656 252434 129668
rect 257522 129656 257528 129668
rect 252428 129628 257528 129656
rect 252428 129616 252434 129628
rect 257522 129616 257528 129628
rect 257580 129616 257586 129668
rect 252186 129412 252192 129464
rect 252244 129452 252250 129464
rect 257430 129452 257436 129464
rect 252244 129424 257436 129452
rect 252244 129412 252250 129424
rect 257430 129412 257436 129424
rect 257488 129412 257494 129464
rect 297358 128392 297364 128444
rect 297416 128432 297422 128444
rect 307570 128432 307576 128444
rect 297416 128404 307576 128432
rect 297416 128392 297422 128404
rect 307570 128392 307576 128404
rect 307628 128392 307634 128444
rect 273990 128324 273996 128376
rect 274048 128364 274054 128376
rect 307662 128364 307668 128376
rect 274048 128336 307668 128364
rect 274048 128324 274054 128336
rect 307662 128324 307668 128336
rect 307720 128324 307726 128376
rect 252370 128256 252376 128308
rect 252428 128296 252434 128308
rect 287790 128296 287796 128308
rect 252428 128268 287796 128296
rect 252428 128256 252434 128268
rect 287790 128256 287796 128268
rect 287848 128256 287854 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 338206 128296 338212 128308
rect 324372 128268 338212 128296
rect 324372 128256 324378 128268
rect 338206 128256 338212 128268
rect 338264 128256 338270 128308
rect 382918 128256 382924 128308
rect 382976 128296 382982 128308
rect 417602 128296 417608 128308
rect 382976 128268 417608 128296
rect 382976 128256 382982 128268
rect 417602 128256 417608 128268
rect 417660 128256 417666 128308
rect 496814 128256 496820 128308
rect 496872 128296 496878 128308
rect 507854 128296 507860 128308
rect 496872 128268 507860 128296
rect 496872 128256 496878 128268
rect 507854 128256 507860 128268
rect 507912 128256 507918 128308
rect 252278 128188 252284 128240
rect 252336 128228 252342 128240
rect 271322 128228 271328 128240
rect 252336 128200 271328 128228
rect 252336 128188 252342 128200
rect 271322 128188 271328 128200
rect 271380 128188 271386 128240
rect 324406 128188 324412 128240
rect 324464 128228 324470 128240
rect 330110 128228 330116 128240
rect 324464 128200 330116 128228
rect 324464 128188 324470 128200
rect 330110 128188 330116 128200
rect 330168 128188 330174 128240
rect 252462 128120 252468 128172
rect 252520 128160 252526 128172
rect 261478 128160 261484 128172
rect 252520 128132 261484 128160
rect 252520 128120 252526 128132
rect 261478 128120 261484 128132
rect 261536 128120 261542 128172
rect 270034 127576 270040 127628
rect 270092 127616 270098 127628
rect 307202 127616 307208 127628
rect 270092 127588 307208 127616
rect 270092 127576 270098 127588
rect 307202 127576 307208 127588
rect 307260 127576 307266 127628
rect 525058 127576 525064 127628
rect 525116 127616 525122 127628
rect 580166 127616 580172 127628
rect 525116 127588 580172 127616
rect 525116 127576 525122 127588
rect 580166 127576 580172 127588
rect 580224 127576 580230 127628
rect 287698 127032 287704 127084
rect 287756 127072 287762 127084
rect 306558 127072 306564 127084
rect 287756 127044 306564 127072
rect 287756 127032 287762 127044
rect 306558 127032 306564 127044
rect 306616 127032 306622 127084
rect 173158 126964 173164 127016
rect 173216 127004 173222 127016
rect 213914 127004 213920 127016
rect 173216 126976 213920 127004
rect 173216 126964 173222 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 271230 126964 271236 127016
rect 271288 127004 271294 127016
rect 307662 127004 307668 127016
rect 271288 126976 307668 127004
rect 271288 126964 271294 126976
rect 307662 126964 307668 126976
rect 307720 126964 307726 127016
rect 252462 126896 252468 126948
rect 252520 126936 252526 126948
rect 268562 126936 268568 126948
rect 252520 126908 268568 126936
rect 252520 126896 252526 126908
rect 268562 126896 268568 126908
rect 268620 126896 268626 126948
rect 251910 126828 251916 126880
rect 251968 126868 251974 126880
rect 254946 126868 254952 126880
rect 251968 126840 254952 126868
rect 251968 126828 251974 126840
rect 254946 126828 254952 126840
rect 255004 126828 255010 126880
rect 496814 126488 496820 126540
rect 496872 126528 496878 126540
rect 499850 126528 499856 126540
rect 496872 126500 499856 126528
rect 496872 126488 496878 126500
rect 499850 126488 499856 126500
rect 499908 126488 499914 126540
rect 292022 125740 292028 125792
rect 292080 125780 292086 125792
rect 307570 125780 307576 125792
rect 292080 125752 307576 125780
rect 292080 125740 292086 125752
rect 307570 125740 307576 125752
rect 307628 125740 307634 125792
rect 176102 125672 176108 125724
rect 176160 125712 176166 125724
rect 213914 125712 213920 125724
rect 176160 125684 213920 125712
rect 176160 125672 176166 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 268470 125672 268476 125724
rect 268528 125712 268534 125724
rect 307662 125712 307668 125724
rect 268528 125684 307668 125712
rect 268528 125672 268534 125684
rect 307662 125672 307668 125684
rect 307720 125672 307726 125724
rect 57790 125604 57796 125656
rect 57848 125644 57854 125656
rect 65150 125644 65156 125656
rect 57848 125616 65156 125644
rect 57848 125604 57854 125616
rect 65150 125604 65156 125616
rect 65208 125604 65214 125656
rect 167638 125604 167644 125656
rect 167696 125644 167702 125656
rect 214006 125644 214012 125656
rect 167696 125616 214012 125644
rect 167696 125604 167702 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 254578 125604 254584 125656
rect 254636 125644 254642 125656
rect 306558 125644 306564 125656
rect 254636 125616 306564 125644
rect 254636 125604 254642 125616
rect 306558 125604 306564 125616
rect 306616 125604 306622 125656
rect 252278 125536 252284 125588
rect 252336 125576 252342 125588
rect 276658 125576 276664 125588
rect 252336 125548 276664 125576
rect 252336 125536 252342 125548
rect 276658 125536 276664 125548
rect 276716 125536 276722 125588
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 347958 125576 347964 125588
rect 324372 125548 347964 125576
rect 324372 125536 324378 125548
rect 347958 125536 347964 125548
rect 348016 125536 348022 125588
rect 496814 125536 496820 125588
rect 496872 125576 496878 125588
rect 517514 125576 517520 125588
rect 496872 125548 517520 125576
rect 496872 125536 496878 125548
rect 517514 125536 517520 125548
rect 517572 125536 517578 125588
rect 252462 125468 252468 125520
rect 252520 125508 252526 125520
rect 269758 125508 269764 125520
rect 252520 125480 269764 125508
rect 252520 125468 252526 125480
rect 269758 125468 269764 125480
rect 269816 125468 269822 125520
rect 324406 125468 324412 125520
rect 324464 125508 324470 125520
rect 343634 125508 343640 125520
rect 324464 125480 343640 125508
rect 324464 125468 324470 125480
rect 343634 125468 343640 125480
rect 343692 125468 343698 125520
rect 252370 125400 252376 125452
rect 252428 125440 252434 125452
rect 253290 125440 253296 125452
rect 252428 125412 253296 125440
rect 252428 125400 252434 125412
rect 253290 125400 253296 125412
rect 253348 125400 253354 125452
rect 252370 124856 252376 124908
rect 252428 124896 252434 124908
rect 305638 124896 305644 124908
rect 252428 124868 305644 124896
rect 252428 124856 252434 124868
rect 305638 124856 305644 124868
rect 305696 124856 305702 124908
rect 302878 124312 302884 124364
rect 302936 124352 302942 124364
rect 307662 124352 307668 124364
rect 302936 124324 307668 124352
rect 302936 124312 302942 124324
rect 307662 124312 307668 124324
rect 307720 124312 307726 124364
rect 193858 124244 193864 124296
rect 193916 124284 193922 124296
rect 214006 124284 214012 124296
rect 193916 124256 214012 124284
rect 193916 124244 193922 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 280798 124244 280804 124296
rect 280856 124284 280862 124296
rect 307570 124284 307576 124296
rect 280856 124256 307576 124284
rect 280856 124244 280862 124256
rect 307570 124244 307576 124256
rect 307628 124244 307634 124296
rect 185670 124176 185676 124228
rect 185728 124216 185734 124228
rect 213914 124216 213920 124228
rect 185728 124188 213920 124216
rect 185728 124176 185734 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 279418 124176 279424 124228
rect 279476 124216 279482 124228
rect 307294 124216 307300 124228
rect 279476 124188 307300 124216
rect 279476 124176 279482 124188
rect 307294 124176 307300 124188
rect 307352 124176 307358 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 274082 124148 274088 124160
rect 252520 124120 274088 124148
rect 252520 124108 252526 124120
rect 274082 124108 274088 124120
rect 274140 124108 274146 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 357434 124148 357440 124160
rect 324372 124120 357440 124148
rect 324372 124108 324378 124120
rect 357434 124108 357440 124120
rect 357492 124108 357498 124160
rect 496906 124108 496912 124160
rect 496964 124148 496970 124160
rect 505094 124148 505100 124160
rect 496964 124120 505100 124148
rect 496964 124108 496970 124120
rect 505094 124108 505100 124120
rect 505152 124108 505158 124160
rect 324406 124040 324412 124092
rect 324464 124080 324470 124092
rect 343910 124080 343916 124092
rect 324464 124052 343916 124080
rect 324464 124040 324470 124052
rect 343910 124040 343916 124052
rect 343968 124040 343974 124092
rect 496814 124040 496820 124092
rect 496872 124080 496878 124092
rect 499758 124080 499764 124092
rect 496872 124052 499764 124080
rect 496872 124040 496878 124052
rect 499758 124040 499764 124052
rect 499816 124040 499822 124092
rect 252094 123156 252100 123208
rect 252152 123196 252158 123208
rect 256234 123196 256240 123208
rect 252152 123168 256240 123196
rect 252152 123156 252158 123168
rect 256234 123156 256240 123168
rect 256292 123156 256298 123208
rect 272610 122952 272616 123004
rect 272668 122992 272674 123004
rect 307570 122992 307576 123004
rect 272668 122964 307576 122992
rect 272668 122952 272674 122964
rect 307570 122952 307576 122964
rect 307628 122952 307634 123004
rect 184290 122884 184296 122936
rect 184348 122924 184354 122936
rect 214006 122924 214012 122936
rect 184348 122896 214012 122924
rect 184348 122884 184354 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 298830 122884 298836 122936
rect 298888 122924 298894 122936
rect 307662 122924 307668 122936
rect 298888 122896 307668 122924
rect 298888 122884 298894 122896
rect 307662 122884 307668 122896
rect 307720 122884 307726 122936
rect 56502 122816 56508 122868
rect 56560 122856 56566 122868
rect 66070 122856 66076 122868
rect 56560 122828 66076 122856
rect 56560 122816 56566 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 170582 122816 170588 122868
rect 170640 122856 170646 122868
rect 213914 122856 213920 122868
rect 170640 122828 213920 122856
rect 170640 122816 170646 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 304258 122788 304264 122800
rect 252520 122760 304264 122788
rect 252520 122748 252526 122760
rect 304258 122748 304264 122760
rect 304316 122748 304322 122800
rect 324406 122748 324412 122800
rect 324464 122788 324470 122800
rect 347866 122788 347872 122800
rect 324464 122760 347872 122788
rect 324464 122748 324470 122760
rect 347866 122748 347872 122760
rect 347924 122748 347930 122800
rect 382182 122748 382188 122800
rect 382240 122788 382246 122800
rect 416774 122788 416780 122800
rect 382240 122760 416780 122788
rect 382240 122748 382246 122760
rect 416774 122748 416780 122760
rect 416832 122748 416838 122800
rect 496814 122748 496820 122800
rect 496872 122788 496878 122800
rect 521654 122788 521660 122800
rect 496872 122760 521660 122788
rect 496872 122748 496878 122760
rect 521654 122748 521660 122760
rect 521712 122748 521718 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 278130 122720 278136 122732
rect 252428 122692 278136 122720
rect 252428 122680 252434 122692
rect 278130 122680 278136 122692
rect 278188 122680 278194 122732
rect 324314 122680 324320 122732
rect 324372 122720 324378 122732
rect 345290 122720 345296 122732
rect 324372 122692 345296 122720
rect 324372 122680 324378 122692
rect 345290 122680 345296 122692
rect 345348 122680 345354 122732
rect 252278 122612 252284 122664
rect 252336 122652 252342 122664
rect 262950 122652 262956 122664
rect 252336 122624 262956 122652
rect 252336 122612 252342 122624
rect 262950 122612 262956 122624
rect 263008 122612 263014 122664
rect 182910 121524 182916 121576
rect 182968 121564 182974 121576
rect 213914 121564 213920 121576
rect 182968 121536 213920 121564
rect 182968 121524 182974 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 293310 121524 293316 121576
rect 293368 121564 293374 121576
rect 307570 121564 307576 121576
rect 293368 121536 307576 121564
rect 293368 121524 293374 121536
rect 307570 121524 307576 121536
rect 307628 121524 307634 121576
rect 167822 121456 167828 121508
rect 167880 121496 167886 121508
rect 214006 121496 214012 121508
rect 167880 121468 214012 121496
rect 167880 121456 167886 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 285122 121456 285128 121508
rect 285180 121496 285186 121508
rect 307662 121496 307668 121508
rect 285180 121468 307668 121496
rect 285180 121456 285186 121468
rect 307662 121456 307668 121468
rect 307720 121456 307726 121508
rect 252462 121388 252468 121440
rect 252520 121428 252526 121440
rect 301498 121428 301504 121440
rect 252520 121400 301504 121428
rect 252520 121388 252526 121400
rect 301498 121388 301504 121400
rect 301556 121388 301562 121440
rect 324406 121388 324412 121440
rect 324464 121428 324470 121440
rect 356054 121428 356060 121440
rect 324464 121400 356060 121428
rect 324464 121388 324470 121400
rect 356054 121388 356060 121400
rect 356112 121388 356118 121440
rect 388438 121388 388444 121440
rect 388496 121428 388502 121440
rect 416774 121428 416780 121440
rect 388496 121400 416780 121428
rect 388496 121388 388502 121400
rect 416774 121388 416780 121400
rect 416832 121388 416838 121440
rect 252370 121320 252376 121372
rect 252428 121360 252434 121372
rect 264330 121360 264336 121372
rect 252428 121332 264336 121360
rect 252428 121320 252434 121332
rect 264330 121320 264336 121332
rect 264388 121320 264394 121372
rect 324314 121320 324320 121372
rect 324372 121360 324378 121372
rect 328638 121360 328644 121372
rect 324372 121332 328644 121360
rect 324372 121320 324378 121332
rect 328638 121320 328644 121332
rect 328696 121320 328702 121372
rect 252278 121252 252284 121304
rect 252336 121292 252342 121304
rect 253474 121292 253480 121304
rect 252336 121264 253480 121292
rect 252336 121252 252342 121264
rect 253474 121252 253480 121264
rect 253532 121252 253538 121304
rect 304442 120232 304448 120284
rect 304500 120272 304506 120284
rect 307570 120272 307576 120284
rect 304500 120244 307576 120272
rect 304500 120232 304506 120244
rect 307570 120232 307576 120244
rect 307628 120232 307634 120284
rect 178862 120164 178868 120216
rect 178920 120204 178926 120216
rect 213914 120204 213920 120216
rect 178920 120176 213920 120204
rect 178920 120164 178926 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 276658 120164 276664 120216
rect 276716 120204 276722 120216
rect 307662 120204 307668 120216
rect 276716 120176 307668 120204
rect 276716 120164 276722 120176
rect 307662 120164 307668 120176
rect 307720 120164 307726 120216
rect 174722 120096 174728 120148
rect 174780 120136 174786 120148
rect 214006 120136 214012 120148
rect 174780 120108 214012 120136
rect 174780 120096 174786 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 253290 120096 253296 120148
rect 253348 120136 253354 120148
rect 307478 120136 307484 120148
rect 253348 120108 307484 120136
rect 253348 120096 253354 120108
rect 307478 120096 307484 120108
rect 307536 120096 307542 120148
rect 252462 120028 252468 120080
rect 252520 120068 252526 120080
rect 293402 120068 293408 120080
rect 252520 120040 293408 120068
rect 252520 120028 252526 120040
rect 293402 120028 293408 120040
rect 293460 120028 293466 120080
rect 496814 119620 496820 119672
rect 496872 119660 496878 119672
rect 499574 119660 499580 119672
rect 496872 119632 499580 119660
rect 496872 119620 496878 119632
rect 499574 119620 499580 119632
rect 499632 119620 499638 119672
rect 252370 119552 252376 119604
rect 252428 119592 252434 119604
rect 258810 119592 258816 119604
rect 252428 119564 258816 119592
rect 252428 119552 252434 119564
rect 258810 119552 258816 119564
rect 258868 119552 258874 119604
rect 170674 118804 170680 118856
rect 170732 118844 170738 118856
rect 214006 118844 214012 118856
rect 170732 118816 214012 118844
rect 170732 118804 170738 118816
rect 214006 118804 214012 118816
rect 214064 118804 214070 118856
rect 172054 118736 172060 118788
rect 172112 118776 172118 118788
rect 213914 118776 213920 118788
rect 172112 118748 213920 118776
rect 172112 118736 172118 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 300394 118736 300400 118788
rect 300452 118776 300458 118788
rect 307662 118776 307668 118788
rect 300452 118748 307668 118776
rect 300452 118736 300458 118748
rect 307662 118736 307668 118748
rect 307720 118736 307726 118788
rect 251910 118668 251916 118720
rect 251968 118708 251974 118720
rect 254854 118708 254860 118720
rect 251968 118680 254860 118708
rect 251968 118668 251974 118680
rect 254854 118668 254860 118680
rect 254912 118668 254918 118720
rect 293218 118668 293224 118720
rect 293276 118708 293282 118720
rect 307570 118708 307576 118720
rect 293276 118680 307576 118708
rect 293276 118668 293282 118680
rect 307570 118668 307576 118680
rect 307628 118668 307634 118720
rect 252462 118600 252468 118652
rect 252520 118640 252526 118652
rect 287882 118640 287888 118652
rect 252520 118612 287888 118640
rect 252520 118600 252526 118612
rect 287882 118600 287888 118612
rect 287940 118600 287946 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 345198 118640 345204 118652
rect 324464 118612 345204 118640
rect 324464 118600 324470 118612
rect 345198 118600 345204 118612
rect 345256 118600 345262 118652
rect 252370 118532 252376 118584
rect 252428 118572 252434 118584
rect 266998 118572 267004 118584
rect 252428 118544 267004 118572
rect 252428 118532 252434 118544
rect 266998 118532 267004 118544
rect 267056 118532 267062 118584
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 343818 118572 343824 118584
rect 324372 118544 343824 118572
rect 324372 118532 324378 118544
rect 343818 118532 343824 118544
rect 343876 118532 343882 118584
rect 496814 118396 496820 118448
rect 496872 118436 496878 118448
rect 501138 118436 501144 118448
rect 496872 118408 501144 118436
rect 496872 118396 496878 118408
rect 501138 118396 501144 118408
rect 501196 118396 501202 118448
rect 171778 117920 171784 117972
rect 171836 117960 171842 117972
rect 209130 117960 209136 117972
rect 171836 117932 209136 117960
rect 171836 117920 171842 117932
rect 209130 117920 209136 117932
rect 209188 117920 209194 117972
rect 252002 117920 252008 117972
rect 252060 117960 252066 117972
rect 300302 117960 300308 117972
rect 252060 117932 300308 117960
rect 252060 117920 252066 117932
rect 300302 117920 300308 117932
rect 300360 117920 300366 117972
rect 496814 117648 496820 117700
rect 496872 117688 496878 117700
rect 500954 117688 500960 117700
rect 496872 117660 500960 117688
rect 496872 117648 496878 117660
rect 500954 117648 500960 117660
rect 501012 117648 501018 117700
rect 287790 117512 287796 117564
rect 287848 117552 287854 117564
rect 306742 117552 306748 117564
rect 287848 117524 306748 117552
rect 287848 117512 287854 117524
rect 306742 117512 306748 117524
rect 306800 117512 306806 117564
rect 301682 117444 301688 117496
rect 301740 117484 301746 117496
rect 307570 117484 307576 117496
rect 301740 117456 307576 117484
rect 301740 117444 301746 117456
rect 307570 117444 307576 117456
rect 307628 117444 307634 117496
rect 173434 117376 173440 117428
rect 173492 117416 173498 117428
rect 214006 117416 214012 117428
rect 173492 117388 214012 117416
rect 173492 117376 173498 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 292114 117376 292120 117428
rect 292172 117416 292178 117428
rect 307478 117416 307484 117428
rect 292172 117388 307484 117416
rect 292172 117376 292178 117388
rect 307478 117376 307484 117388
rect 307536 117376 307542 117428
rect 169110 117308 169116 117360
rect 169168 117348 169174 117360
rect 213914 117348 213920 117360
rect 169168 117320 213920 117348
rect 169168 117308 169174 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 304258 117308 304264 117360
rect 304316 117348 304322 117360
rect 307662 117348 307668 117360
rect 304316 117320 307668 117348
rect 304316 117308 304322 117320
rect 307662 117308 307668 117320
rect 307720 117308 307726 117360
rect 252278 117240 252284 117292
rect 252336 117280 252342 117292
rect 285030 117280 285036 117292
rect 252336 117252 285036 117280
rect 252336 117240 252342 117252
rect 285030 117240 285036 117252
rect 285088 117240 285094 117292
rect 324406 117240 324412 117292
rect 324464 117280 324470 117292
rect 334066 117280 334072 117292
rect 324464 117252 334072 117280
rect 324464 117240 324470 117252
rect 334066 117240 334072 117252
rect 334124 117240 334130 117292
rect 342898 117240 342904 117292
rect 342956 117280 342962 117292
rect 416774 117280 416780 117292
rect 342956 117252 416780 117280
rect 342956 117240 342962 117252
rect 416774 117240 416780 117252
rect 416832 117240 416838 117292
rect 496906 117240 496912 117292
rect 496964 117280 496970 117292
rect 510706 117280 510712 117292
rect 496964 117252 510712 117280
rect 496964 117240 496970 117252
rect 510706 117240 510712 117252
rect 510764 117240 510770 117292
rect 252462 117172 252468 117224
rect 252520 117212 252526 117224
rect 272794 117212 272800 117224
rect 252520 117184 272800 117212
rect 252520 117172 252526 117184
rect 272794 117172 272800 117184
rect 272852 117172 272858 117224
rect 324314 117172 324320 117224
rect 324372 117212 324378 117224
rect 345106 117212 345112 117224
rect 324372 117184 345112 117212
rect 324372 117172 324378 117184
rect 345106 117172 345112 117184
rect 345164 117172 345170 117224
rect 252370 117104 252376 117156
rect 252428 117144 252434 117156
rect 260190 117144 260196 117156
rect 252428 117116 260196 117144
rect 252428 117104 252434 117116
rect 260190 117104 260196 117116
rect 260248 117104 260254 117156
rect 301498 116084 301504 116136
rect 301556 116124 301562 116136
rect 307478 116124 307484 116136
rect 301556 116096 307484 116124
rect 301556 116084 301562 116096
rect 307478 116084 307484 116096
rect 307536 116084 307542 116136
rect 198274 116016 198280 116068
rect 198332 116056 198338 116068
rect 214006 116056 214012 116068
rect 198332 116028 214012 116056
rect 198332 116016 198338 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 272518 116016 272524 116068
rect 272576 116056 272582 116068
rect 307570 116056 307576 116068
rect 272576 116028 307576 116056
rect 272576 116016 272582 116028
rect 307570 116016 307576 116028
rect 307628 116016 307634 116068
rect 192570 115948 192576 116000
rect 192628 115988 192634 116000
rect 213914 115988 213920 116000
rect 192628 115960 213920 115988
rect 192628 115948 192634 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 269850 115948 269856 116000
rect 269908 115988 269914 116000
rect 307662 115988 307668 116000
rect 269908 115960 307668 115988
rect 269908 115948 269914 115960
rect 307662 115948 307668 115960
rect 307720 115948 307726 116000
rect 252462 115880 252468 115932
rect 252520 115920 252526 115932
rect 272702 115920 272708 115932
rect 252520 115892 272708 115920
rect 252520 115880 252526 115892
rect 272702 115880 272708 115892
rect 272760 115880 272766 115932
rect 324314 115880 324320 115932
rect 324372 115920 324378 115932
rect 339494 115920 339500 115932
rect 324372 115892 339500 115920
rect 324372 115880 324378 115892
rect 339494 115880 339500 115892
rect 339552 115880 339558 115932
rect 252370 115812 252376 115864
rect 252428 115852 252434 115864
rect 262858 115852 262864 115864
rect 252428 115824 262864 115852
rect 252428 115812 252434 115824
rect 262858 115812 262864 115824
rect 262916 115812 262922 115864
rect 324406 115812 324412 115864
rect 324464 115852 324470 115864
rect 336734 115852 336740 115864
rect 324464 115824 336740 115852
rect 324464 115812 324470 115824
rect 336734 115812 336740 115824
rect 336792 115812 336798 115864
rect 196802 114588 196808 114640
rect 196860 114628 196866 114640
rect 214006 114628 214012 114640
rect 196860 114600 214012 114628
rect 196860 114588 196866 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 296254 114588 296260 114640
rect 296312 114628 296318 114640
rect 307570 114628 307576 114640
rect 296312 114600 307576 114628
rect 296312 114588 296318 114600
rect 307570 114588 307576 114600
rect 307628 114588 307634 114640
rect 177574 114520 177580 114572
rect 177632 114560 177638 114572
rect 213914 114560 213920 114572
rect 177632 114532 213920 114560
rect 177632 114520 177638 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 278130 114520 278136 114572
rect 278188 114560 278194 114572
rect 307662 114560 307668 114572
rect 278188 114532 307668 114560
rect 278188 114520 278194 114532
rect 307662 114520 307668 114532
rect 307720 114520 307726 114572
rect 252278 114452 252284 114504
rect 252336 114492 252342 114504
rect 298738 114492 298744 114504
rect 252336 114464 298744 114492
rect 252336 114452 252342 114464
rect 298738 114452 298744 114464
rect 298796 114452 298802 114504
rect 324314 114452 324320 114504
rect 324372 114492 324378 114504
rect 340966 114492 340972 114504
rect 324372 114464 340972 114492
rect 324372 114452 324378 114464
rect 340966 114452 340972 114464
rect 341024 114452 341030 114504
rect 252462 114384 252468 114436
rect 252520 114424 252526 114436
rect 267090 114424 267096 114436
rect 252520 114396 267096 114424
rect 252520 114384 252526 114396
rect 267090 114384 267096 114396
rect 267148 114384 267154 114436
rect 324406 114384 324412 114436
rect 324464 114424 324470 114436
rect 336826 114424 336832 114436
rect 324464 114396 336832 114424
rect 324464 114384 324470 114396
rect 336826 114384 336832 114396
rect 336884 114384 336890 114436
rect 252370 114316 252376 114368
rect 252428 114356 252434 114368
rect 261754 114356 261760 114368
rect 252428 114328 261760 114356
rect 252428 114316 252434 114328
rect 261754 114316 261760 114328
rect 261812 114316 261818 114368
rect 251818 113772 251824 113824
rect 251876 113812 251882 113824
rect 254762 113812 254768 113824
rect 251876 113784 254768 113812
rect 251876 113772 251882 113784
rect 254762 113772 254768 113784
rect 254820 113772 254826 113824
rect 300302 113296 300308 113348
rect 300360 113336 300366 113348
rect 307662 113336 307668 113348
rect 300360 113308 307668 113336
rect 300360 113296 300366 113308
rect 307662 113296 307668 113308
rect 307720 113296 307726 113348
rect 196894 113228 196900 113280
rect 196952 113268 196958 113280
rect 213914 113268 213920 113280
rect 196952 113240 213920 113268
rect 196952 113228 196958 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 266998 113228 267004 113280
rect 267056 113268 267062 113280
rect 306742 113268 306748 113280
rect 267056 113240 306748 113268
rect 267056 113228 267062 113240
rect 306742 113228 306748 113240
rect 306800 113228 306806 113280
rect 169294 113160 169300 113212
rect 169352 113200 169358 113212
rect 214006 113200 214012 113212
rect 169352 113172 214012 113200
rect 169352 113160 169358 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 261478 113160 261484 113212
rect 261536 113200 261542 113212
rect 307570 113200 307576 113212
rect 261536 113172 307576 113200
rect 261536 113160 261542 113172
rect 307570 113160 307576 113172
rect 307628 113160 307634 113212
rect 252462 113092 252468 113144
rect 252520 113132 252526 113144
rect 302970 113132 302976 113144
rect 252520 113104 302976 113132
rect 252520 113092 252526 113104
rect 302970 113092 302976 113104
rect 303028 113092 303034 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 335354 113132 335360 113144
rect 324372 113104 335360 113132
rect 324372 113092 324378 113104
rect 335354 113092 335360 113104
rect 335412 113092 335418 113144
rect 349246 113092 349252 113144
rect 349304 113132 349310 113144
rect 367738 113132 367744 113144
rect 349304 113104 367744 113132
rect 349304 113092 349310 113104
rect 367738 113092 367744 113104
rect 367796 113092 367802 113144
rect 395338 113092 395344 113144
rect 395396 113132 395402 113144
rect 416774 113132 416780 113144
rect 395396 113104 416780 113132
rect 395396 113092 395402 113104
rect 416774 113092 416780 113104
rect 416832 113092 416838 113144
rect 252370 113024 252376 113076
rect 252428 113064 252434 113076
rect 276842 113064 276848 113076
rect 252428 113036 276848 113064
rect 252428 113024 252434 113036
rect 276842 113024 276848 113036
rect 276900 113024 276906 113076
rect 252462 112888 252468 112940
rect 252520 112928 252526 112940
rect 256142 112928 256148 112940
rect 252520 112900 256148 112928
rect 252520 112888 252526 112900
rect 256142 112888 256148 112900
rect 256200 112888 256206 112940
rect 322934 112412 322940 112464
rect 322992 112452 322998 112464
rect 349246 112452 349252 112464
rect 322992 112424 349252 112452
rect 322992 112412 322998 112424
rect 349246 112412 349252 112424
rect 349304 112412 349310 112464
rect 200942 111868 200948 111920
rect 201000 111908 201006 111920
rect 213914 111908 213920 111920
rect 201000 111880 213920 111908
rect 201000 111868 201006 111880
rect 213914 111868 213920 111880
rect 213972 111868 213978 111920
rect 286410 111868 286416 111920
rect 286468 111908 286474 111920
rect 307570 111908 307576 111920
rect 286468 111880 307576 111908
rect 286468 111868 286474 111880
rect 307570 111868 307576 111880
rect 307628 111868 307634 111920
rect 174814 111800 174820 111852
rect 174872 111840 174878 111852
rect 214006 111840 214012 111852
rect 174872 111812 214012 111840
rect 174872 111800 174878 111812
rect 214006 111800 214012 111812
rect 214064 111800 214070 111852
rect 276750 111800 276756 111852
rect 276808 111840 276814 111852
rect 307662 111840 307668 111852
rect 276808 111812 307668 111840
rect 276808 111800 276814 111812
rect 307662 111800 307668 111812
rect 307720 111800 307726 111852
rect 496906 111800 496912 111852
rect 496964 111840 496970 111852
rect 499574 111840 499580 111852
rect 496964 111812 499580 111840
rect 496964 111800 496970 111812
rect 499574 111800 499580 111812
rect 499632 111800 499638 111852
rect 167914 111732 167920 111784
rect 167972 111772 167978 111784
rect 196710 111772 196716 111784
rect 167972 111744 196716 111772
rect 167972 111732 167978 111744
rect 196710 111732 196716 111744
rect 196768 111732 196774 111784
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 308490 111772 308496 111784
rect 252520 111744 308496 111772
rect 252520 111732 252526 111744
rect 308490 111732 308496 111744
rect 308548 111732 308554 111784
rect 371878 111732 371884 111784
rect 371936 111772 371942 111784
rect 416774 111772 416780 111784
rect 371936 111744 416780 111772
rect 371936 111732 371942 111744
rect 416774 111732 416780 111744
rect 416832 111732 416838 111784
rect 496814 111732 496820 111784
rect 496872 111772 496878 111784
rect 506474 111772 506480 111784
rect 496872 111744 506480 111772
rect 496872 111732 496878 111744
rect 506474 111732 506480 111744
rect 506532 111732 506538 111784
rect 252370 111664 252376 111716
rect 252428 111704 252434 111716
rect 257614 111704 257620 111716
rect 252428 111676 257620 111704
rect 252428 111664 252434 111676
rect 257614 111664 257620 111676
rect 257672 111664 257678 111716
rect 3418 110984 3424 111036
rect 3476 111024 3482 111036
rect 7558 111024 7564 111036
rect 3476 110996 7564 111024
rect 3476 110984 3482 110996
rect 7558 110984 7564 110996
rect 7616 110984 7622 111036
rect 252462 110644 252468 110696
rect 252520 110684 252526 110696
rect 258718 110684 258724 110696
rect 252520 110656 258724 110684
rect 252520 110644 252526 110656
rect 258718 110644 258724 110656
rect 258776 110644 258782 110696
rect 289354 110576 289360 110628
rect 289412 110616 289418 110628
rect 307478 110616 307484 110628
rect 289412 110588 307484 110616
rect 289412 110576 289418 110588
rect 307478 110576 307484 110588
rect 307536 110576 307542 110628
rect 173342 110508 173348 110560
rect 173400 110548 173406 110560
rect 213914 110548 213920 110560
rect 173400 110520 213920 110548
rect 173400 110508 173406 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 257430 110508 257436 110560
rect 257488 110548 257494 110560
rect 307570 110548 307576 110560
rect 257488 110520 307576 110548
rect 257488 110508 257494 110520
rect 307570 110508 307576 110520
rect 307628 110508 307634 110560
rect 166350 110440 166356 110492
rect 166408 110480 166414 110492
rect 214006 110480 214012 110492
rect 166408 110452 214012 110480
rect 166408 110440 166414 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 250438 110440 250444 110492
rect 250496 110480 250502 110492
rect 307662 110480 307668 110492
rect 250496 110452 307668 110480
rect 250496 110440 250502 110452
rect 307662 110440 307668 110452
rect 307720 110440 307726 110492
rect 252278 110372 252284 110424
rect 252336 110412 252342 110424
rect 303062 110412 303068 110424
rect 252336 110384 303068 110412
rect 252336 110372 252342 110384
rect 303062 110372 303068 110384
rect 303120 110372 303126 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 332870 110412 332876 110424
rect 324372 110384 332876 110412
rect 324372 110372 324378 110384
rect 332870 110372 332876 110384
rect 332928 110372 332934 110424
rect 377398 110372 377404 110424
rect 377456 110412 377462 110424
rect 416774 110412 416780 110424
rect 377456 110384 416780 110412
rect 377456 110372 377462 110384
rect 416774 110372 416780 110384
rect 416832 110372 416838 110424
rect 496814 110372 496820 110424
rect 496872 110412 496878 110424
rect 510614 110412 510620 110424
rect 496872 110384 510620 110412
rect 496872 110372 496878 110384
rect 510614 110372 510620 110384
rect 510672 110372 510678 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 289262 110344 289268 110356
rect 252520 110316 289268 110344
rect 252520 110304 252526 110316
rect 289262 110304 289268 110316
rect 289320 110304 289326 110356
rect 252370 110236 252376 110288
rect 252428 110276 252434 110288
rect 264238 110276 264244 110288
rect 252428 110248 264244 110276
rect 252428 110236 252434 110248
rect 264238 110236 264244 110248
rect 264296 110236 264302 110288
rect 324406 109692 324412 109744
rect 324464 109732 324470 109744
rect 329834 109732 329840 109744
rect 324464 109704 329840 109732
rect 324464 109692 324470 109704
rect 329834 109692 329840 109704
rect 329892 109692 329898 109744
rect 302970 109148 302976 109200
rect 303028 109188 303034 109200
rect 306742 109188 306748 109200
rect 303028 109160 306748 109188
rect 303028 109148 303034 109160
rect 306742 109148 306748 109160
rect 306800 109148 306806 109200
rect 178954 109080 178960 109132
rect 179012 109120 179018 109132
rect 213914 109120 213920 109132
rect 179012 109092 213920 109120
rect 179012 109080 179018 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 294690 109080 294696 109132
rect 294748 109120 294754 109132
rect 307570 109120 307576 109132
rect 294748 109092 307576 109120
rect 294748 109080 294754 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 166442 109012 166448 109064
rect 166500 109052 166506 109064
rect 214006 109052 214012 109064
rect 166500 109024 214012 109052
rect 166500 109012 166506 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 285030 109012 285036 109064
rect 285088 109052 285094 109064
rect 307662 109052 307668 109064
rect 285088 109024 307668 109052
rect 285088 109012 285094 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 252278 108944 252284 108996
rect 252336 108984 252342 108996
rect 287974 108984 287980 108996
rect 252336 108956 287980 108984
rect 252336 108944 252342 108956
rect 287974 108944 287980 108956
rect 288032 108944 288038 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 279510 108916 279516 108928
rect 252520 108888 279516 108916
rect 252520 108876 252526 108888
rect 279510 108876 279516 108888
rect 279568 108876 279574 108928
rect 252370 108808 252376 108860
rect 252428 108848 252434 108860
rect 265710 108848 265716 108860
rect 252428 108820 265716 108848
rect 252428 108808 252434 108820
rect 265710 108808 265716 108820
rect 265768 108808 265774 108860
rect 324314 108740 324320 108792
rect 324372 108780 324378 108792
rect 327166 108780 327172 108792
rect 324372 108752 327172 108780
rect 324372 108740 324378 108752
rect 327166 108740 327172 108752
rect 327224 108740 327230 108792
rect 282362 107856 282368 107908
rect 282420 107896 282426 107908
rect 307478 107896 307484 107908
rect 282420 107868 307484 107896
rect 282420 107856 282426 107868
rect 307478 107856 307484 107868
rect 307536 107856 307542 107908
rect 169202 107720 169208 107772
rect 169260 107760 169266 107772
rect 213914 107760 213920 107772
rect 169260 107732 213920 107760
rect 169260 107720 169266 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 287882 107720 287888 107772
rect 287940 107760 287946 107772
rect 307662 107760 307668 107772
rect 287940 107732 307668 107760
rect 287940 107720 287946 107732
rect 307662 107720 307668 107732
rect 307720 107720 307726 107772
rect 167914 107652 167920 107704
rect 167972 107692 167978 107704
rect 214006 107692 214012 107704
rect 167972 107664 214012 107692
rect 167972 107652 167978 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 303062 107652 303068 107704
rect 303120 107692 303126 107704
rect 306926 107692 306932 107704
rect 303120 107664 306932 107692
rect 303120 107652 303126 107664
rect 306926 107652 306932 107664
rect 306984 107652 306990 107704
rect 252462 107584 252468 107636
rect 252520 107624 252526 107636
rect 286594 107624 286600 107636
rect 252520 107596 286600 107624
rect 252520 107584 252526 107596
rect 286594 107584 286600 107596
rect 286652 107584 286658 107636
rect 324314 107584 324320 107636
rect 324372 107624 324378 107636
rect 340874 107624 340880 107636
rect 324372 107596 340880 107624
rect 324372 107584 324378 107596
rect 340874 107584 340880 107596
rect 340932 107584 340938 107636
rect 403710 107584 403716 107636
rect 403768 107624 403774 107636
rect 416774 107624 416780 107636
rect 403768 107596 416780 107624
rect 403768 107584 403774 107596
rect 416774 107584 416780 107596
rect 416832 107584 416838 107636
rect 252370 107516 252376 107568
rect 252428 107556 252434 107568
rect 257338 107556 257344 107568
rect 252428 107528 257344 107556
rect 252428 107516 252434 107528
rect 257338 107516 257344 107528
rect 257396 107516 257402 107568
rect 290550 106428 290556 106480
rect 290608 106468 290614 106480
rect 307570 106468 307576 106480
rect 290608 106440 307576 106468
rect 290608 106428 290614 106440
rect 307570 106428 307576 106440
rect 307628 106428 307634 106480
rect 181622 106360 181628 106412
rect 181680 106400 181686 106412
rect 213914 106400 213920 106412
rect 181680 106372 213920 106400
rect 181680 106360 181686 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 269758 106360 269764 106412
rect 269816 106400 269822 106412
rect 307478 106400 307484 106412
rect 269816 106372 307484 106400
rect 269816 106360 269822 106372
rect 307478 106360 307484 106372
rect 307536 106360 307542 106412
rect 169018 106292 169024 106344
rect 169076 106332 169082 106344
rect 214006 106332 214012 106344
rect 169076 106304 214012 106332
rect 169076 106292 169082 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 249058 106292 249064 106344
rect 249116 106332 249122 106344
rect 307662 106332 307668 106344
rect 249116 106304 307668 106332
rect 249116 106292 249122 106304
rect 307662 106292 307668 106304
rect 307720 106292 307726 106344
rect 252462 106224 252468 106276
rect 252520 106264 252526 106276
rect 255958 106264 255964 106276
rect 252520 106236 255964 106264
rect 252520 106224 252526 106236
rect 255958 106224 255964 106236
rect 256016 106224 256022 106276
rect 341518 106224 341524 106276
rect 341576 106264 341582 106276
rect 416774 106264 416780 106276
rect 341576 106236 416780 106264
rect 341576 106224 341582 106236
rect 416774 106224 416780 106236
rect 416832 106224 416838 106276
rect 496814 106224 496820 106276
rect 496872 106264 496878 106276
rect 507946 106264 507952 106276
rect 496872 106236 507952 106264
rect 496872 106224 496878 106236
rect 507946 106224 507952 106236
rect 508004 106224 508010 106276
rect 252186 105612 252192 105664
rect 252244 105652 252250 105664
rect 283742 105652 283748 105664
rect 252244 105624 283748 105652
rect 252244 105612 252250 105624
rect 283742 105612 283748 105624
rect 283800 105612 283806 105664
rect 252278 105544 252284 105596
rect 252336 105584 252342 105596
rect 296162 105584 296168 105596
rect 252336 105556 296168 105584
rect 252336 105544 252342 105556
rect 296162 105544 296168 105556
rect 296220 105544 296226 105596
rect 300210 105000 300216 105052
rect 300268 105040 300274 105052
rect 307478 105040 307484 105052
rect 300268 105012 307484 105040
rect 300268 105000 300274 105012
rect 307478 105000 307484 105012
rect 307536 105000 307542 105052
rect 283650 104932 283656 104984
rect 283708 104972 283714 104984
rect 307570 104972 307576 104984
rect 283708 104944 307576 104972
rect 283708 104932 283714 104944
rect 307570 104932 307576 104944
rect 307628 104932 307634 104984
rect 202414 104864 202420 104916
rect 202472 104904 202478 104916
rect 213914 104904 213920 104916
rect 202472 104876 213920 104904
rect 202472 104864 202478 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 264330 104864 264336 104916
rect 264388 104904 264394 104916
rect 307662 104904 307668 104916
rect 264388 104876 307668 104904
rect 264388 104864 264394 104876
rect 307662 104864 307668 104876
rect 307720 104864 307726 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 269942 104836 269948 104848
rect 252520 104808 269948 104836
rect 252520 104796 252526 104808
rect 269942 104796 269948 104808
rect 270000 104796 270006 104848
rect 359458 104796 359464 104848
rect 359516 104836 359522 104848
rect 416774 104836 416780 104848
rect 359516 104808 416780 104836
rect 359516 104796 359522 104808
rect 416774 104796 416780 104808
rect 416832 104796 416838 104848
rect 252370 104728 252376 104780
rect 252428 104768 252434 104780
rect 264514 104768 264520 104780
rect 252428 104740 264520 104768
rect 252428 104728 252434 104740
rect 264514 104728 264520 104740
rect 264572 104728 264578 104780
rect 267090 103640 267096 103692
rect 267148 103680 267154 103692
rect 306742 103680 306748 103692
rect 267148 103652 306748 103680
rect 267148 103640 267154 103652
rect 306742 103640 306748 103652
rect 306800 103640 306806 103692
rect 264238 103572 264244 103624
rect 264296 103612 264302 103624
rect 307570 103612 307576 103624
rect 264296 103584 307576 103612
rect 264296 103572 264302 103584
rect 307570 103572 307576 103584
rect 307628 103572 307634 103624
rect 188430 103504 188436 103556
rect 188488 103544 188494 103556
rect 213914 103544 213920 103556
rect 188488 103516 213920 103544
rect 188488 103504 188494 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 264422 103504 264428 103556
rect 264480 103544 264486 103556
rect 307662 103544 307668 103556
rect 264480 103516 307668 103544
rect 264480 103504 264486 103516
rect 307662 103504 307668 103516
rect 307720 103504 307726 103556
rect 407758 103436 407764 103488
rect 407816 103476 407822 103488
rect 416774 103476 416780 103488
rect 407816 103448 416780 103476
rect 407816 103436 407822 103448
rect 416774 103436 416780 103448
rect 416832 103436 416838 103488
rect 252462 103368 252468 103420
rect 252520 103408 252526 103420
rect 275278 103408 275284 103420
rect 252520 103380 275284 103408
rect 252520 103368 252526 103380
rect 275278 103368 275284 103380
rect 275336 103368 275342 103420
rect 252370 103300 252376 103352
rect 252428 103340 252434 103352
rect 280890 103340 280896 103352
rect 252428 103312 280896 103340
rect 252428 103300 252434 103312
rect 280890 103300 280896 103312
rect 280948 103300 280954 103352
rect 251174 102892 251180 102944
rect 251232 102932 251238 102944
rect 253382 102932 253388 102944
rect 251232 102904 253388 102932
rect 251232 102892 251238 102904
rect 253382 102892 253388 102904
rect 253440 102892 253446 102944
rect 330478 102756 330484 102808
rect 330536 102796 330542 102808
rect 376018 102796 376024 102808
rect 330536 102768 376024 102796
rect 330536 102756 330542 102768
rect 376018 102756 376024 102768
rect 376076 102756 376082 102808
rect 296162 102280 296168 102332
rect 296220 102320 296226 102332
rect 306742 102320 306748 102332
rect 296220 102292 306748 102320
rect 296220 102280 296226 102292
rect 306742 102280 306748 102292
rect 306800 102280 306806 102332
rect 207842 102212 207848 102264
rect 207900 102252 207906 102264
rect 213914 102252 213920 102264
rect 207900 102224 213920 102252
rect 207900 102212 207906 102224
rect 213914 102212 213920 102224
rect 213972 102212 213978 102264
rect 280982 102212 280988 102264
rect 281040 102252 281046 102264
rect 307662 102252 307668 102264
rect 281040 102224 307668 102252
rect 281040 102212 281046 102224
rect 307662 102212 307668 102224
rect 307720 102212 307726 102264
rect 192662 102144 192668 102196
rect 192720 102184 192726 102196
rect 214006 102184 214012 102196
rect 192720 102156 214012 102184
rect 192720 102144 192726 102156
rect 214006 102144 214012 102156
rect 214064 102144 214070 102196
rect 262858 102144 262864 102196
rect 262916 102184 262922 102196
rect 307570 102184 307576 102196
rect 262916 102156 307576 102184
rect 262916 102144 262922 102156
rect 307570 102144 307576 102156
rect 307628 102144 307634 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 276934 102116 276940 102128
rect 252520 102088 276940 102116
rect 252520 102076 252526 102088
rect 276934 102076 276940 102088
rect 276992 102076 276998 102128
rect 252186 101396 252192 101448
rect 252244 101436 252250 101448
rect 256050 101436 256056 101448
rect 252244 101408 256056 101436
rect 252244 101396 252250 101408
rect 256050 101396 256056 101408
rect 256108 101396 256114 101448
rect 298738 100852 298744 100904
rect 298796 100892 298802 100904
rect 307570 100892 307576 100904
rect 298796 100864 307576 100892
rect 298796 100852 298802 100864
rect 307570 100852 307576 100864
rect 307628 100852 307634 100904
rect 206554 100784 206560 100836
rect 206612 100824 206618 100836
rect 214006 100824 214012 100836
rect 206612 100796 214012 100824
rect 206612 100784 206618 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 260190 100784 260196 100836
rect 260248 100824 260254 100836
rect 307662 100824 307668 100836
rect 260248 100796 307668 100824
rect 260248 100784 260254 100796
rect 307662 100784 307668 100796
rect 307720 100784 307726 100836
rect 200850 100716 200856 100768
rect 200908 100756 200914 100768
rect 213914 100756 213920 100768
rect 200908 100728 213920 100756
rect 200908 100716 200914 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 258718 100716 258724 100768
rect 258776 100756 258782 100768
rect 306926 100756 306932 100768
rect 258776 100728 306932 100756
rect 258776 100716 258782 100728
rect 306926 100716 306932 100728
rect 306984 100716 306990 100768
rect 252370 100648 252376 100700
rect 252428 100688 252434 100700
rect 290642 100688 290648 100700
rect 252428 100660 290648 100688
rect 252428 100648 252434 100660
rect 290642 100648 290648 100660
rect 290700 100648 290706 100700
rect 360194 100648 360200 100700
rect 360252 100688 360258 100700
rect 370498 100688 370504 100700
rect 360252 100660 370504 100688
rect 360252 100648 360258 100660
rect 370498 100648 370504 100660
rect 370556 100648 370562 100700
rect 378778 100648 378784 100700
rect 378836 100688 378842 100700
rect 494054 100688 494060 100700
rect 378836 100660 494060 100688
rect 378836 100648 378842 100660
rect 494054 100648 494060 100660
rect 494112 100648 494118 100700
rect 519538 100648 519544 100700
rect 519596 100688 519602 100700
rect 580166 100688 580172 100700
rect 519596 100660 580172 100688
rect 519596 100648 519602 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 270034 100620 270040 100632
rect 252520 100592 270040 100620
rect 252520 100580 252526 100592
rect 270034 100580 270040 100592
rect 270092 100580 270098 100632
rect 406378 100580 406384 100632
rect 406436 100620 406442 100632
rect 496814 100620 496820 100632
rect 406436 100592 496820 100620
rect 406436 100580 406442 100592
rect 496814 100580 496820 100592
rect 496872 100580 496878 100632
rect 252278 100512 252284 100564
rect 252336 100552 252342 100564
rect 260466 100552 260472 100564
rect 252336 100524 260472 100552
rect 252336 100512 252342 100524
rect 260466 100512 260472 100524
rect 260524 100512 260530 100564
rect 167730 99968 167736 100020
rect 167788 100008 167794 100020
rect 214558 100008 214564 100020
rect 167788 99980 214564 100008
rect 167788 99968 167794 99980
rect 214558 99968 214564 99980
rect 214616 99968 214622 100020
rect 325694 99968 325700 100020
rect 325752 100008 325758 100020
rect 360194 100008 360200 100020
rect 325752 99980 360200 100008
rect 325752 99968 325758 99980
rect 360194 99968 360200 99980
rect 360252 99968 360258 100020
rect 254762 99492 254768 99544
rect 254820 99532 254826 99544
rect 307570 99532 307576 99544
rect 254820 99504 307576 99532
rect 254820 99492 254826 99504
rect 307570 99492 307576 99504
rect 307628 99492 307634 99544
rect 275278 99424 275284 99476
rect 275336 99464 275342 99476
rect 307662 99464 307668 99476
rect 275336 99436 307668 99464
rect 275336 99424 275342 99436
rect 307662 99424 307668 99436
rect 307720 99424 307726 99476
rect 164878 99356 164884 99408
rect 164936 99396 164942 99408
rect 213914 99396 213920 99408
rect 164936 99368 213920 99396
rect 164936 99356 164942 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 252462 99288 252468 99340
rect 252520 99328 252526 99340
rect 261662 99328 261668 99340
rect 252520 99300 261668 99328
rect 252520 99288 252526 99300
rect 261662 99288 261668 99300
rect 261720 99288 261726 99340
rect 419626 99288 419632 99340
rect 419684 99328 419690 99340
rect 580258 99328 580264 99340
rect 419684 99300 580264 99328
rect 419684 99288 419690 99300
rect 580258 99288 580264 99300
rect 580316 99288 580322 99340
rect 251910 99220 251916 99272
rect 251968 99260 251974 99272
rect 254946 99260 254952 99272
rect 251968 99232 254952 99260
rect 251968 99220 251974 99232
rect 254946 99220 254952 99232
rect 255004 99220 255010 99272
rect 400858 99220 400864 99272
rect 400916 99260 400922 99272
rect 493962 99260 493968 99272
rect 400916 99232 493968 99260
rect 400916 99220 400922 99232
rect 493962 99220 493968 99232
rect 494020 99220 494026 99272
rect 410610 99152 410616 99204
rect 410668 99192 410674 99204
rect 496906 99192 496912 99204
rect 410668 99164 496912 99192
rect 410668 99152 410674 99164
rect 496906 99152 496912 99164
rect 496964 99152 496970 99204
rect 171778 98608 171784 98660
rect 171836 98648 171842 98660
rect 214006 98648 214012 98660
rect 171836 98620 214012 98648
rect 171836 98608 171842 98620
rect 214006 98608 214012 98620
rect 214064 98608 214070 98660
rect 324406 98608 324412 98660
rect 324464 98648 324470 98660
rect 331582 98648 331588 98660
rect 324464 98620 331588 98648
rect 324464 98608 324470 98620
rect 331582 98608 331588 98620
rect 331640 98608 331646 98660
rect 264514 98064 264520 98116
rect 264572 98104 264578 98116
rect 307662 98104 307668 98116
rect 264572 98076 307668 98104
rect 264572 98064 264578 98076
rect 307662 98064 307668 98076
rect 307720 98064 307726 98116
rect 212442 97996 212448 98048
rect 212500 98036 212506 98048
rect 213914 98036 213920 98048
rect 212500 98008 213920 98036
rect 212500 97996 212506 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 251910 97996 251916 98048
rect 251968 98036 251974 98048
rect 306742 98036 306748 98048
rect 251968 98008 306748 98036
rect 251968 97996 251974 98008
rect 306742 97996 306748 98008
rect 306800 97996 306806 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 17218 97968 17224 97980
rect 3476 97940 17224 97968
rect 3476 97928 3482 97940
rect 17218 97928 17224 97940
rect 17276 97928 17282 97980
rect 324314 97928 324320 97980
rect 324372 97968 324378 97980
rect 346394 97968 346400 97980
rect 324372 97940 346400 97968
rect 324372 97928 324378 97940
rect 346394 97928 346400 97940
rect 346452 97928 346458 97980
rect 399478 97928 399484 97980
rect 399536 97968 399542 97980
rect 494330 97968 494336 97980
rect 399536 97940 494336 97968
rect 399536 97928 399542 97940
rect 494330 97928 494336 97940
rect 494388 97928 494394 97980
rect 413278 97860 413284 97912
rect 413336 97900 413342 97912
rect 496998 97900 497004 97912
rect 413336 97872 497004 97900
rect 413336 97860 413342 97872
rect 496998 97860 497004 97872
rect 497056 97860 497062 97912
rect 420178 97316 420184 97368
rect 420236 97356 420242 97368
rect 427722 97356 427728 97368
rect 420236 97328 427728 97356
rect 420236 97316 420242 97328
rect 427722 97316 427728 97328
rect 427780 97316 427786 97368
rect 166534 97248 166540 97300
rect 166592 97288 166598 97300
rect 214650 97288 214656 97300
rect 166592 97260 214656 97288
rect 166592 97248 166598 97260
rect 214650 97248 214656 97260
rect 214708 97248 214714 97300
rect 252002 97248 252008 97300
rect 252060 97288 252066 97300
rect 259362 97288 259368 97300
rect 252060 97260 259368 97288
rect 252060 97248 252066 97260
rect 259362 97248 259368 97260
rect 259420 97288 259426 97300
rect 308398 97288 308404 97300
rect 259420 97260 308404 97288
rect 259420 97248 259426 97260
rect 308398 97248 308404 97260
rect 308456 97248 308462 97300
rect 421558 97248 421564 97300
rect 421616 97288 421622 97300
rect 458910 97288 458916 97300
rect 421616 97260 458916 97288
rect 421616 97248 421622 97260
rect 458910 97248 458916 97260
rect 458968 97248 458974 97300
rect 467098 97248 467104 97300
rect 467156 97288 467162 97300
rect 492490 97288 492496 97300
rect 467156 97260 492496 97288
rect 467156 97248 467162 97260
rect 492490 97248 492496 97260
rect 492548 97248 492554 97300
rect 439498 96908 439504 96960
rect 439556 96948 439562 96960
rect 440878 96948 440884 96960
rect 439556 96920 440884 96948
rect 439556 96908 439562 96920
rect 440878 96908 440884 96920
rect 440936 96908 440942 96960
rect 454034 96908 454040 96960
rect 454092 96948 454098 96960
rect 455046 96948 455052 96960
rect 454092 96920 455052 96948
rect 454092 96908 454098 96920
rect 455046 96908 455052 96920
rect 455104 96908 455110 96960
rect 461578 96908 461584 96960
rect 461636 96948 461642 96960
rect 464890 96948 464896 96960
rect 461636 96920 464896 96948
rect 461636 96908 461642 96920
rect 464890 96908 464896 96920
rect 464948 96908 464954 96960
rect 465718 96908 465724 96960
rect 465776 96948 465782 96960
rect 467282 96948 467288 96960
rect 465776 96920 467288 96948
rect 465776 96908 465782 96920
rect 467282 96908 467288 96920
rect 467340 96908 467346 96960
rect 472618 96908 472624 96960
rect 472676 96948 472682 96960
rect 474550 96948 474556 96960
rect 472676 96920 474556 96948
rect 472676 96908 472682 96920
rect 474550 96908 474556 96920
rect 474608 96908 474614 96960
rect 481634 96908 481640 96960
rect 481692 96948 481698 96960
rect 482646 96948 482652 96960
rect 481692 96920 482652 96948
rect 481692 96908 481698 96920
rect 482646 96908 482652 96920
rect 482704 96908 482710 96960
rect 486418 96908 486424 96960
rect 486476 96948 486482 96960
rect 487706 96948 487712 96960
rect 486476 96920 487712 96948
rect 486476 96908 486482 96920
rect 487706 96908 487712 96920
rect 487764 96908 487770 96960
rect 289262 96772 289268 96824
rect 289320 96812 289326 96824
rect 307662 96812 307668 96824
rect 289320 96784 307668 96812
rect 289320 96772 289326 96784
rect 307662 96772 307668 96784
rect 307720 96772 307726 96824
rect 417418 96772 417424 96824
rect 417476 96812 417482 96824
rect 420546 96812 420552 96824
rect 417476 96784 420552 96812
rect 417476 96772 417482 96784
rect 420546 96772 420552 96784
rect 420604 96772 420610 96824
rect 258810 96704 258816 96756
rect 258868 96744 258874 96756
rect 306926 96744 306932 96756
rect 258868 96716 306932 96744
rect 258868 96704 258874 96716
rect 306926 96704 306932 96716
rect 306984 96704 306990 96756
rect 253382 96636 253388 96688
rect 253440 96676 253446 96688
rect 307570 96676 307576 96688
rect 253440 96648 307576 96676
rect 253440 96636 253446 96648
rect 307570 96636 307576 96648
rect 307628 96636 307634 96688
rect 186222 96568 186228 96620
rect 186280 96608 186286 96620
rect 321462 96608 321468 96620
rect 186280 96580 321468 96608
rect 186280 96568 186286 96580
rect 321462 96568 321468 96580
rect 321520 96568 321526 96620
rect 350534 96568 350540 96620
rect 350592 96608 350598 96620
rect 351178 96608 351184 96620
rect 350592 96580 351184 96608
rect 350592 96568 350598 96580
rect 351178 96568 351184 96580
rect 351236 96608 351242 96620
rect 501046 96608 501052 96620
rect 351236 96580 501052 96608
rect 351236 96568 351242 96580
rect 501046 96568 501052 96580
rect 501104 96568 501110 96620
rect 282178 96500 282184 96552
rect 282236 96540 282242 96552
rect 321554 96540 321560 96552
rect 282236 96512 321560 96540
rect 282236 96500 282242 96512
rect 321554 96500 321560 96512
rect 321612 96500 321618 96552
rect 309778 96432 309784 96484
rect 309836 96472 309842 96484
rect 321646 96472 321652 96484
rect 309836 96444 321652 96472
rect 309836 96432 309842 96444
rect 321646 96432 321652 96444
rect 321704 96432 321710 96484
rect 203610 95208 203616 95260
rect 203668 95248 203674 95260
rect 213914 95248 213920 95260
rect 203668 95220 213920 95248
rect 203668 95208 203674 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 247678 95208 247684 95260
rect 247736 95248 247742 95260
rect 307662 95248 307668 95260
rect 247736 95220 307668 95248
rect 247736 95208 247742 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 203518 95140 203524 95192
rect 203576 95180 203582 95192
rect 321370 95180 321376 95192
rect 203576 95152 321376 95180
rect 203576 95140 203582 95152
rect 321370 95140 321376 95152
rect 321428 95140 321434 95192
rect 389818 95140 389824 95192
rect 389876 95180 389882 95192
rect 499574 95180 499580 95192
rect 389876 95152 499580 95180
rect 389876 95140 389882 95152
rect 499574 95140 499580 95152
rect 499632 95140 499638 95192
rect 204162 95072 204168 95124
rect 204220 95112 204226 95124
rect 321830 95112 321836 95124
rect 204220 95084 321836 95112
rect 204220 95072 204226 95084
rect 321830 95072 321836 95084
rect 321888 95072 321894 95124
rect 206278 95004 206284 95056
rect 206336 95044 206342 95056
rect 321738 95044 321744 95056
rect 206336 95016 321744 95044
rect 206336 95004 206342 95016
rect 321738 95004 321744 95016
rect 321796 95004 321802 95056
rect 290458 94936 290464 94988
rect 290516 94976 290522 94988
rect 323026 94976 323032 94988
rect 290516 94948 323032 94976
rect 290516 94936 290522 94948
rect 323026 94936 323032 94948
rect 323084 94936 323090 94988
rect 296070 94868 296076 94920
rect 296128 94908 296134 94920
rect 323210 94908 323216 94920
rect 296128 94880 323216 94908
rect 296128 94868 296134 94880
rect 323210 94868 323216 94880
rect 323268 94868 323274 94920
rect 304902 94800 304908 94852
rect 304960 94840 304966 94852
rect 324498 94840 324504 94852
rect 304960 94812 324504 94840
rect 304960 94800 304966 94812
rect 324498 94800 324504 94812
rect 324556 94800 324562 94852
rect 129550 94460 129556 94512
rect 129608 94500 129614 94512
rect 214006 94500 214012 94512
rect 129608 94472 214012 94500
rect 129608 94460 129614 94472
rect 214006 94460 214012 94472
rect 214064 94460 214070 94512
rect 333974 94460 333980 94512
rect 334032 94500 334038 94512
rect 494238 94500 494244 94512
rect 334032 94472 494244 94500
rect 334032 94460 334038 94472
rect 494238 94460 494244 94472
rect 494296 94460 494302 94512
rect 124490 94052 124496 94104
rect 124548 94092 124554 94104
rect 174630 94092 174636 94104
rect 124548 94064 174636 94092
rect 124548 94052 124554 94064
rect 174630 94052 174636 94064
rect 174688 94052 174694 94104
rect 112346 93984 112352 94036
rect 112404 94024 112410 94036
rect 172054 94024 172060 94036
rect 112404 93996 172060 94024
rect 112404 93984 112410 93996
rect 172054 93984 172060 93996
rect 172112 93984 172118 94036
rect 122834 93916 122840 93968
rect 122892 93956 122898 93968
rect 185670 93956 185676 93968
rect 122892 93928 185676 93956
rect 122892 93916 122898 93928
rect 185670 93916 185676 93928
rect 185728 93916 185734 93968
rect 85574 93848 85580 93900
rect 85632 93888 85638 93900
rect 212442 93888 212448 93900
rect 85632 93860 212448 93888
rect 85632 93848 85638 93860
rect 212442 93848 212448 93860
rect 212500 93848 212506 93900
rect 56502 93780 56508 93832
rect 56560 93820 56566 93832
rect 192662 93820 192668 93832
rect 56560 93792 192668 93820
rect 56560 93780 56566 93792
rect 192662 93780 192668 93792
rect 192720 93780 192726 93832
rect 308398 93780 308404 93832
rect 308456 93820 308462 93832
rect 420914 93820 420920 93832
rect 308456 93792 420920 93820
rect 308456 93780 308462 93792
rect 420914 93780 420920 93792
rect 420972 93780 420978 93832
rect 57790 93712 57796 93764
rect 57848 93752 57854 93764
rect 188430 93752 188436 93764
rect 57848 93724 188436 93752
rect 57848 93712 57854 93724
rect 188430 93712 188436 93724
rect 188488 93712 188494 93764
rect 291930 93712 291936 93764
rect 291988 93752 291994 93764
rect 323118 93752 323124 93764
rect 291988 93724 323124 93752
rect 291988 93712 291994 93724
rect 323118 93712 323124 93724
rect 323176 93712 323182 93764
rect 151722 93304 151728 93356
rect 151780 93344 151786 93356
rect 166258 93344 166264 93356
rect 151780 93316 166264 93344
rect 151780 93304 151786 93316
rect 166258 93304 166264 93316
rect 166316 93304 166322 93356
rect 123202 93236 123208 93288
rect 123260 93276 123266 93288
rect 170398 93276 170404 93288
rect 123260 93248 170404 93276
rect 123260 93236 123266 93248
rect 170398 93236 170404 93248
rect 170456 93236 170462 93288
rect 134702 93168 134708 93220
rect 134760 93208 134766 93220
rect 214742 93208 214748 93220
rect 134760 93180 214748 93208
rect 134760 93168 134766 93180
rect 214742 93168 214748 93180
rect 214800 93168 214806 93220
rect 320818 93168 320824 93220
rect 320876 93208 320882 93220
rect 420178 93208 420184 93220
rect 320876 93180 420184 93208
rect 320876 93168 320882 93180
rect 420178 93168 420184 93180
rect 420236 93168 420242 93220
rect 100570 93100 100576 93152
rect 100628 93140 100634 93152
rect 200942 93140 200948 93152
rect 100628 93112 200948 93140
rect 100628 93100 100634 93112
rect 200942 93100 200948 93112
rect 201000 93100 201006 93152
rect 419166 93100 419172 93152
rect 419224 93140 419230 93152
rect 580258 93140 580264 93152
rect 419224 93112 580264 93140
rect 419224 93100 419230 93112
rect 580258 93100 580264 93112
rect 580316 93100 580322 93152
rect 88058 92420 88064 92472
rect 88116 92460 88122 92472
rect 171778 92460 171784 92472
rect 88116 92432 171784 92460
rect 88116 92420 88122 92432
rect 171778 92420 171784 92432
rect 171836 92420 171842 92472
rect 202138 92420 202144 92472
rect 202196 92460 202202 92472
rect 324590 92460 324596 92472
rect 202196 92432 324596 92460
rect 202196 92420 202202 92432
rect 324590 92420 324596 92432
rect 324648 92420 324654 92472
rect 119338 92352 119344 92404
rect 119396 92392 119402 92404
rect 202322 92392 202328 92404
rect 119396 92364 202328 92392
rect 119396 92352 119402 92364
rect 202322 92352 202328 92364
rect 202380 92352 202386 92404
rect 86770 92284 86776 92336
rect 86828 92324 86834 92336
rect 129550 92324 129556 92336
rect 86828 92296 129556 92324
rect 86828 92284 86834 92296
rect 129550 92284 129556 92296
rect 129608 92284 129614 92336
rect 133138 92284 133144 92336
rect 133196 92324 133202 92336
rect 176010 92324 176016 92336
rect 133196 92296 176016 92324
rect 133196 92284 133202 92296
rect 176010 92284 176016 92296
rect 176068 92284 176074 92336
rect 129458 92216 129464 92268
rect 129516 92256 129522 92268
rect 166534 92256 166540 92268
rect 129516 92228 166540 92256
rect 129516 92216 129522 92228
rect 166534 92216 166540 92228
rect 166592 92216 166598 92268
rect 110690 92148 110696 92200
rect 110748 92188 110754 92200
rect 134702 92188 134708 92200
rect 110748 92160 134708 92188
rect 110748 92148 110754 92160
rect 134702 92148 134708 92160
rect 134760 92148 134766 92200
rect 152090 92148 152096 92200
rect 152148 92188 152154 92200
rect 189718 92188 189724 92200
rect 152148 92160 189724 92188
rect 152148 92148 152154 92160
rect 189718 92148 189724 92160
rect 189776 92148 189782 92200
rect 136082 92080 136088 92132
rect 136140 92120 136146 92132
rect 167730 92120 167736 92132
rect 136140 92092 167736 92120
rect 136140 92080 136146 92092
rect 167730 92080 167736 92092
rect 167788 92080 167794 92132
rect 199470 91740 199476 91792
rect 199528 91780 199534 91792
rect 313274 91780 313280 91792
rect 199528 91752 313280 91780
rect 199528 91740 199534 91752
rect 313274 91740 313280 91752
rect 313332 91740 313338 91792
rect 84838 91128 84844 91180
rect 84896 91168 84902 91180
rect 111150 91168 111156 91180
rect 84896 91140 111156 91168
rect 84896 91128 84902 91140
rect 111150 91128 111156 91140
rect 111208 91128 111214 91180
rect 74810 91060 74816 91112
rect 74868 91100 74874 91112
rect 111058 91100 111064 91112
rect 74868 91072 111064 91100
rect 74868 91060 74874 91072
rect 111058 91060 111064 91072
rect 111116 91060 111122 91112
rect 67634 90992 67640 91044
rect 67692 91032 67698 91044
rect 206554 91032 206560 91044
rect 67692 91004 206560 91032
rect 67692 90992 67698 91004
rect 206554 90992 206560 91004
rect 206612 90992 206618 91044
rect 210418 90992 210424 91044
rect 210476 91032 210482 91044
rect 333974 91032 333980 91044
rect 210476 91004 333980 91032
rect 210476 90992 210482 91004
rect 333974 90992 333980 91004
rect 334032 90992 334038 91044
rect 110046 90924 110052 90976
rect 110104 90964 110110 90976
rect 198274 90964 198280 90976
rect 110104 90936 198280 90964
rect 110104 90924 110110 90936
rect 198274 90924 198280 90936
rect 198332 90924 198338 90976
rect 113818 90856 113824 90908
rect 113876 90896 113882 90908
rect 178770 90896 178776 90908
rect 113876 90868 178776 90896
rect 113876 90856 113882 90868
rect 178770 90856 178776 90868
rect 178828 90856 178834 90908
rect 119890 90788 119896 90840
rect 119948 90828 119954 90840
rect 167822 90828 167828 90840
rect 119948 90800 167828 90828
rect 119948 90788 119954 90800
rect 167822 90788 167828 90800
rect 167880 90788 167886 90840
rect 151538 90720 151544 90772
rect 151596 90760 151602 90772
rect 174538 90760 174544 90772
rect 151596 90732 174544 90760
rect 151596 90720 151602 90732
rect 174538 90720 174544 90732
rect 174596 90720 174602 90772
rect 289170 90312 289176 90364
rect 289228 90352 289234 90364
rect 321554 90352 321560 90364
rect 289228 90324 321560 90352
rect 289228 90312 289234 90324
rect 321554 90312 321560 90324
rect 321612 90352 321618 90364
rect 465074 90352 465080 90364
rect 321612 90324 465080 90352
rect 321612 90312 321618 90324
rect 465074 90312 465080 90324
rect 465132 90312 465138 90364
rect 88978 89632 88984 89684
rect 89036 89672 89042 89684
rect 164878 89672 164884 89684
rect 89036 89644 164884 89672
rect 89036 89632 89042 89644
rect 164878 89632 164884 89644
rect 164936 89632 164942 89684
rect 134886 89564 134892 89616
rect 134944 89604 134950 89616
rect 209222 89604 209228 89616
rect 134944 89576 209228 89604
rect 134944 89564 134950 89576
rect 209222 89564 209228 89576
rect 209280 89564 209286 89616
rect 102042 89496 102048 89548
rect 102100 89536 102106 89548
rect 174814 89536 174820 89548
rect 102100 89508 174820 89536
rect 102100 89496 102106 89508
rect 174814 89496 174820 89508
rect 174872 89496 174878 89548
rect 111610 89428 111616 89480
rect 111668 89468 111674 89480
rect 173434 89468 173440 89480
rect 111668 89440 173440 89468
rect 111668 89428 111674 89440
rect 173434 89428 173440 89440
rect 173492 89428 173498 89480
rect 118050 89360 118056 89412
rect 118108 89400 118114 89412
rect 170490 89400 170496 89412
rect 118108 89372 170496 89400
rect 118108 89360 118114 89372
rect 170490 89360 170496 89372
rect 170548 89360 170554 89412
rect 120902 89292 120908 89344
rect 120960 89332 120966 89344
rect 170582 89332 170588 89344
rect 120960 89304 170588 89332
rect 120960 89292 120966 89304
rect 170582 89292 170588 89304
rect 170640 89292 170646 89344
rect 170398 88952 170404 89004
rect 170456 88992 170462 89004
rect 307294 88992 307300 89004
rect 170456 88964 307300 88992
rect 170456 88952 170462 88964
rect 307294 88952 307300 88964
rect 307352 88952 307358 89004
rect 316034 88952 316040 89004
rect 316092 88992 316098 89004
rect 333238 88992 333244 89004
rect 316092 88964 333244 88992
rect 316092 88952 316098 88964
rect 333238 88952 333244 88964
rect 333296 88952 333302 89004
rect 334710 88952 334716 89004
rect 334768 88992 334774 89004
rect 462314 88992 462320 89004
rect 334768 88964 462320 88992
rect 334768 88952 334774 88964
rect 462314 88952 462320 88964
rect 462372 88952 462378 89004
rect 122098 88272 122104 88324
rect 122156 88312 122162 88324
rect 210510 88312 210516 88324
rect 122156 88284 210516 88312
rect 122156 88272 122162 88284
rect 210510 88272 210516 88284
rect 210568 88272 210574 88324
rect 124122 88204 124128 88256
rect 124180 88244 124186 88256
rect 193858 88244 193864 88256
rect 124180 88216 193864 88244
rect 124180 88204 124186 88216
rect 193858 88204 193864 88216
rect 193916 88204 193922 88256
rect 97442 88136 97448 88188
rect 97500 88176 97506 88188
rect 166442 88176 166448 88188
rect 97500 88148 166448 88176
rect 97500 88136 97506 88148
rect 166442 88136 166448 88148
rect 166500 88136 166506 88188
rect 104434 88068 104440 88120
rect 104492 88108 104498 88120
rect 169294 88108 169300 88120
rect 104492 88080 169300 88108
rect 104492 88068 104498 88080
rect 169294 88068 169300 88080
rect 169352 88068 169358 88120
rect 151630 88000 151636 88052
rect 151688 88040 151694 88052
rect 213362 88040 213368 88052
rect 151688 88012 213368 88040
rect 151688 88000 151694 88012
rect 213362 88000 213368 88012
rect 213420 88000 213426 88052
rect 115290 87932 115296 87984
rect 115348 87972 115354 87984
rect 170674 87972 170680 87984
rect 115348 87944 170680 87972
rect 115348 87932 115354 87944
rect 170674 87932 170680 87944
rect 170732 87932 170738 87984
rect 318794 87660 318800 87712
rect 318852 87700 318858 87712
rect 352650 87700 352656 87712
rect 318852 87672 352656 87700
rect 318852 87660 318858 87672
rect 352650 87660 352656 87672
rect 352708 87660 352714 87712
rect 352558 87592 352564 87644
rect 352616 87632 352622 87644
rect 456794 87632 456800 87644
rect 352616 87604 456800 87632
rect 352616 87592 352622 87604
rect 456794 87592 456800 87604
rect 456852 87592 456858 87644
rect 90634 86912 90640 86964
rect 90692 86952 90698 86964
rect 202414 86952 202420 86964
rect 90692 86924 202420 86952
rect 90692 86912 90698 86924
rect 202414 86912 202420 86924
rect 202472 86912 202478 86964
rect 353294 86912 353300 86964
rect 353352 86952 353358 86964
rect 421558 86952 421564 86964
rect 353352 86924 421564 86952
rect 353352 86912 353358 86924
rect 421558 86912 421564 86924
rect 421616 86912 421622 86964
rect 504358 86912 504364 86964
rect 504416 86952 504422 86964
rect 580166 86952 580172 86964
rect 504416 86924 580172 86952
rect 504416 86912 504422 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 126054 86844 126060 86896
rect 126112 86884 126118 86896
rect 211890 86884 211896 86896
rect 126112 86856 211896 86884
rect 126112 86844 126118 86856
rect 211890 86844 211896 86856
rect 211948 86844 211954 86896
rect 107930 86776 107936 86828
rect 107988 86816 107994 86828
rect 192570 86816 192576 86828
rect 107988 86788 192576 86816
rect 107988 86776 107994 86788
rect 192570 86776 192576 86788
rect 192628 86776 192634 86828
rect 97074 86708 97080 86760
rect 97132 86748 97138 86760
rect 173158 86748 173164 86760
rect 97132 86720 173164 86748
rect 97132 86708 97138 86720
rect 173158 86708 173164 86720
rect 173216 86708 173222 86760
rect 115750 86640 115756 86692
rect 115808 86680 115814 86692
rect 178862 86680 178868 86692
rect 115808 86652 178868 86680
rect 115808 86640 115814 86652
rect 178862 86640 178868 86652
rect 178920 86640 178926 86692
rect 342254 86300 342260 86352
rect 342312 86340 342318 86352
rect 353294 86340 353300 86352
rect 342312 86312 353300 86340
rect 342312 86300 342318 86312
rect 353294 86300 353300 86312
rect 353352 86300 353358 86352
rect 178678 86232 178684 86284
rect 178736 86272 178742 86284
rect 253198 86272 253204 86284
rect 178736 86244 253204 86272
rect 178736 86232 178742 86244
rect 253198 86232 253204 86244
rect 253256 86232 253262 86284
rect 311894 86232 311900 86284
rect 311952 86272 311958 86284
rect 342346 86272 342352 86284
rect 311952 86244 342352 86272
rect 311952 86232 311958 86244
rect 342346 86232 342352 86244
rect 342404 86232 342410 86284
rect 349798 86232 349804 86284
rect 349856 86272 349862 86284
rect 455414 86272 455420 86284
rect 349856 86244 455420 86272
rect 349856 86232 349862 86244
rect 455414 86232 455420 86244
rect 455472 86232 455478 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 32398 85524 32404 85536
rect 3200 85496 32404 85524
rect 3200 85484 3206 85496
rect 32398 85484 32404 85496
rect 32456 85484 32462 85536
rect 67726 85484 67732 85536
rect 67784 85524 67790 85536
rect 214834 85524 214840 85536
rect 67784 85496 214840 85524
rect 67784 85484 67790 85496
rect 214834 85484 214840 85496
rect 214892 85484 214898 85536
rect 104618 85416 104624 85468
rect 104676 85456 104682 85468
rect 171962 85456 171968 85468
rect 104676 85428 171968 85456
rect 104676 85416 104682 85428
rect 171962 85416 171968 85428
rect 172020 85416 172026 85468
rect 100110 85348 100116 85400
rect 100168 85388 100174 85400
rect 166350 85388 166356 85400
rect 100168 85360 166356 85388
rect 100168 85348 100174 85360
rect 166350 85348 166356 85360
rect 166408 85348 166414 85400
rect 110138 85280 110144 85332
rect 110196 85320 110202 85332
rect 169110 85320 169116 85332
rect 110196 85292 169116 85320
rect 110196 85280 110202 85292
rect 169110 85280 169116 85292
rect 169168 85280 169174 85332
rect 117130 85212 117136 85264
rect 117188 85252 117194 85264
rect 174722 85252 174728 85264
rect 117188 85224 174728 85252
rect 117188 85212 117194 85224
rect 174722 85212 174728 85224
rect 174780 85212 174786 85264
rect 126698 85144 126704 85196
rect 126756 85184 126762 85196
rect 181530 85184 181536 85196
rect 126756 85156 181536 85184
rect 126756 85144 126762 85156
rect 181530 85144 181536 85156
rect 181588 85144 181594 85196
rect 336090 84804 336096 84856
rect 336148 84844 336154 84856
rect 460934 84844 460940 84856
rect 336148 84816 460940 84844
rect 336148 84804 336154 84816
rect 460934 84804 460940 84816
rect 460992 84804 460998 84856
rect 66070 84124 66076 84176
rect 66128 84164 66134 84176
rect 214558 84164 214564 84176
rect 66128 84136 214564 84164
rect 66128 84124 66134 84136
rect 214558 84124 214564 84136
rect 214616 84124 214622 84176
rect 103330 84056 103336 84108
rect 103388 84096 103394 84108
rect 196894 84096 196900 84108
rect 103388 84068 196900 84096
rect 103388 84056 103394 84068
rect 196894 84056 196900 84068
rect 196952 84056 196958 84108
rect 92382 83988 92388 84040
rect 92440 84028 92446 84040
rect 181622 84028 181628 84040
rect 92440 84000 181628 84028
rect 92440 83988 92446 84000
rect 181622 83988 181628 84000
rect 181680 83988 181686 84040
rect 125502 83920 125508 83972
rect 125560 83960 125566 83972
rect 176102 83960 176108 83972
rect 125560 83932 176108 83960
rect 125560 83920 125566 83932
rect 176102 83920 176108 83932
rect 176160 83920 176166 83972
rect 131022 83852 131028 83904
rect 131080 83892 131086 83904
rect 171870 83892 171876 83904
rect 131080 83864 171876 83892
rect 131080 83852 131086 83864
rect 171870 83852 171876 83864
rect 171928 83852 171934 83904
rect 192478 83444 192484 83496
rect 192536 83484 192542 83496
rect 315298 83484 315304 83496
rect 192536 83456 315304 83484
rect 192536 83444 192542 83456
rect 315298 83444 315304 83456
rect 315356 83444 315362 83496
rect 332042 83444 332048 83496
rect 332100 83484 332106 83496
rect 463694 83484 463700 83496
rect 332100 83456 463700 83484
rect 332100 83444 332106 83456
rect 463694 83444 463700 83456
rect 463752 83444 463758 83496
rect 103422 82764 103428 82816
rect 103480 82804 103486 82816
rect 205082 82804 205088 82816
rect 103480 82776 205088 82804
rect 103480 82764 103486 82776
rect 205082 82764 205088 82776
rect 205140 82764 205146 82816
rect 95050 82696 95056 82748
rect 95108 82736 95114 82748
rect 169202 82736 169208 82748
rect 95108 82708 169208 82736
rect 95108 82696 95114 82708
rect 169202 82696 169208 82708
rect 169260 82696 169266 82748
rect 106182 82628 106188 82680
rect 106240 82668 106246 82680
rect 177574 82668 177580 82680
rect 106240 82640 177580 82668
rect 106240 82628 106246 82640
rect 177574 82628 177580 82640
rect 177632 82628 177638 82680
rect 122742 82560 122748 82612
rect 122800 82600 122806 82612
rect 184290 82600 184296 82612
rect 122800 82572 184296 82600
rect 122800 82560 122806 82572
rect 184290 82560 184296 82572
rect 184348 82560 184354 82612
rect 126882 82492 126888 82544
rect 126940 82532 126946 82544
rect 167638 82532 167644 82544
rect 126940 82504 167644 82532
rect 126940 82492 126946 82504
rect 167638 82492 167644 82504
rect 167696 82492 167702 82544
rect 216030 82220 216036 82272
rect 216088 82260 216094 82272
rect 239398 82260 239404 82272
rect 216088 82232 239404 82260
rect 216088 82220 216094 82232
rect 239398 82220 239404 82232
rect 239456 82220 239462 82272
rect 207658 82152 207664 82204
rect 207716 82192 207722 82204
rect 232498 82192 232504 82204
rect 207716 82164 232504 82192
rect 207716 82152 207722 82164
rect 232498 82152 232504 82164
rect 232556 82152 232562 82204
rect 195330 82084 195336 82136
rect 195388 82124 195394 82136
rect 246298 82124 246304 82136
rect 195388 82096 246304 82124
rect 195388 82084 195394 82096
rect 246298 82084 246304 82096
rect 246356 82084 246362 82136
rect 324314 82084 324320 82136
rect 324372 82124 324378 82136
rect 461578 82124 461584 82136
rect 324372 82096 461584 82124
rect 324372 82084 324378 82096
rect 461578 82084 461584 82096
rect 461636 82084 461642 82136
rect 107470 81336 107476 81388
rect 107528 81376 107534 81388
rect 196802 81376 196808 81388
rect 107528 81348 196808 81376
rect 107528 81336 107534 81348
rect 196802 81336 196808 81348
rect 196860 81336 196866 81388
rect 351914 81336 351920 81388
rect 351972 81376 351978 81388
rect 465718 81376 465724 81388
rect 351972 81348 465724 81376
rect 351972 81336 351978 81348
rect 465718 81336 465724 81348
rect 465776 81336 465782 81388
rect 121362 81268 121368 81320
rect 121420 81308 121426 81320
rect 206462 81308 206468 81320
rect 121420 81280 206468 81308
rect 121420 81268 121426 81280
rect 206462 81268 206468 81280
rect 206520 81268 206526 81320
rect 95142 81200 95148 81252
rect 95200 81240 95206 81252
rect 167914 81240 167920 81252
rect 95200 81212 167920 81240
rect 95200 81200 95206 81212
rect 167914 81200 167920 81212
rect 167972 81200 167978 81252
rect 118602 81132 118608 81184
rect 118660 81172 118666 81184
rect 182910 81172 182916 81184
rect 118660 81144 182916 81172
rect 118660 81132 118666 81144
rect 182910 81132 182916 81144
rect 182968 81132 182974 81184
rect 187050 80656 187056 80708
rect 187108 80696 187114 80708
rect 307110 80696 307116 80708
rect 187108 80668 307116 80696
rect 187108 80656 187114 80668
rect 307110 80656 307116 80668
rect 307168 80656 307174 80708
rect 317414 80656 317420 80708
rect 317472 80696 317478 80708
rect 351914 80696 351920 80708
rect 317472 80668 351920 80696
rect 317472 80656 317478 80668
rect 351914 80656 351920 80668
rect 351972 80656 351978 80708
rect 114370 79976 114376 80028
rect 114428 80016 114434 80028
rect 213454 80016 213460 80028
rect 114428 79988 213460 80016
rect 114428 79976 114434 79988
rect 213454 79976 213460 79988
rect 213512 79976 213518 80028
rect 96522 79908 96528 79960
rect 96580 79948 96586 79960
rect 178954 79948 178960 79960
rect 96580 79920 178960 79948
rect 96580 79908 96586 79920
rect 178954 79908 178960 79920
rect 179012 79908 179018 79960
rect 93762 79840 93768 79892
rect 93820 79880 93826 79892
rect 169018 79880 169024 79892
rect 93820 79852 169024 79880
rect 93820 79840 93826 79852
rect 169018 79840 169024 79852
rect 169076 79840 169082 79892
rect 101950 79772 101956 79824
rect 102008 79812 102014 79824
rect 173250 79812 173256 79824
rect 102008 79784 173256 79812
rect 102008 79772 102014 79784
rect 173250 79772 173256 79784
rect 173308 79772 173314 79824
rect 209038 79432 209044 79484
rect 209096 79472 209102 79484
rect 238018 79472 238024 79484
rect 209096 79444 238024 79472
rect 209096 79432 209102 79444
rect 238018 79432 238024 79444
rect 238076 79432 238082 79484
rect 198090 79364 198096 79416
rect 198148 79404 198154 79416
rect 244918 79404 244924 79416
rect 198148 79376 244924 79404
rect 198148 79364 198154 79376
rect 244918 79364 244924 79376
rect 244976 79364 244982 79416
rect 173158 79296 173164 79348
rect 173216 79336 173222 79348
rect 307202 79336 307208 79348
rect 173216 79308 307208 79336
rect 173216 79296 173222 79308
rect 307202 79296 307208 79308
rect 307260 79296 307266 79348
rect 309778 79296 309784 79348
rect 309836 79336 309842 79348
rect 470594 79336 470600 79348
rect 309836 79308 470600 79336
rect 309836 79296 309842 79308
rect 470594 79296 470600 79308
rect 470652 79296 470658 79348
rect 110322 78616 110328 78668
rect 110380 78656 110386 78668
rect 177482 78656 177488 78668
rect 110380 78628 177488 78656
rect 110380 78616 110386 78628
rect 177482 78616 177488 78628
rect 177540 78616 177546 78668
rect 339402 78616 339408 78668
rect 339460 78656 339466 78668
rect 471974 78656 471980 78668
rect 339460 78628 471980 78656
rect 339460 78616 339466 78628
rect 471974 78616 471980 78628
rect 472032 78616 472038 78668
rect 128262 78548 128268 78600
rect 128320 78588 128326 78600
rect 187142 78588 187148 78600
rect 128320 78560 187148 78588
rect 128320 78548 128326 78560
rect 187142 78548 187148 78560
rect 187200 78548 187206 78600
rect 269942 78072 269948 78124
rect 270000 78112 270006 78124
rect 334618 78112 334624 78124
rect 270000 78084 334624 78112
rect 270000 78072 270006 78084
rect 334618 78072 334624 78084
rect 334676 78072 334682 78124
rect 196618 78004 196624 78056
rect 196676 78044 196682 78056
rect 279510 78044 279516 78056
rect 196676 78016 279516 78044
rect 196676 78004 196682 78016
rect 279510 78004 279516 78016
rect 279568 78004 279574 78056
rect 45554 77936 45560 77988
rect 45612 77976 45618 77988
rect 297542 77976 297548 77988
rect 45612 77948 297548 77976
rect 45612 77936 45618 77948
rect 297542 77936 297548 77948
rect 297600 77936 297606 77988
rect 303614 77256 303620 77308
rect 303672 77296 303678 77308
rect 339402 77296 339408 77308
rect 303672 77268 339408 77296
rect 303672 77256 303678 77268
rect 339402 77256 339408 77268
rect 339460 77256 339466 77308
rect 111150 77188 111156 77240
rect 111208 77228 111214 77240
rect 200850 77228 200856 77240
rect 111208 77200 200856 77228
rect 111208 77188 111214 77200
rect 200850 77188 200856 77200
rect 200908 77188 200914 77240
rect 99282 77120 99288 77172
rect 99340 77160 99346 77172
rect 173342 77160 173348 77172
rect 99340 77132 173348 77160
rect 99340 77120 99346 77132
rect 173342 77120 173348 77132
rect 173400 77120 173406 77172
rect 199378 76644 199384 76696
rect 199436 76684 199442 76696
rect 199436 76656 287054 76684
rect 199436 76644 199442 76656
rect 287026 76628 287054 76656
rect 86954 76576 86960 76628
rect 87012 76616 87018 76628
rect 285122 76616 285128 76628
rect 87012 76588 285128 76616
rect 87012 76576 87018 76588
rect 285122 76576 285128 76588
rect 285180 76576 285186 76628
rect 287026 76588 287060 76628
rect 287054 76576 287060 76588
rect 287112 76616 287118 76628
rect 335998 76616 336004 76628
rect 287112 76588 336004 76616
rect 287112 76576 287118 76588
rect 335998 76576 336004 76588
rect 336056 76576 336062 76628
rect 2774 76508 2780 76560
rect 2832 76548 2838 76560
rect 294782 76548 294788 76560
rect 2832 76520 294788 76548
rect 2832 76508 2838 76520
rect 294782 76508 294788 76520
rect 294840 76508 294846 76560
rect 14 75828 20 75880
rect 72 75868 78 75880
rect 1302 75868 1308 75880
rect 72 75840 1308 75868
rect 72 75828 78 75840
rect 1302 75828 1308 75840
rect 1360 75868 1366 75880
rect 249150 75868 249156 75880
rect 1360 75840 249156 75868
rect 1360 75828 1366 75840
rect 249150 75828 249156 75840
rect 249208 75828 249214 75880
rect 111058 75760 111064 75812
rect 111116 75800 111122 75812
rect 203610 75800 203616 75812
rect 111116 75772 203616 75800
rect 111116 75760 111122 75772
rect 203610 75760 203616 75772
rect 203668 75760 203674 75812
rect 69014 75216 69020 75268
rect 69072 75256 69078 75268
rect 300394 75256 300400 75268
rect 69072 75228 300400 75256
rect 69072 75216 69078 75228
rect 300394 75216 300400 75228
rect 300452 75216 300458 75268
rect 63402 75148 63408 75200
rect 63460 75188 63466 75200
rect 309870 75188 309876 75200
rect 63460 75160 309876 75188
rect 63460 75148 63466 75160
rect 309870 75148 309876 75160
rect 309928 75148 309934 75200
rect 312538 75148 312544 75200
rect 312596 75188 312602 75200
rect 469214 75188 469220 75200
rect 312596 75160 469220 75188
rect 312596 75148 312602 75160
rect 469214 75148 469220 75160
rect 469272 75148 469278 75200
rect 343726 74468 343732 74520
rect 343784 74508 343790 74520
rect 459554 74508 459560 74520
rect 343784 74480 459560 74508
rect 343784 74468 343790 74480
rect 459554 74468 459560 74480
rect 459612 74468 459618 74520
rect 110414 73924 110420 73976
rect 110472 73964 110478 73976
rect 257430 73964 257436 73976
rect 110472 73936 257436 73964
rect 110472 73924 110478 73936
rect 257430 73924 257436 73936
rect 257488 73924 257494 73976
rect 80054 73856 80060 73908
rect 80112 73896 80118 73908
rect 304442 73896 304448 73908
rect 80112 73868 304448 73896
rect 80112 73856 80118 73868
rect 304442 73856 304448 73868
rect 304500 73856 304506 73908
rect 61930 73788 61936 73840
rect 61988 73828 61994 73840
rect 338850 73828 338856 73840
rect 61988 73800 338856 73828
rect 61988 73788 61994 73800
rect 338850 73788 338856 73800
rect 338908 73788 338914 73840
rect 339494 73176 339500 73228
rect 339552 73216 339558 73228
rect 343726 73216 343732 73228
rect 339552 73188 343732 73216
rect 339552 73176 339558 73188
rect 343726 73176 343732 73188
rect 343784 73176 343790 73228
rect 419350 73108 419356 73160
rect 419408 73148 419414 73160
rect 579982 73148 579988 73160
rect 419408 73120 579988 73148
rect 419408 73108 419414 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 352098 73040 352104 73092
rect 352156 73080 352162 73092
rect 426526 73080 426532 73092
rect 352156 73052 426532 73080
rect 352156 73040 352162 73052
rect 426526 73040 426532 73052
rect 426584 73040 426590 73092
rect 114554 72564 114560 72616
rect 114612 72604 114618 72616
rect 289354 72604 289360 72616
rect 114612 72576 289360 72604
rect 114612 72564 114618 72576
rect 289354 72564 289360 72576
rect 289412 72564 289418 72616
rect 44082 72496 44088 72548
rect 44140 72536 44146 72548
rect 240778 72536 240784 72548
rect 44140 72508 240784 72536
rect 44140 72496 44146 72508
rect 240778 72496 240784 72508
rect 240836 72496 240842 72548
rect 59354 72428 59360 72480
rect 59412 72468 59418 72480
rect 301682 72468 301688 72480
rect 59412 72440 301688 72468
rect 59412 72428 59418 72440
rect 301682 72428 301688 72440
rect 301740 72428 301746 72480
rect 345750 71748 345756 71800
rect 345808 71788 345814 71800
rect 352098 71788 352104 71800
rect 345808 71760 352104 71788
rect 345808 71748 345814 71760
rect 352098 71748 352104 71760
rect 352156 71748 352162 71800
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 52362 71720 52368 71732
rect 3476 71692 52368 71720
rect 3476 71680 3482 71692
rect 52362 71680 52368 71692
rect 52420 71720 52426 71732
rect 495710 71720 495716 71732
rect 52420 71692 495716 71720
rect 52420 71680 52426 71692
rect 495710 71680 495716 71692
rect 495768 71680 495774 71732
rect 41322 71612 41328 71664
rect 41380 71652 41386 71664
rect 332042 71652 332048 71664
rect 41380 71624 332048 71652
rect 41380 71612 41386 71624
rect 332042 71612 332048 71624
rect 332100 71612 332106 71664
rect 186958 71068 186964 71120
rect 187016 71108 187022 71120
rect 333238 71108 333244 71120
rect 187016 71080 333244 71108
rect 187016 71068 187022 71080
rect 333238 71068 333244 71080
rect 333296 71068 333302 71120
rect 84194 71000 84200 71052
rect 84252 71040 84258 71052
rect 253290 71040 253296 71052
rect 84252 71012 253296 71040
rect 84252 71000 84258 71012
rect 253290 71000 253296 71012
rect 253348 71000 253354 71052
rect 331306 70524 331312 70576
rect 331364 70564 331370 70576
rect 332042 70564 332048 70576
rect 331364 70536 332048 70564
rect 331364 70524 331370 70536
rect 332042 70524 332048 70536
rect 332100 70524 332106 70576
rect 333238 70388 333244 70440
rect 333296 70428 333302 70440
rect 334710 70428 334716 70440
rect 333296 70400 334716 70428
rect 333296 70388 333302 70400
rect 334710 70388 334716 70400
rect 334768 70388 334774 70440
rect 204990 69776 204996 69828
rect 205048 69816 205054 69828
rect 289814 69816 289820 69828
rect 205048 69788 289820 69816
rect 205048 69776 205054 69788
rect 289814 69776 289820 69788
rect 289872 69776 289878 69828
rect 63310 69708 63316 69760
rect 63368 69748 63374 69760
rect 292574 69748 292580 69760
rect 63368 69720 292580 69748
rect 63368 69708 63374 69720
rect 292574 69708 292580 69720
rect 292632 69708 292638 69760
rect 40034 69640 40040 69692
rect 40092 69680 40098 69692
rect 280982 69680 280988 69692
rect 40092 69652 280988 69680
rect 40092 69640 40098 69652
rect 280982 69640 280988 69652
rect 281040 69640 281046 69692
rect 297542 69640 297548 69692
rect 297600 69680 297606 69692
rect 472618 69680 472624 69692
rect 297600 69652 472624 69680
rect 297600 69640 297606 69652
rect 472618 69640 472624 69652
rect 472676 69640 472682 69692
rect 60550 68960 60556 69012
rect 60608 69000 60614 69012
rect 335354 69000 335360 69012
rect 60608 68972 335360 69000
rect 60608 68960 60614 68972
rect 335354 68960 335360 68972
rect 335412 69000 335418 69012
rect 336090 69000 336096 69012
rect 335412 68972 336096 69000
rect 335412 68960 335418 68972
rect 336090 68960 336096 68972
rect 336148 68960 336154 69012
rect 292574 68892 292580 68944
rect 292632 68932 292638 68944
rect 474734 68932 474740 68944
rect 292632 68904 474740 68932
rect 292632 68892 292638 68904
rect 474734 68892 474740 68904
rect 474792 68892 474798 68944
rect 93854 68348 93860 68400
rect 93912 68388 93918 68400
rect 293310 68388 293316 68400
rect 93912 68360 293316 68388
rect 93912 68348 93918 68360
rect 293310 68348 293316 68360
rect 293368 68348 293374 68400
rect 20714 68280 20720 68332
rect 20772 68320 20778 68332
rect 254762 68320 254768 68332
rect 20772 68292 254768 68320
rect 20772 68280 20778 68292
rect 254762 68280 254768 68292
rect 254820 68280 254826 68332
rect 2682 67532 2688 67584
rect 2740 67572 2746 67584
rect 5442 67572 5448 67584
rect 2740 67544 5448 67572
rect 2740 67532 2746 67544
rect 5442 67532 5448 67544
rect 5500 67572 5506 67584
rect 251358 67572 251364 67584
rect 5500 67544 251364 67572
rect 5500 67532 5506 67544
rect 251358 67532 251364 67544
rect 251416 67532 251422 67584
rect 289814 67532 289820 67584
rect 289872 67572 289878 67584
rect 476114 67572 476120 67584
rect 289872 67544 476120 67572
rect 289872 67532 289878 67544
rect 476114 67532 476120 67544
rect 476172 67532 476178 67584
rect 180150 66920 180156 66972
rect 180208 66960 180214 66972
rect 257338 66960 257344 66972
rect 180208 66932 257344 66960
rect 180208 66920 180214 66932
rect 257338 66920 257344 66932
rect 257396 66920 257402 66972
rect 262214 66920 262220 66972
rect 262272 66960 262278 66972
rect 338758 66960 338764 66972
rect 262272 66932 338764 66960
rect 262272 66920 262278 66932
rect 338758 66920 338764 66932
rect 338816 66920 338822 66972
rect 62114 66852 62120 66904
rect 62172 66892 62178 66904
rect 292114 66892 292120 66904
rect 62172 66864 292120 66892
rect 62172 66852 62178 66864
rect 292114 66852 292120 66864
rect 292172 66852 292178 66904
rect 61838 66172 61844 66224
rect 61896 66212 61902 66224
rect 269114 66212 269120 66224
rect 61896 66184 269120 66212
rect 61896 66172 61902 66184
rect 269114 66172 269120 66184
rect 269172 66212 269178 66224
rect 269942 66212 269948 66224
rect 269172 66184 269948 66212
rect 269172 66172 269178 66184
rect 269942 66172 269948 66184
rect 270000 66172 270006 66224
rect 285674 66172 285680 66224
rect 285732 66212 285738 66224
rect 286318 66212 286324 66224
rect 285732 66184 286324 66212
rect 285732 66172 285738 66184
rect 286318 66172 286324 66184
rect 286376 66212 286382 66224
rect 477494 66212 477500 66224
rect 286376 66184 477500 66212
rect 286376 66172 286382 66184
rect 477494 66172 477500 66184
rect 477552 66172 477558 66224
rect 121454 65560 121460 65612
rect 121512 65600 121518 65612
rect 305914 65600 305920 65612
rect 121512 65572 305920 65600
rect 121512 65560 121518 65572
rect 305914 65560 305920 65572
rect 305972 65560 305978 65612
rect 31754 65492 31760 65544
rect 31812 65532 31818 65544
rect 273990 65532 273996 65544
rect 31812 65504 273996 65532
rect 31812 65492 31818 65504
rect 273990 65492 273996 65504
rect 274048 65492 274054 65544
rect 60642 64812 60648 64864
rect 60700 64852 60706 64864
rect 273254 64852 273260 64864
rect 60700 64824 273260 64852
rect 60700 64812 60706 64824
rect 273254 64812 273260 64824
rect 273312 64812 273318 64864
rect 279510 64812 279516 64864
rect 279568 64852 279574 64864
rect 480254 64852 480260 64864
rect 279568 64824 480260 64852
rect 279568 64812 279574 64824
rect 480254 64812 480260 64824
rect 480312 64812 480318 64864
rect 273254 64404 273260 64456
rect 273312 64444 273318 64456
rect 274082 64444 274088 64456
rect 273312 64416 274088 64444
rect 273312 64404 273318 64416
rect 274082 64404 274088 64416
rect 274140 64404 274146 64456
rect 73154 64132 73160 64184
rect 73212 64172 73218 64184
rect 293218 64172 293224 64184
rect 73212 64144 293224 64172
rect 73212 64132 73218 64144
rect 293218 64132 293224 64144
rect 293276 64132 293282 64184
rect 278774 63520 278780 63572
rect 278832 63560 278838 63572
rect 279510 63560 279516 63572
rect 278832 63532 279516 63560
rect 278832 63520 278838 63532
rect 279510 63520 279516 63532
rect 279568 63520 279574 63572
rect 97994 62840 98000 62892
rect 98052 62880 98058 62892
rect 298830 62880 298836 62892
rect 98052 62852 298836 62880
rect 98052 62840 98058 62852
rect 298830 62840 298836 62852
rect 298888 62840 298894 62892
rect 278222 62772 278228 62824
rect 278280 62812 278286 62824
rect 481726 62812 481732 62824
rect 278280 62784 481732 62812
rect 278280 62772 278286 62784
rect 481726 62772 481732 62784
rect 481784 62772 481790 62824
rect 274634 62024 274640 62076
rect 274692 62064 274698 62076
rect 481634 62064 481640 62076
rect 274692 62036 481640 62064
rect 274692 62024 274698 62036
rect 481634 62024 481640 62036
rect 481692 62024 481698 62076
rect 104894 61480 104900 61532
rect 104952 61520 104958 61532
rect 272610 61520 272616 61532
rect 104952 61492 272616 61520
rect 104952 61480 104958 61492
rect 272610 61480 272616 61492
rect 272668 61480 272674 61532
rect 59170 61412 59176 61464
rect 59228 61452 59234 61464
rect 285122 61452 285128 61464
rect 59228 61424 285128 61452
rect 59228 61412 59234 61424
rect 285122 61412 285128 61424
rect 285180 61412 285186 61464
rect 17954 61344 17960 61396
rect 18012 61384 18018 61396
rect 300302 61384 300308 61396
rect 18012 61356 300308 61384
rect 18012 61344 18018 61356
rect 300302 61344 300308 61356
rect 300360 61344 300366 61396
rect 271874 60732 271880 60784
rect 271932 60772 271938 60784
rect 274634 60772 274640 60784
rect 271932 60744 274640 60772
rect 271932 60732 271938 60744
rect 274634 60732 274640 60744
rect 274692 60732 274698 60784
rect 513282 60664 513288 60716
rect 513340 60704 513346 60716
rect 580166 60704 580172 60716
rect 513340 60676 580172 60704
rect 513340 60664 513346 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 118694 60052 118700 60104
rect 118752 60092 118758 60104
rect 279418 60092 279424 60104
rect 118752 60064 279424 60092
rect 118752 60052 118758 60064
rect 279418 60052 279424 60064
rect 279476 60052 279482 60104
rect 15194 59984 15200 60036
rect 15252 60024 15258 60036
rect 258810 60024 258816 60036
rect 15252 59996 258816 60024
rect 15252 59984 15258 59996
rect 258810 59984 258816 59996
rect 258868 59984 258874 60036
rect 268562 59984 268568 60036
rect 268620 60024 268626 60036
rect 483014 60024 483020 60036
rect 268620 59996 483020 60024
rect 268620 59984 268626 59996
rect 483014 59984 483020 59996
rect 483072 59984 483078 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 25498 59344 25504 59356
rect 3108 59316 25504 59344
rect 3108 59304 3114 59316
rect 25498 59304 25504 59316
rect 25556 59304 25562 59356
rect 211798 58828 211804 58880
rect 211856 58868 211862 58880
rect 264974 58868 264980 58880
rect 211856 58840 264980 58868
rect 211856 58828 211862 58840
rect 264974 58828 264980 58840
rect 265032 58868 265038 58880
rect 265032 58840 267734 58868
rect 265032 58828 265038 58840
rect 74534 58760 74540 58812
rect 74592 58800 74598 58812
rect 254670 58800 254676 58812
rect 74592 58772 254676 58800
rect 74592 58760 74598 58772
rect 254670 58760 254676 58772
rect 254728 58760 254734 58812
rect 267706 58800 267734 58840
rect 484394 58800 484400 58812
rect 267706 58772 484400 58800
rect 484394 58760 484400 58772
rect 484452 58760 484458 58812
rect 56594 58692 56600 58744
rect 56652 58732 56658 58744
rect 278038 58732 278044 58744
rect 56652 58704 278044 58732
rect 56652 58692 56658 58704
rect 278038 58692 278044 58704
rect 278096 58692 278102 58744
rect 57882 58624 57888 58676
rect 57940 58664 57946 58676
rect 332594 58664 332600 58676
rect 57940 58636 332600 58664
rect 57940 58624 57946 58636
rect 332594 58624 332600 58636
rect 332652 58624 332658 58676
rect 261662 57876 261668 57928
rect 261720 57916 261726 57928
rect 485774 57916 485780 57928
rect 261720 57888 485780 57916
rect 261720 57876 261726 57888
rect 485774 57876 485780 57888
rect 485832 57876 485838 57928
rect 414658 57848 414664 57860
rect 335326 57820 414664 57848
rect 332594 57740 332600 57792
rect 332652 57780 332658 57792
rect 335326 57780 335354 57820
rect 414658 57808 414664 57820
rect 414716 57808 414722 57860
rect 332652 57752 335354 57780
rect 332652 57740 332658 57752
rect 260834 57672 260840 57724
rect 260892 57712 260898 57724
rect 261662 57712 261668 57724
rect 260892 57684 261668 57712
rect 260892 57672 260898 57684
rect 261662 57672 261668 57684
rect 261720 57672 261726 57724
rect 102134 57332 102140 57384
rect 102192 57372 102198 57384
rect 305822 57372 305828 57384
rect 102192 57344 305828 57372
rect 102192 57332 102198 57344
rect 305822 57332 305828 57344
rect 305880 57332 305886 57384
rect 52454 57264 52460 57316
rect 52512 57304 52518 57316
rect 261570 57304 261576 57316
rect 52512 57276 261576 57304
rect 52512 57264 52518 57276
rect 261570 57264 261576 57276
rect 261628 57264 261634 57316
rect 6914 57196 6920 57248
rect 6972 57236 6978 57248
rect 264514 57236 264520 57248
rect 6972 57208 264520 57236
rect 6972 57196 6978 57208
rect 264514 57196 264520 57208
rect 264572 57196 264578 57248
rect 209130 56040 209136 56092
rect 209188 56080 209194 56092
rect 253934 56080 253940 56092
rect 209188 56052 253940 56080
rect 209188 56040 209194 56052
rect 253934 56040 253940 56052
rect 253992 56040 253998 56092
rect 51074 55972 51080 56024
rect 51132 56012 51138 56024
rect 264422 56012 264428 56024
rect 51132 55984 264428 56012
rect 51132 55972 51138 55984
rect 264422 55972 264428 55984
rect 264480 55972 264486 56024
rect 67634 55904 67640 55956
rect 67692 55944 67698 55956
rect 297450 55944 297456 55956
rect 67692 55916 297456 55944
rect 67692 55904 67698 55916
rect 297450 55904 297456 55916
rect 297508 55904 297514 55956
rect 117314 55836 117320 55888
rect 117372 55876 117378 55888
rect 250622 55876 250628 55888
rect 117372 55848 250628 55876
rect 117372 55836 117378 55848
rect 250622 55836 250628 55848
rect 250680 55836 250686 55888
rect 253934 55836 253940 55888
rect 253992 55876 253998 55888
rect 488534 55876 488540 55888
rect 253992 55848 488540 55876
rect 253992 55836 253998 55848
rect 488534 55836 488540 55848
rect 488592 55836 488598 55888
rect 78674 54680 78680 54732
rect 78732 54720 78738 54732
rect 290550 54720 290556 54732
rect 78732 54692 290556 54720
rect 78732 54680 78738 54692
rect 290550 54680 290556 54692
rect 290608 54680 290614 54732
rect 70394 54612 70400 54664
rect 70452 54652 70458 54664
rect 304350 54652 304356 54664
rect 70452 54624 304356 54652
rect 70452 54612 70458 54624
rect 304350 54612 304356 54624
rect 304408 54612 304414 54664
rect 253014 54544 253020 54596
rect 253072 54584 253078 54596
rect 489914 54584 489920 54596
rect 253072 54556 489920 54584
rect 253072 54544 253078 54556
rect 489914 54544 489920 54556
rect 489972 54544 489978 54596
rect 11054 54476 11060 54528
rect 11112 54516 11118 54528
rect 253382 54516 253388 54528
rect 11112 54488 253388 54516
rect 11112 54476 11118 54488
rect 253382 54476 253388 54488
rect 253440 54476 253446 54528
rect 60734 53184 60740 53236
rect 60792 53224 60798 53236
rect 264330 53224 264336 53236
rect 60792 53196 264336 53224
rect 60792 53184 60798 53196
rect 264330 53184 264336 53196
rect 264388 53184 264394 53236
rect 4154 53116 4160 53168
rect 4212 53156 4218 53168
rect 247678 53156 247684 53168
rect 4212 53128 247684 53156
rect 4212 53116 4218 53128
rect 247678 53116 247684 53128
rect 247736 53116 247742 53168
rect 247770 53116 247776 53168
rect 247828 53156 247834 53168
rect 491294 53156 491300 53168
rect 247828 53128 491300 53156
rect 247828 53116 247834 53128
rect 491294 53116 491300 53128
rect 491352 53116 491358 53168
rect 37274 53048 37280 53100
rect 37332 53088 37338 53100
rect 296254 53088 296260 53100
rect 37332 53060 296260 53088
rect 37332 53048 37338 53060
rect 296254 53048 296260 53060
rect 296312 53048 296318 53100
rect 243538 52368 243544 52420
rect 243596 52408 243602 52420
rect 467098 52408 467104 52420
rect 243596 52380 467104 52408
rect 243596 52368 243602 52380
rect 467098 52368 467104 52380
rect 467156 52368 467162 52420
rect 35802 52300 35808 52352
rect 35860 52340 35866 52352
rect 252646 52340 252652 52352
rect 35860 52312 252652 52340
rect 35860 52300 35866 52312
rect 252646 52300 252652 52312
rect 252704 52340 252710 52352
rect 253014 52340 253020 52352
rect 252704 52312 253020 52340
rect 252704 52300 252710 52312
rect 253014 52300 253020 52312
rect 253072 52300 253078 52352
rect 202230 52232 202236 52284
rect 202288 52272 202294 52284
rect 247034 52272 247040 52284
rect 202288 52244 247040 52272
rect 202288 52232 202294 52244
rect 247034 52232 247040 52244
rect 247092 52272 247098 52284
rect 247770 52272 247776 52284
rect 247092 52244 247776 52272
rect 247092 52232 247098 52244
rect 247770 52232 247776 52244
rect 247828 52232 247834 52284
rect 69106 51688 69112 51740
rect 69164 51728 69170 51740
rect 300210 51728 300216 51740
rect 69164 51700 300216 51728
rect 69164 51688 69170 51700
rect 300210 51688 300216 51700
rect 300268 51688 300274 51740
rect 242894 51076 242900 51128
rect 242952 51116 242958 51128
rect 243538 51116 243544 51128
rect 242952 51088 243544 51116
rect 242952 51076 242958 51088
rect 243538 51076 243544 51088
rect 243596 51076 243602 51128
rect 240778 51008 240784 51060
rect 240836 51048 240842 51060
rect 492674 51048 492680 51060
rect 240836 51020 492680 51048
rect 240836 51008 240842 51020
rect 492674 51008 492680 51020
rect 492732 51008 492738 51060
rect 240134 50532 240140 50584
rect 240192 50572 240198 50584
rect 240778 50572 240784 50584
rect 240192 50544 240784 50572
rect 240192 50532 240198 50544
rect 240778 50532 240784 50544
rect 240836 50532 240842 50584
rect 71774 50464 71780 50516
rect 71832 50504 71838 50516
rect 249058 50504 249064 50516
rect 71832 50476 249064 50504
rect 71832 50464 71838 50476
rect 249058 50464 249064 50476
rect 249116 50464 249122 50516
rect 85574 50396 85580 50448
rect 85632 50436 85638 50448
rect 300118 50436 300124 50448
rect 85632 50408 300124 50436
rect 85632 50396 85638 50408
rect 300118 50396 300124 50408
rect 300176 50396 300182 50448
rect 41414 50328 41420 50380
rect 41472 50368 41478 50380
rect 269850 50368 269856 50380
rect 41472 50340 269856 50368
rect 41472 50328 41478 50340
rect 269850 50328 269856 50340
rect 269908 50328 269914 50380
rect 311158 49648 311164 49700
rect 311216 49688 311222 49700
rect 312538 49688 312544 49700
rect 311216 49660 312544 49688
rect 311216 49648 311222 49660
rect 312538 49648 312544 49660
rect 312596 49648 312602 49700
rect 124214 49104 124220 49156
rect 124272 49144 124278 49156
rect 260098 49144 260104 49156
rect 124272 49116 260104 49144
rect 124272 49104 124278 49116
rect 260098 49104 260104 49116
rect 260156 49104 260162 49156
rect 267182 49104 267188 49156
rect 267240 49144 267246 49156
rect 353938 49144 353944 49156
rect 267240 49116 353944 49144
rect 267240 49104 267246 49116
rect 353938 49104 353944 49116
rect 353996 49104 354002 49156
rect 64598 49036 64604 49088
rect 64656 49076 64662 49088
rect 311158 49076 311164 49088
rect 64656 49048 311164 49076
rect 64656 49036 64662 49048
rect 311158 49036 311164 49048
rect 311216 49036 311222 49088
rect 9674 48968 9680 49020
rect 9732 49008 9738 49020
rect 292022 49008 292028 49020
rect 9732 48980 292028 49008
rect 9732 48968 9738 48980
rect 292022 48968 292028 48980
rect 292080 48968 292086 49020
rect 349154 48968 349160 49020
rect 349212 49008 349218 49020
rect 495618 49008 495624 49020
rect 349212 48980 495624 49008
rect 349212 48968 349218 48980
rect 495618 48968 495624 48980
rect 495676 48968 495682 49020
rect 367830 48220 367836 48272
rect 367888 48260 367894 48272
rect 495526 48260 495532 48272
rect 367888 48232 495532 48260
rect 367888 48220 367894 48232
rect 495526 48220 495532 48232
rect 495584 48220 495590 48272
rect 122834 47676 122840 47728
rect 122892 47716 122898 47728
rect 268470 47716 268476 47728
rect 122892 47688 268476 47716
rect 122892 47676 122898 47688
rect 268470 47676 268476 47688
rect 268528 47676 268534 47728
rect 273898 47676 273904 47728
rect 273956 47716 273962 47728
rect 276014 47716 276020 47728
rect 273956 47688 276020 47716
rect 273956 47676 273962 47688
rect 276014 47676 276020 47688
rect 276072 47716 276078 47728
rect 345658 47716 345664 47728
rect 276072 47688 345664 47716
rect 276072 47676 276078 47688
rect 345658 47676 345664 47688
rect 345716 47676 345722 47728
rect 34514 47608 34520 47660
rect 34572 47648 34578 47660
rect 278130 47648 278136 47660
rect 34572 47620 278136 47648
rect 34572 47608 34578 47620
rect 278130 47608 278136 47620
rect 278188 47608 278194 47660
rect 64690 47540 64696 47592
rect 64748 47580 64754 47592
rect 327718 47580 327724 47592
rect 64748 47552 327724 47580
rect 64748 47540 64754 47552
rect 327718 47540 327724 47552
rect 327776 47540 327782 47592
rect 345014 47540 345020 47592
rect 345072 47580 345078 47592
rect 367094 47580 367100 47592
rect 345072 47552 367100 47580
rect 345072 47540 345078 47552
rect 367094 47540 367100 47552
rect 367152 47580 367158 47592
rect 367830 47580 367836 47592
rect 367152 47552 367836 47580
rect 367152 47540 367158 47552
rect 367830 47540 367836 47552
rect 367888 47540 367894 47592
rect 206370 46860 206376 46912
rect 206428 46900 206434 46912
rect 349154 46900 349160 46912
rect 206428 46872 349160 46900
rect 206428 46860 206434 46872
rect 349154 46860 349160 46872
rect 349212 46860 349218 46912
rect 555418 46860 555424 46912
rect 555476 46900 555482 46912
rect 580166 46900 580172 46912
rect 555476 46872 580172 46900
rect 555476 46860 555482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 45462 46248 45468 46300
rect 45520 46288 45526 46300
rect 291194 46288 291200 46300
rect 45520 46260 291200 46288
rect 45520 46248 45526 46260
rect 291194 46248 291200 46260
rect 291252 46288 291258 46300
rect 356790 46288 356796 46300
rect 291252 46260 356796 46288
rect 291252 46248 291258 46260
rect 356790 46248 356796 46260
rect 356848 46248 356854 46300
rect 2866 46180 2872 46232
rect 2924 46220 2930 46232
rect 289262 46220 289268 46232
rect 2924 46192 289268 46220
rect 2924 46180 2930 46192
rect 289262 46180 289268 46192
rect 289320 46180 289326 46232
rect 340874 46180 340880 46232
rect 340932 46220 340938 46232
rect 494146 46220 494152 46232
rect 340932 46192 494152 46220
rect 340932 46180 340938 46192
rect 494146 46180 494152 46192
rect 494204 46180 494210 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 22738 45540 22744 45552
rect 3476 45512 22744 45540
rect 3476 45500 3482 45512
rect 22738 45500 22744 45512
rect 22796 45500 22802 45552
rect 67174 45500 67180 45552
rect 67232 45540 67238 45552
rect 320174 45540 320180 45552
rect 67232 45512 320180 45540
rect 67232 45500 67238 45512
rect 320174 45500 320180 45512
rect 320232 45500 320238 45552
rect 362954 45500 362960 45552
rect 363012 45540 363018 45552
rect 498194 45540 498200 45552
rect 363012 45512 498200 45540
rect 363012 45500 363018 45512
rect 498194 45500 498200 45512
rect 498252 45500 498258 45552
rect 338850 45432 338856 45484
rect 338908 45472 338914 45484
rect 422294 45472 422300 45484
rect 338908 45444 422300 45472
rect 338908 45432 338914 45444
rect 422294 45432 422300 45444
rect 422352 45432 422358 45484
rect 320174 45228 320180 45280
rect 320232 45268 320238 45280
rect 320818 45268 320824 45280
rect 320232 45240 320824 45268
rect 320232 45228 320238 45240
rect 320818 45228 320824 45240
rect 320876 45228 320882 45280
rect 115934 44888 115940 44940
rect 115992 44928 115998 44940
rect 280798 44928 280804 44940
rect 115992 44900 280804 44928
rect 115992 44888 115998 44900
rect 280798 44888 280804 44900
rect 280856 44888 280862 44940
rect 62022 44820 62028 44872
rect 62080 44860 62086 44872
rect 282178 44860 282184 44872
rect 62080 44832 282184 44860
rect 62080 44820 62086 44832
rect 282178 44820 282184 44832
rect 282236 44820 282242 44872
rect 343634 44820 343640 44872
rect 343692 44860 343698 44872
rect 362954 44860 362960 44872
rect 343692 44832 362960 44860
rect 343692 44820 343698 44832
rect 362954 44820 362960 44832
rect 363012 44820 363018 44872
rect 338114 44140 338120 44192
rect 338172 44180 338178 44192
rect 338850 44180 338856 44192
rect 338172 44152 338856 44180
rect 338172 44140 338178 44152
rect 338850 44140 338856 44152
rect 338908 44140 338914 44192
rect 106274 43460 106280 43512
rect 106332 43500 106338 43512
rect 250530 43500 250536 43512
rect 106332 43472 250536 43500
rect 106332 43460 106338 43472
rect 250530 43460 250536 43472
rect 250588 43460 250594 43512
rect 85666 43392 85672 43444
rect 85724 43432 85730 43444
rect 287882 43432 287888 43444
rect 85724 43404 287888 43432
rect 85724 43392 85730 43404
rect 287882 43392 287888 43404
rect 287940 43392 287946 43444
rect 317322 43392 317328 43444
rect 317380 43432 317386 43444
rect 427814 43432 427820 43444
rect 317380 43404 427820 43432
rect 317380 43392 317386 43404
rect 427814 43392 427820 43404
rect 427872 43392 427878 43444
rect 195238 42712 195244 42764
rect 195296 42752 195302 42764
rect 266354 42752 266360 42764
rect 195296 42724 266360 42752
rect 195296 42712 195302 42724
rect 266354 42712 266360 42724
rect 266412 42712 266418 42764
rect 266354 42100 266360 42152
rect 266412 42140 266418 42152
rect 267182 42140 267188 42152
rect 266412 42112 267188 42140
rect 266412 42100 266418 42112
rect 267182 42100 267188 42112
rect 267240 42100 267246 42152
rect 304994 42100 305000 42152
rect 305052 42140 305058 42152
rect 369854 42140 369860 42152
rect 305052 42112 369860 42140
rect 305052 42100 305058 42112
rect 369854 42100 369860 42112
rect 369912 42100 369918 42152
rect 313918 42032 313924 42084
rect 313976 42072 313982 42084
rect 429194 42072 429200 42084
rect 313976 42044 429200 42072
rect 313976 42032 313982 42044
rect 429194 42032 429200 42044
rect 429252 42032 429258 42084
rect 284294 41352 284300 41404
rect 284352 41392 284358 41404
rect 285122 41392 285128 41404
rect 284352 41364 285128 41392
rect 284352 41352 284358 41364
rect 285122 41352 285128 41364
rect 285180 41392 285186 41404
rect 331858 41392 331864 41404
rect 285180 41364 331864 41392
rect 285180 41352 285186 41364
rect 331858 41352 331864 41364
rect 331916 41352 331922 41404
rect 113174 40740 113180 40792
rect 113232 40780 113238 40792
rect 286502 40780 286508 40792
rect 113232 40752 286508 40780
rect 113232 40740 113238 40752
rect 286502 40740 286508 40752
rect 286560 40740 286566 40792
rect 96614 40672 96620 40724
rect 96672 40712 96678 40724
rect 285030 40712 285036 40724
rect 96672 40684 285036 40712
rect 96672 40672 96678 40684
rect 285030 40672 285036 40684
rect 285088 40672 285094 40724
rect 309870 40672 309876 40724
rect 309928 40712 309934 40724
rect 430574 40712 430580 40724
rect 309928 40684 430580 40712
rect 309928 40672 309934 40684
rect 430574 40672 430580 40684
rect 430632 40672 430638 40724
rect 34422 39448 34428 39500
rect 34480 39488 34486 39500
rect 133138 39488 133144 39500
rect 34480 39460 133144 39488
rect 34480 39448 34486 39460
rect 133138 39448 133144 39460
rect 133196 39448 133202 39500
rect 185578 39448 185584 39500
rect 185636 39488 185642 39500
rect 299566 39488 299572 39500
rect 185636 39460 299572 39488
rect 185636 39448 185642 39460
rect 299566 39448 299572 39460
rect 299624 39488 299630 39500
rect 300670 39488 300676 39500
rect 299624 39460 300676 39488
rect 299624 39448 299630 39460
rect 300670 39448 300676 39460
rect 300728 39448 300734 39500
rect 110506 39380 110512 39432
rect 110564 39420 110570 39432
rect 268378 39420 268384 39432
rect 110564 39392 268384 39420
rect 110564 39380 110570 39392
rect 268378 39380 268384 39392
rect 268436 39380 268442 39432
rect 302234 39380 302240 39432
rect 302292 39420 302298 39432
rect 433334 39420 433340 39432
rect 302292 39392 433340 39420
rect 302292 39380 302298 39392
rect 433334 39380 433340 39392
rect 433392 39380 433398 39432
rect 89714 39312 89720 39364
rect 89772 39352 89778 39364
rect 305730 39352 305736 39364
rect 89772 39324 305736 39352
rect 89772 39312 89778 39324
rect 305730 39312 305736 39324
rect 305788 39312 305794 39364
rect 182818 38564 182824 38616
rect 182876 38604 182882 38616
rect 296714 38604 296720 38616
rect 182876 38576 296720 38604
rect 182876 38564 182882 38576
rect 296714 38564 296720 38576
rect 296772 38604 296778 38616
rect 297542 38604 297548 38616
rect 296772 38576 297548 38604
rect 296772 38564 296778 38576
rect 297542 38564 297548 38576
rect 297600 38564 297606 38616
rect 434714 38604 434720 38616
rect 316006 38576 434720 38604
rect 239398 38496 239404 38548
rect 239456 38536 239462 38548
rect 302234 38536 302240 38548
rect 239456 38508 302240 38536
rect 239456 38496 239462 38508
rect 302234 38496 302240 38508
rect 302292 38496 302298 38548
rect 313274 38496 313280 38548
rect 313332 38536 313338 38548
rect 316006 38536 316034 38576
rect 434714 38564 434720 38576
rect 434772 38564 434778 38616
rect 313332 38508 316034 38536
rect 313332 38496 313338 38508
rect 299474 37952 299480 38004
rect 299532 37992 299538 38004
rect 313274 37992 313280 38004
rect 299532 37964 313280 37992
rect 299532 37952 299538 37964
rect 313274 37952 313280 37964
rect 313332 37952 313338 38004
rect 93946 37884 93952 37936
rect 94004 37924 94010 37936
rect 303062 37924 303068 37936
rect 94004 37896 303068 37924
rect 94004 37884 94010 37896
rect 303062 37884 303068 37896
rect 303120 37884 303126 37936
rect 213270 36660 213276 36712
rect 213328 36700 213334 36712
rect 295334 36700 295340 36712
rect 213328 36672 295340 36700
rect 213328 36660 213334 36672
rect 295334 36660 295340 36672
rect 295392 36700 295398 36712
rect 295392 36672 296714 36700
rect 295392 36660 295398 36672
rect 28994 36592 29000 36644
rect 29052 36632 29058 36644
rect 260190 36632 260196 36644
rect 29052 36604 260196 36632
rect 29052 36592 29058 36604
rect 260190 36592 260196 36604
rect 260248 36592 260254 36644
rect 296686 36632 296714 36672
rect 436186 36632 436192 36644
rect 296686 36604 436192 36632
rect 436186 36592 436192 36604
rect 436244 36592 436250 36644
rect 44174 36524 44180 36576
rect 44232 36564 44238 36576
rect 296162 36564 296168 36576
rect 44232 36536 296168 36564
rect 44232 36524 44238 36536
rect 296162 36524 296168 36536
rect 296220 36524 296226 36576
rect 22094 35164 22100 35216
rect 22152 35204 22158 35216
rect 261478 35204 261484 35216
rect 22152 35176 261484 35204
rect 22152 35164 22158 35176
rect 261478 35164 261484 35176
rect 261536 35164 261542 35216
rect 295426 35164 295432 35216
rect 295484 35204 295490 35216
rect 436278 35204 436284 35216
rect 295484 35176 436284 35204
rect 295484 35164 295490 35176
rect 436278 35164 436284 35176
rect 436336 35164 436342 35216
rect 289170 34416 289176 34468
rect 289228 34456 289234 34468
rect 437474 34456 437480 34468
rect 289228 34428 437480 34456
rect 289228 34416 289234 34428
rect 437474 34416 437480 34428
rect 437532 34416 437538 34468
rect 53834 33804 53840 33856
rect 53892 33844 53898 33856
rect 267090 33844 267096 33856
rect 53892 33816 267096 33844
rect 53892 33804 53898 33816
rect 267090 33804 267096 33816
rect 267148 33804 267154 33856
rect 60826 33736 60832 33788
rect 60884 33776 60890 33788
rect 301590 33776 301596 33788
rect 60884 33748 301596 33776
rect 60884 33736 60890 33748
rect 301590 33736 301596 33748
rect 301648 33736 301654 33788
rect 288434 33124 288440 33176
rect 288492 33164 288498 33176
rect 289170 33164 289176 33176
rect 288492 33136 289176 33164
rect 288492 33124 288498 33136
rect 289170 33124 289176 33136
rect 289228 33124 289234 33176
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 47578 33096 47584 33108
rect 3568 33068 47584 33096
rect 3568 33056 3574 33068
rect 47578 33056 47584 33068
rect 47636 33056 47642 33108
rect 184198 33056 184204 33108
rect 184256 33096 184262 33108
rect 313918 33096 313924 33108
rect 184256 33068 313924 33096
rect 184256 33056 184262 33068
rect 313918 33056 313924 33068
rect 313976 33056 313982 33108
rect 327718 33056 327724 33108
rect 327776 33096 327782 33108
rect 425054 33096 425060 33108
rect 327776 33068 425060 33096
rect 327776 33056 327782 33068
rect 425054 33056 425060 33068
rect 425112 33056 425118 33108
rect 99374 32444 99380 32496
rect 99432 32484 99438 32496
rect 265618 32484 265624 32496
rect 99432 32456 265624 32484
rect 99432 32444 99438 32456
rect 265618 32444 265624 32456
rect 265676 32444 265682 32496
rect 291838 32444 291844 32496
rect 291896 32484 291902 32496
rect 293954 32484 293960 32496
rect 291896 32456 293960 32484
rect 291896 32444 291902 32456
rect 293954 32444 293960 32456
rect 294012 32484 294018 32496
rect 360838 32484 360844 32496
rect 294012 32456 360844 32484
rect 294012 32444 294018 32456
rect 360838 32444 360844 32456
rect 360896 32444 360902 32496
rect 103514 32376 103520 32428
rect 103572 32416 103578 32428
rect 294690 32416 294696 32428
rect 103572 32388 294696 32416
rect 103572 32376 103578 32388
rect 294690 32376 294696 32388
rect 294748 32376 294754 32428
rect 313274 32036 313280 32088
rect 313332 32076 313338 32088
rect 313918 32076 313924 32088
rect 313332 32048 313924 32076
rect 313332 32036 313338 32048
rect 313918 32036 313924 32048
rect 313976 32036 313982 32088
rect 327074 31764 327080 31816
rect 327132 31804 327138 31816
rect 327718 31804 327724 31816
rect 327132 31776 327724 31804
rect 327132 31764 327138 31776
rect 327718 31764 327724 31776
rect 327776 31764 327782 31816
rect 238018 31152 238024 31204
rect 238076 31192 238082 31204
rect 284386 31192 284392 31204
rect 238076 31164 284392 31192
rect 238076 31152 238082 31164
rect 284386 31152 284392 31164
rect 284444 31152 284450 31204
rect 100754 31084 100760 31136
rect 100812 31124 100818 31136
rect 302970 31124 302976 31136
rect 100812 31096 302976 31124
rect 100812 31084 100818 31096
rect 302970 31084 302976 31096
rect 303028 31084 303034 31136
rect 19334 31016 19340 31068
rect 19392 31056 19398 31068
rect 271230 31056 271236 31068
rect 19392 31028 271236 31056
rect 19392 31016 19398 31028
rect 271230 31016 271236 31028
rect 271288 31016 271294 31068
rect 284386 31016 284392 31068
rect 284444 31056 284450 31068
rect 438854 31056 438860 31068
rect 284444 31028 438860 31056
rect 284444 31016 284450 31028
rect 438854 31016 438860 31028
rect 438912 31016 438918 31068
rect 175918 30268 175924 30320
rect 175976 30308 175982 30320
rect 241514 30308 241520 30320
rect 175976 30280 241520 30308
rect 175976 30268 175982 30280
rect 241514 30268 241520 30280
rect 241572 30308 241578 30320
rect 242158 30308 242164 30320
rect 241572 30280 242164 30308
rect 241572 30268 241578 30280
rect 242158 30268 242164 30280
rect 242216 30268 242222 30320
rect 277394 30268 277400 30320
rect 277452 30308 277458 30320
rect 278038 30308 278044 30320
rect 277452 30280 278044 30308
rect 277452 30268 277458 30280
rect 278038 30268 278044 30280
rect 278096 30308 278102 30320
rect 441614 30308 441620 30320
rect 278096 30280 441620 30308
rect 278096 30268 278102 30280
rect 441614 30268 441620 30280
rect 441672 30268 441678 30320
rect 82814 29656 82820 29708
rect 82872 29696 82878 29708
rect 282362 29696 282368 29708
rect 82872 29668 282368 29696
rect 82872 29656 82878 29668
rect 282362 29656 282368 29668
rect 282420 29656 282426 29708
rect 95234 29588 95240 29640
rect 95292 29628 95298 29640
rect 295978 29628 295984 29640
rect 95292 29600 295984 29628
rect 95292 29588 95298 29600
rect 295978 29588 295984 29600
rect 296036 29588 296042 29640
rect 246298 28364 246304 28416
rect 246356 28404 246362 28416
rect 274634 28404 274640 28416
rect 246356 28376 274640 28404
rect 246356 28364 246362 28376
rect 274634 28364 274640 28376
rect 274692 28404 274698 28416
rect 274692 28376 277394 28404
rect 274692 28364 274698 28376
rect 44266 28296 44272 28348
rect 44324 28336 44330 28348
rect 272518 28336 272524 28348
rect 44324 28308 272524 28336
rect 44324 28296 44330 28308
rect 272518 28296 272524 28308
rect 272576 28296 272582 28348
rect 277366 28336 277394 28376
rect 442994 28336 443000 28348
rect 277366 28308 443000 28336
rect 442994 28296 443000 28308
rect 443052 28296 443058 28348
rect 59262 28228 59268 28280
rect 59320 28268 59326 28280
rect 298830 28268 298836 28280
rect 59320 28240 298836 28268
rect 59320 28228 59326 28240
rect 298830 28228 298836 28240
rect 298888 28228 298894 28280
rect 188338 27548 188344 27600
rect 188396 27588 188402 27600
rect 329834 27588 329840 27600
rect 188396 27560 329840 27588
rect 188396 27548 188402 27560
rect 329834 27548 329840 27560
rect 329892 27588 329898 27600
rect 330478 27588 330484 27600
rect 329892 27560 330484 27588
rect 329892 27548 329898 27560
rect 330478 27548 330484 27560
rect 330536 27548 330542 27600
rect 39850 27004 39856 27056
rect 39908 27044 39914 27056
rect 128354 27044 128360 27056
rect 39908 27016 128360 27044
rect 39908 27004 39914 27016
rect 128354 27004 128360 27016
rect 128412 27004 128418 27056
rect 118786 26936 118792 26988
rect 118844 26976 118850 26988
rect 276750 26976 276756 26988
rect 118844 26948 276756 26976
rect 118844 26936 118850 26948
rect 276750 26936 276756 26948
rect 276808 26936 276814 26988
rect 276934 26936 276940 26988
rect 276992 26976 276998 26988
rect 444374 26976 444380 26988
rect 276992 26948 444380 26976
rect 276992 26936 276998 26948
rect 444374 26936 444380 26948
rect 444432 26936 444438 26988
rect 92474 26868 92480 26920
rect 92532 26908 92538 26920
rect 283558 26908 283564 26920
rect 92532 26880 283564 26908
rect 92532 26868 92538 26880
rect 283558 26868 283564 26880
rect 283616 26868 283622 26920
rect 271138 26188 271144 26240
rect 271196 26228 271202 26240
rect 276934 26228 276940 26240
rect 271196 26200 276940 26228
rect 271196 26188 271202 26200
rect 276934 26188 276940 26200
rect 276992 26188 276998 26240
rect 204898 25576 204904 25628
rect 204956 25616 204962 25628
rect 267734 25616 267740 25628
rect 204956 25588 267740 25616
rect 204956 25576 204962 25588
rect 267734 25576 267740 25588
rect 267792 25616 267798 25628
rect 445846 25616 445852 25628
rect 267792 25588 445852 25616
rect 267792 25576 267798 25588
rect 445846 25576 445852 25588
rect 445904 25576 445910 25628
rect 77386 25508 77392 25560
rect 77444 25548 77450 25560
rect 276658 25548 276664 25560
rect 77444 25520 276664 25548
rect 77444 25508 77450 25520
rect 276658 25508 276664 25520
rect 276716 25508 276722 25560
rect 81434 24216 81440 24268
rect 81492 24256 81498 24268
rect 282270 24256 282276 24268
rect 81492 24228 282276 24256
rect 81492 24216 81498 24228
rect 282270 24216 282276 24228
rect 282328 24216 282334 24268
rect 57974 24148 57980 24200
rect 58032 24188 58038 24200
rect 264238 24188 264244 24200
rect 58032 24160 264244 24188
rect 58032 24148 58038 24160
rect 264238 24148 264244 24160
rect 264296 24148 264302 24200
rect 264330 24148 264336 24200
rect 264388 24188 264394 24200
rect 445938 24188 445944 24200
rect 264388 24160 445944 24188
rect 264388 24148 264394 24160
rect 445938 24148 445944 24160
rect 445996 24148 446002 24200
rect 52546 24080 52552 24132
rect 52604 24120 52610 24132
rect 304258 24120 304264 24132
rect 52604 24092 304264 24120
rect 52604 24080 52610 24092
rect 304258 24080 304264 24092
rect 304316 24080 304322 24132
rect 244918 22924 244924 22976
rect 244976 22964 244982 22976
rect 262306 22964 262312 22976
rect 244976 22936 262312 22964
rect 244976 22924 244982 22936
rect 262306 22924 262312 22936
rect 262364 22964 262370 22976
rect 447134 22964 447140 22976
rect 262364 22936 447140 22964
rect 262364 22924 262370 22936
rect 447134 22924 447140 22936
rect 447192 22924 447198 22976
rect 111794 22856 111800 22908
rect 111852 22896 111858 22908
rect 302878 22896 302884 22908
rect 111852 22868 302884 22896
rect 111852 22856 111858 22868
rect 302878 22856 302884 22868
rect 302936 22856 302942 22908
rect 46934 22788 46940 22840
rect 46992 22828 46998 22840
rect 262858 22828 262864 22840
rect 46992 22800 262864 22828
rect 46992 22788 46998 22800
rect 262858 22788 262864 22800
rect 262916 22788 262922 22840
rect 63494 22720 63500 22772
rect 63552 22760 63558 22772
rect 289078 22760 289084 22772
rect 63552 22732 289084 22760
rect 63552 22720 63558 22732
rect 289078 22720 289084 22732
rect 289136 22720 289142 22772
rect 253198 22040 253204 22092
rect 253256 22080 253262 22092
rect 449894 22080 449900 22092
rect 253256 22052 449900 22080
rect 253256 22040 253262 22052
rect 449894 22040 449900 22052
rect 449952 22040 449958 22092
rect 252554 21564 252560 21616
rect 252612 21604 252618 21616
rect 253198 21604 253204 21616
rect 252612 21576 253204 21604
rect 252612 21564 252618 21576
rect 253198 21564 253204 21576
rect 253256 21564 253262 21616
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 254578 21468 254584 21480
rect 13872 21440 254584 21468
rect 13872 21428 13878 21440
rect 254578 21428 254584 21440
rect 254636 21428 254642 21480
rect 12434 21360 12440 21412
rect 12492 21400 12498 21412
rect 266998 21400 267004 21412
rect 12492 21372 267004 21400
rect 12492 21360 12498 21372
rect 266998 21360 267004 21372
rect 267056 21360 267062 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 11698 20652 11704 20664
rect 3476 20624 11704 20652
rect 3476 20612 3482 20624
rect 11698 20612 11704 20624
rect 11756 20612 11762 20664
rect 507762 20612 507768 20664
rect 507820 20652 507826 20664
rect 579982 20652 579988 20664
rect 507820 20624 579988 20652
rect 507820 20612 507826 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 250530 20000 250536 20052
rect 250588 20040 250594 20052
rect 451274 20040 451280 20052
rect 250588 20012 451280 20040
rect 250588 20000 250594 20012
rect 451274 20000 451280 20012
rect 451332 20000 451338 20052
rect 49694 19932 49700 19984
rect 49752 19972 49758 19984
rect 294598 19972 294604 19984
rect 49752 19944 294604 19972
rect 49752 19932 49758 19944
rect 294598 19932 294604 19944
rect 294656 19932 294662 19984
rect 298830 19252 298836 19304
rect 298888 19292 298894 19304
rect 359550 19292 359556 19304
rect 298888 19264 359556 19292
rect 298888 19252 298894 19264
rect 359550 19252 359556 19264
rect 359608 19252 359614 19304
rect 75914 18708 75920 18760
rect 75972 18748 75978 18760
rect 269758 18748 269764 18760
rect 75972 18720 269764 18748
rect 75972 18708 75978 18720
rect 269758 18708 269764 18720
rect 269816 18708 269822 18760
rect 246298 18640 246304 18692
rect 246356 18680 246362 18692
rect 452654 18680 452660 18692
rect 246356 18652 452660 18680
rect 246356 18640 246362 18652
rect 452654 18640 452660 18652
rect 452712 18640 452718 18692
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 251818 18612 251824 18624
rect 24912 18584 251824 18612
rect 24912 18572 24918 18584
rect 251818 18572 251824 18584
rect 251876 18572 251882 18624
rect 298094 18028 298100 18080
rect 298152 18068 298158 18080
rect 298830 18068 298836 18080
rect 298152 18040 298836 18068
rect 298152 18028 298158 18040
rect 298830 18028 298836 18040
rect 298888 18028 298894 18080
rect 215938 17280 215944 17332
rect 215996 17320 216002 17332
rect 242986 17320 242992 17332
rect 215996 17292 242992 17320
rect 215996 17280 216002 17292
rect 242986 17280 242992 17292
rect 243044 17320 243050 17332
rect 454126 17320 454132 17332
rect 243044 17292 454132 17320
rect 243044 17280 243050 17292
rect 454126 17280 454132 17292
rect 454184 17280 454190 17332
rect 26234 17212 26240 17264
rect 26292 17252 26298 17264
rect 258718 17252 258724 17264
rect 26292 17224 258724 17252
rect 26292 17212 26298 17224
rect 258718 17212 258724 17224
rect 258776 17212 258782 17264
rect 89162 15988 89168 16040
rect 89220 16028 89226 16040
rect 284938 16028 284944 16040
rect 89220 16000 284944 16028
rect 89220 15988 89226 16000
rect 284938 15988 284944 16000
rect 284996 15988 285002 16040
rect 36722 15920 36728 15972
rect 36780 15960 36786 15972
rect 298738 15960 298744 15972
rect 36780 15932 298744 15960
rect 36780 15920 36786 15932
rect 298738 15920 298744 15932
rect 298796 15920 298802 15972
rect 11882 15852 11888 15904
rect 11940 15892 11946 15904
rect 275278 15892 275284 15904
rect 11940 15864 275284 15892
rect 11940 15852 11946 15864
rect 275278 15852 275284 15864
rect 275336 15852 275342 15904
rect 282270 15852 282276 15904
rect 282328 15892 282334 15904
rect 454034 15892 454040 15904
rect 282328 15864 454040 15892
rect 282328 15852 282334 15864
rect 454034 15852 454040 15864
rect 454092 15852 454098 15904
rect 164418 14492 164424 14544
rect 164476 14532 164482 14544
rect 417418 14532 417424 14544
rect 164476 14504 417424 14532
rect 164476 14492 164482 14504
rect 417418 14492 417424 14504
rect 417476 14492 417482 14544
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 305638 14464 305644 14476
rect 17092 14436 305644 14464
rect 17092 14424 17098 14436
rect 305638 14424 305644 14436
rect 305696 14424 305702 14476
rect 314654 13744 314660 13796
rect 314712 13784 314718 13796
rect 315298 13784 315304 13796
rect 314712 13756 315304 13784
rect 314712 13744 314718 13756
rect 315298 13744 315304 13756
rect 315356 13784 315362 13796
rect 467834 13784 467840 13796
rect 315356 13756 467840 13784
rect 315356 13744 315362 13756
rect 467834 13744 467840 13756
rect 467892 13744 467898 13796
rect 213178 13132 213184 13184
rect 213236 13172 213242 13184
rect 245194 13172 245200 13184
rect 213236 13144 245200 13172
rect 213236 13132 213242 13144
rect 245194 13132 245200 13144
rect 245252 13172 245258 13184
rect 340138 13172 340144 13184
rect 245252 13144 340144 13172
rect 245252 13132 245258 13144
rect 340138 13132 340144 13144
rect 340196 13132 340202 13184
rect 48498 13064 48504 13116
rect 48556 13104 48562 13116
rect 301498 13104 301504 13116
rect 48556 13076 301504 13104
rect 48556 13064 48562 13076
rect 301498 13064 301504 13076
rect 301556 13064 301562 13116
rect 64782 12384 64788 12436
rect 64840 12424 64846 12436
rect 264146 12424 264152 12436
rect 64840 12396 264152 12424
rect 64840 12384 64846 12396
rect 264146 12384 264152 12396
rect 264204 12384 264210 12436
rect 249058 12316 249064 12368
rect 249116 12356 249122 12368
rect 358078 12356 358084 12368
rect 249116 12328 358084 12356
rect 249116 12316 249122 12328
rect 358078 12316 358084 12328
rect 358136 12316 358142 12368
rect 248414 11908 248420 11960
rect 248472 11948 248478 11960
rect 249058 11948 249064 11960
rect 248472 11920 249064 11948
rect 248472 11908 248478 11920
rect 249058 11908 249064 11920
rect 249116 11908 249122 11960
rect 242894 11772 242900 11824
rect 242952 11812 242958 11824
rect 244090 11812 244096 11824
rect 242952 11784 244096 11812
rect 242952 11772 242958 11784
rect 244090 11772 244096 11784
rect 244148 11772 244154 11824
rect 181438 11704 181444 11756
rect 181496 11744 181502 11756
rect 283098 11744 283104 11756
rect 181496 11716 283104 11744
rect 181496 11704 181502 11716
rect 283098 11704 283104 11716
rect 283156 11744 283162 11756
rect 478874 11744 478880 11756
rect 283156 11716 478880 11744
rect 283156 11704 283162 11716
rect 478874 11704 478880 11716
rect 478932 11704 478938 11756
rect 238018 10412 238024 10464
rect 238076 10452 238082 10464
rect 251266 10452 251272 10464
rect 238076 10424 251272 10452
rect 238076 10412 238082 10424
rect 251266 10412 251272 10424
rect 251324 10412 251330 10464
rect 197998 10344 198004 10396
rect 198056 10384 198062 10396
rect 258258 10384 258264 10396
rect 198056 10356 258264 10384
rect 198056 10344 198062 10356
rect 258258 10344 258264 10356
rect 258316 10384 258322 10396
rect 486418 10384 486424 10396
rect 258316 10356 486424 10384
rect 258316 10344 258322 10356
rect 486418 10344 486424 10356
rect 486476 10344 486482 10396
rect 56042 10276 56048 10328
rect 56100 10316 56106 10328
rect 287790 10316 287796 10328
rect 56100 10288 287796 10316
rect 56100 10276 56106 10288
rect 287790 10276 287796 10288
rect 287848 10276 287854 10328
rect 308398 9596 308404 9648
rect 308456 9636 308462 9648
rect 309042 9636 309048 9648
rect 308456 9608 309048 9636
rect 308456 9596 308462 9608
rect 309042 9596 309048 9608
rect 309100 9636 309106 9648
rect 309100 9608 316034 9636
rect 309100 9596 309106 9608
rect 316006 9568 316034 9608
rect 331582 9596 331588 9648
rect 331640 9636 331646 9648
rect 423674 9636 423680 9648
rect 331640 9608 423680 9636
rect 331640 9596 331646 9608
rect 423674 9596 423680 9608
rect 423732 9596 423738 9648
rect 356698 9568 356704 9580
rect 316006 9540 356704 9568
rect 356698 9528 356704 9540
rect 356756 9528 356762 9580
rect 91554 8984 91560 9036
rect 91612 9024 91618 9036
rect 307018 9024 307024 9036
rect 91612 8996 307024 9024
rect 91612 8984 91618 8996
rect 307018 8984 307024 8996
rect 307076 8984 307082 9036
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 29638 8956 29644 8968
rect 3384 8928 29644 8956
rect 3384 8916 3390 8928
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 65518 8916 65524 8968
rect 65576 8956 65582 8968
rect 283650 8956 283656 8968
rect 65576 8928 283656 8956
rect 65576 8916 65582 8928
rect 283650 8916 283656 8928
rect 283708 8916 283714 8968
rect 332594 8848 332600 8900
rect 332652 8888 332658 8900
rect 333882 8888 333888 8900
rect 332652 8860 333888 8888
rect 332652 8848 332658 8860
rect 333882 8848 333888 8860
rect 333940 8848 333946 8900
rect 232498 7692 232504 7744
rect 232556 7732 232562 7744
rect 232556 7704 306374 7732
rect 232556 7692 232562 7704
rect 39942 7624 39948 7676
rect 40000 7664 40006 7676
rect 301498 7664 301504 7676
rect 40000 7636 301504 7664
rect 40000 7624 40006 7636
rect 301498 7624 301504 7636
rect 301556 7624 301562 7676
rect 8754 7556 8760 7608
rect 8812 7596 8818 7608
rect 286410 7596 286416 7608
rect 8812 7568 286416 7596
rect 8812 7556 8818 7568
rect 286410 7556 286416 7568
rect 286468 7556 286474 7608
rect 306346 7596 306374 7704
rect 306742 7596 306748 7608
rect 306346 7568 306748 7596
rect 306742 7556 306748 7568
rect 306800 7596 306806 7608
rect 431954 7596 431960 7608
rect 306800 7568 431960 7596
rect 306800 7556 306806 7568
rect 431954 7556 431960 7568
rect 432012 7556 432018 7608
rect 281902 6808 281908 6860
rect 281960 6848 281966 6860
rect 439498 6848 439504 6860
rect 281960 6820 439504 6848
rect 281960 6808 281966 6820
rect 439498 6808 439504 6820
rect 439556 6808 439562 6860
rect 542998 6808 543004 6860
rect 543056 6848 543062 6860
rect 580166 6848 580172 6860
rect 543056 6820 580172 6848
rect 543056 6808 543062 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 301498 6740 301504 6792
rect 301556 6780 301562 6792
rect 363598 6780 363604 6792
rect 301556 6752 363604 6780
rect 301556 6740 301562 6752
rect 363598 6740 363604 6752
rect 363656 6740 363662 6792
rect 308490 6672 308496 6724
rect 308548 6712 308554 6724
rect 309778 6712 309784 6724
rect 308548 6684 309784 6712
rect 308548 6672 308554 6684
rect 309778 6672 309784 6684
rect 309836 6672 309842 6724
rect 34330 6264 34336 6316
rect 34388 6304 34394 6316
rect 132954 6304 132960 6316
rect 34388 6276 132960 6304
rect 34388 6264 34394 6276
rect 132954 6264 132960 6276
rect 133012 6264 133018 6316
rect 108114 6196 108120 6248
rect 108172 6236 108178 6248
rect 250438 6236 250444 6248
rect 108172 6208 250444 6236
rect 108172 6196 108178 6208
rect 250438 6196 250444 6208
rect 250496 6196 250502 6248
rect 28902 6128 28908 6180
rect 28960 6168 28966 6180
rect 287698 6168 287704 6180
rect 28960 6140 287704 6168
rect 28960 6128 28966 6140
rect 287698 6128 287704 6140
rect 287756 6128 287762 6180
rect 257062 5448 257068 5500
rect 257120 5488 257126 5500
rect 257338 5488 257344 5500
rect 257120 5460 257344 5488
rect 257120 5448 257126 5460
rect 257338 5448 257344 5460
rect 257396 5488 257402 5500
rect 448514 5488 448520 5500
rect 257396 5460 448520 5488
rect 257396 5448 257402 5460
rect 448514 5448 448520 5460
rect 448572 5448 448578 5500
rect 180058 4768 180064 4820
rect 180116 4808 180122 4820
rect 239214 4808 239220 4820
rect 180116 4780 239220 4808
rect 180116 4768 180122 4780
rect 239214 4768 239220 4780
rect 239272 4768 239278 4820
rect 177390 4088 177396 4140
rect 177448 4128 177454 4140
rect 249978 4128 249984 4140
rect 177448 4100 249984 4128
rect 177448 4088 177454 4100
rect 249978 4088 249984 4100
rect 250036 4128 250042 4140
rect 250530 4128 250536 4140
rect 250036 4100 250536 4128
rect 250036 4088 250042 4100
rect 250530 4088 250536 4100
rect 250588 4088 250594 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 333238 4128 333244 4140
rect 332744 4100 333244 4128
rect 332744 4088 332750 4100
rect 333238 4088 333244 4100
rect 333296 4088 333302 4140
rect 346946 4088 346952 4140
rect 347004 4128 347010 4140
rect 352558 4128 352564 4140
rect 347004 4100 352564 4128
rect 347004 4088 347010 4100
rect 352558 4088 352564 4100
rect 352616 4088 352622 4140
rect 191098 4020 191104 4072
rect 191156 4060 191162 4072
rect 246390 4060 246396 4072
rect 191156 4032 246396 4060
rect 191156 4020 191162 4032
rect 246390 4020 246396 4032
rect 246448 4020 246454 4072
rect 239214 3952 239220 4004
rect 239272 3992 239278 4004
rect 282270 3992 282276 4004
rect 239272 3964 282276 3992
rect 239272 3952 239278 3964
rect 282270 3952 282276 3964
rect 282328 3952 282334 4004
rect 109310 3612 109316 3664
rect 109368 3652 109374 3664
rect 173158 3652 173164 3664
rect 109368 3624 173164 3652
rect 109368 3612 109374 3624
rect 173158 3612 173164 3624
rect 173216 3612 173222 3664
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 66772 3556 74534 3584
rect 66772 3544 66778 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 60734 3476 60740 3528
rect 60792 3516 60798 3528
rect 61654 3516 61660 3528
rect 60792 3488 61660 3516
rect 60792 3476 60798 3488
rect 61654 3476 61660 3488
rect 61712 3476 61718 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 74506 3516 74534 3556
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 78214 3584 78220 3596
rect 77352 3556 78220 3584
rect 77352 3544 77358 3556
rect 78214 3544 78220 3556
rect 78272 3544 78278 3596
rect 93854 3544 93860 3596
rect 93912 3584 93918 3596
rect 94774 3584 94780 3596
rect 93912 3556 94780 3584
rect 93912 3544 93918 3556
rect 94774 3544 94780 3556
rect 94832 3544 94838 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 187050 3584 187056 3596
rect 103388 3556 187056 3584
rect 103388 3544 103394 3556
rect 187050 3544 187056 3556
rect 187108 3544 187114 3596
rect 251266 3544 251272 3596
rect 251324 3584 251330 3596
rect 252646 3584 252652 3596
rect 251324 3556 252652 3584
rect 251324 3544 251330 3556
rect 252646 3544 252652 3556
rect 252704 3544 252710 3596
rect 170398 3516 170404 3528
rect 74506 3488 170404 3516
rect 170398 3476 170404 3488
rect 170456 3476 170462 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 252370 3516 252376 3528
rect 251232 3488 252376 3516
rect 251232 3476 251238 3488
rect 252370 3476 252376 3488
rect 252428 3476 252434 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 276842 3516 276848 3528
rect 276072 3488 276848 3516
rect 276072 3476 276078 3488
rect 276842 3476 276848 3488
rect 276900 3476 276906 3528
rect 316678 3476 316684 3528
rect 316736 3516 316742 3528
rect 317322 3516 317328 3528
rect 316736 3488 317328 3516
rect 316736 3476 316742 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 329190 3476 329196 3528
rect 329248 3516 329254 3528
rect 331306 3516 331312 3528
rect 329248 3488 331312 3516
rect 329248 3476 329254 3488
rect 331306 3476 331312 3488
rect 331364 3476 331370 3528
rect 349798 3476 349804 3528
rect 349856 3516 349862 3528
rect 350442 3516 350448 3528
rect 349856 3488 350448 3516
rect 349856 3476 349862 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 17218 3448 17224 3460
rect 6512 3420 17224 3448
rect 6512 3408 6518 3420
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 178678 3448 178684 3460
rect 24268 3420 178684 3448
rect 24268 3408 24274 3420
rect 178678 3408 178684 3420
rect 178736 3408 178742 3460
rect 324406 3408 324412 3460
rect 324464 3448 324470 3460
rect 345750 3448 345756 3460
rect 324464 3420 345756 3448
rect 324464 3408 324470 3420
rect 345750 3408 345756 3420
rect 345808 3408 345814 3460
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 133138 3340 133144 3392
rect 133196 3380 133202 3392
rect 136450 3380 136456 3392
rect 133196 3352 136456 3380
rect 133196 3340 133202 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 260650 3272 260656 3324
rect 260708 3312 260714 3324
rect 262306 3312 262312 3324
rect 260708 3284 262312 3312
rect 260708 3272 260714 3284
rect 262306 3272 262312 3284
rect 262364 3272 262370 3324
rect 235810 3068 235816 3120
rect 235868 3108 235874 3120
rect 238018 3108 238024 3120
rect 235868 3080 238024 3108
rect 235868 3068 235874 3080
rect 238018 3068 238024 3080
rect 238076 3068 238082 3120
rect 292574 3068 292580 3120
rect 292632 3108 292638 3120
rect 295426 3108 295432 3120
rect 292632 3080 295432 3108
rect 292632 3068 292638 3080
rect 295426 3068 295432 3080
rect 295484 3068 295490 3120
rect 171962 3000 171968 3052
rect 172020 3040 172026 3052
rect 177298 3040 177304 3052
rect 172020 3012 177304 3040
rect 172020 3000 172026 3012
rect 177298 3000 177304 3012
rect 177356 3000 177362 3052
rect 35986 2048 35992 2100
rect 36044 2088 36050 2100
rect 297358 2088 297364 2100
rect 36044 2060 297364 2088
rect 36044 2048 36050 2060
rect 297358 2048 297364 2060
rect 297416 2048 297422 2100
<< via1 >>
rect 201500 703332 201552 703384
rect 202788 703332 202840 703384
rect 77944 703264 77996 703316
rect 267648 703264 267700 703316
rect 95148 703196 95200 703248
rect 332508 703196 332560 703248
rect 109684 703128 109736 703180
rect 348792 703128 348844 703180
rect 115204 703060 115256 703112
rect 397460 703060 397512 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 76564 702992 76616 703044
rect 358728 702992 358780 703044
rect 364984 702992 365036 703044
rect 104808 702924 104860 702976
rect 413652 702924 413704 702976
rect 111708 702856 111760 702908
rect 462320 702856 462372 702908
rect 75184 702788 75236 702840
rect 429200 702788 429252 702840
rect 429844 702788 429896 702840
rect 117228 702720 117280 702772
rect 478512 702720 478564 702772
rect 113088 702652 113140 702704
rect 425704 702652 425756 702704
rect 492588 702652 492640 702704
rect 494796 702652 494848 702704
rect 79324 702584 79376 702636
rect 527180 702584 527232 702636
rect 108948 702516 109000 702568
rect 521568 702516 521620 702568
rect 550548 702516 550600 702568
rect 559656 702516 559708 702568
rect 68928 702448 68980 702500
rect 543464 702448 543516 702500
rect 519544 700952 519596 701004
rect 521568 700952 521620 701004
rect 137284 700408 137336 700460
rect 69020 700340 69072 700392
rect 137836 700340 137888 700392
rect 154120 700340 154172 700392
rect 62028 700272 62080 700324
rect 235172 700272 235224 700324
rect 238024 700272 238076 700324
rect 283840 700272 283892 700324
rect 425704 700272 425756 700324
rect 492588 700272 492640 700324
rect 521568 700272 521620 700324
rect 550548 700272 550600 700324
rect 99288 698912 99340 698964
rect 218980 698912 219032 698964
rect 24308 697620 24360 697672
rect 106280 697620 106332 697672
rect 57888 697552 57940 697604
rect 170312 697552 170364 697604
rect 334624 696940 334676 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 15844 683136 15896 683188
rect 320824 683136 320876 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 54484 670692 54536 670744
rect 3424 656888 3476 656940
rect 87604 656888 87656 656940
rect 159364 643084 159416 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 276664 630640 276716 630692
rect 579988 630640 580040 630692
rect 126244 616836 126296 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 35164 605820 35216 605872
rect 6920 598204 6972 598256
rect 53104 598204 53156 598256
rect 53104 597524 53156 597576
rect 85580 597524 85632 597576
rect 15844 596776 15896 596828
rect 50988 596776 51040 596828
rect 50988 596164 51040 596216
rect 71872 596164 71924 596216
rect 68836 594056 68888 594108
rect 238024 594056 238076 594108
rect 81808 592628 81860 592680
rect 580264 592628 580316 592680
rect 40040 592016 40092 592068
rect 48228 592016 48280 592068
rect 74632 592016 74684 592068
rect 580264 592016 580316 592068
rect 582380 592016 582432 592068
rect 385684 590656 385736 590708
rect 579804 590656 579856 590708
rect 3424 588548 3476 588600
rect 57704 588548 57756 588600
rect 88340 588548 88392 588600
rect 118884 588548 118936 588600
rect 57704 587868 57756 587920
rect 95424 587868 95476 587920
rect 97908 586780 97960 586832
rect 113364 586780 113416 586832
rect 52368 586712 52420 586764
rect 85120 586712 85172 586764
rect 100576 586712 100628 586764
rect 121644 586712 121696 586764
rect 49608 586644 49660 586696
rect 81900 586644 81952 586696
rect 92848 586644 92900 586696
rect 117320 586644 117372 586696
rect 48044 586576 48096 586628
rect 84292 586576 84344 586628
rect 94872 586576 94924 586628
rect 123116 586576 123168 586628
rect 42616 586508 42668 586560
rect 80612 586508 80664 586560
rect 89628 586508 89680 586560
rect 123024 586508 123076 586560
rect 68468 585760 68520 585812
rect 137284 585760 137336 585812
rect 99288 585420 99340 585472
rect 109040 585420 109092 585472
rect 87604 585352 87656 585404
rect 110696 585352 110748 585404
rect 53656 585284 53708 585336
rect 74908 585284 74960 585336
rect 94136 585284 94188 585336
rect 46756 585216 46808 585268
rect 83188 585216 83240 585268
rect 41236 585148 41288 585200
rect 78036 585148 78088 585200
rect 98736 585148 98788 585200
rect 99288 585148 99340 585200
rect 118792 585148 118844 585200
rect 103152 584400 103204 584452
rect 104808 584400 104860 584452
rect 112076 584400 112128 584452
rect 55128 584060 55180 584112
rect 73344 584060 73396 584112
rect 45468 583992 45520 584044
rect 78680 583992 78732 584044
rect 88984 583992 89036 584044
rect 111984 583992 112036 584044
rect 59176 583924 59228 583976
rect 76564 583924 76616 583976
rect 77852 583924 77904 583976
rect 79324 583924 79376 583976
rect 101312 583924 101364 583976
rect 113272 583924 113324 583976
rect 70308 583856 70360 583908
rect 83004 583856 83056 583908
rect 103888 583856 103940 583908
rect 120172 583856 120224 583908
rect 47952 583788 48004 583840
rect 77852 583788 77904 583840
rect 96528 583788 96580 583840
rect 118700 583788 118752 583840
rect 65892 583720 65944 583772
rect 70952 583720 71004 583772
rect 105544 583720 105596 583772
rect 114560 583720 114612 583772
rect 56416 582972 56468 583024
rect 71780 582972 71832 583024
rect 92296 582632 92348 582684
rect 110512 582632 110564 582684
rect 70216 582564 70268 582616
rect 84476 582564 84528 582616
rect 97448 582564 97500 582616
rect 116032 582564 116084 582616
rect 50804 582496 50856 582548
rect 76748 582496 76800 582548
rect 99288 582496 99340 582548
rect 120080 582496 120132 582548
rect 3424 582428 3476 582480
rect 107660 582428 107712 582480
rect 69112 582360 69164 582412
rect 580172 582360 580224 582412
rect 65524 581680 65576 581732
rect 75460 581680 75512 581732
rect 79324 581680 79376 581732
rect 90272 581680 90324 581732
rect 39764 581204 39816 581256
rect 67640 581204 67692 581256
rect 59084 581136 59136 581188
rect 43812 581068 43864 581120
rect 65524 581068 65576 581120
rect 37004 581000 37056 581052
rect 70400 581000 70452 581052
rect 104440 581680 104492 581732
rect 104992 581680 105044 581732
rect 114652 581136 114704 581188
rect 126980 581068 127032 581120
rect 121460 581000 121512 581052
rect 108948 579708 109000 579760
rect 128360 579708 128412 579760
rect 3332 579640 3384 579692
rect 15844 579640 15896 579692
rect 52184 579640 52236 579692
rect 69020 579640 69072 579692
rect 57244 578212 57296 578264
rect 67640 578212 67692 578264
rect 108948 578212 109000 578264
rect 134156 578212 134208 578264
rect 356704 577464 356756 577516
rect 429200 577464 429252 577516
rect 108948 576852 109000 576904
rect 129832 576852 129884 576904
rect 108764 575560 108816 575612
rect 131120 575560 131172 575612
rect 34428 575492 34480 575544
rect 67640 575492 67692 575544
rect 108948 575492 109000 575544
rect 122748 575492 122800 575544
rect 429844 575492 429896 575544
rect 59268 574064 59320 574116
rect 67640 574064 67692 574116
rect 108948 574064 109000 574116
rect 124220 574064 124272 574116
rect 65984 573316 66036 573368
rect 68100 573316 68152 573368
rect 108672 573316 108724 573368
rect 130384 573316 130436 573368
rect 61844 572704 61896 572756
rect 67640 572704 67692 572756
rect 64696 571956 64748 572008
rect 67824 571956 67876 572008
rect 105636 571956 105688 572008
rect 110604 571956 110656 572008
rect 108948 571344 109000 571396
rect 133880 571344 133932 571396
rect 108948 569984 109000 570036
rect 120264 569984 120316 570036
rect 41328 569916 41380 569968
rect 67640 569916 67692 569968
rect 108856 569916 108908 569968
rect 142160 569916 142212 569968
rect 64604 568624 64656 568676
rect 67732 568624 67784 568676
rect 61752 568556 61804 568608
rect 67640 568556 67692 568608
rect 108948 568556 109000 568608
rect 129004 568556 129056 568608
rect 106924 567808 106976 567860
rect 117412 567808 117464 567860
rect 66076 567264 66128 567316
rect 67732 567264 67784 567316
rect 108948 567264 109000 567316
rect 117964 567264 118016 567316
rect 63224 567196 63276 567248
rect 67640 567196 67692 567248
rect 108856 567196 108908 567248
rect 125876 567196 125928 567248
rect 108948 565904 109000 565956
rect 113180 565904 113232 565956
rect 3240 565836 3292 565888
rect 25504 565836 25556 565888
rect 64788 565836 64840 565888
rect 67640 565836 67692 565888
rect 108396 565836 108448 565888
rect 111892 565836 111944 565888
rect 429844 565088 429896 565140
rect 497464 565088 497516 565140
rect 504364 565088 504416 565140
rect 41144 564476 41196 564528
rect 67640 564476 67692 564528
rect 108948 564476 109000 564528
rect 123208 564476 123260 564528
rect 108856 564408 108908 564460
rect 133144 564408 133196 564460
rect 155224 564408 155276 564460
rect 108948 564340 109000 564392
rect 117228 564340 117280 564392
rect 117228 563660 117280 563712
rect 138020 563660 138072 563712
rect 504364 563660 504416 563712
rect 580172 563660 580224 563712
rect 49424 563048 49476 563100
rect 67640 563048 67692 563100
rect 61108 562300 61160 562352
rect 62028 562300 62080 562352
rect 67640 562300 67692 562352
rect 60372 561688 60424 561740
rect 67640 561688 67692 561740
rect 56508 561620 56560 561672
rect 61108 561620 61160 561672
rect 60464 560328 60516 560380
rect 67732 560328 67784 560380
rect 108948 560328 109000 560380
rect 116124 560328 116176 560380
rect 57796 560260 57848 560312
rect 67640 560260 67692 560312
rect 108212 560260 108264 560312
rect 140780 560260 140832 560312
rect 136640 559512 136692 559564
rect 201500 559512 201552 559564
rect 108948 558968 109000 559020
rect 135444 558968 135496 559020
rect 42708 558900 42760 558952
rect 67640 558900 67692 558952
rect 108856 558900 108908 558952
rect 136640 558900 136692 558952
rect 66168 558288 66220 558340
rect 68836 558288 68888 558340
rect 56324 557540 56376 557592
rect 67640 557540 67692 557592
rect 108948 557540 109000 557592
rect 115940 557540 115992 557592
rect 108948 556520 109000 556572
rect 113916 556520 113968 556572
rect 43720 556248 43772 556300
rect 67640 556248 67692 556300
rect 37096 556180 37148 556232
rect 67824 556180 67876 556232
rect 55036 556112 55088 556164
rect 57888 556112 57940 556164
rect 67732 556112 67784 556164
rect 108948 556112 109000 556164
rect 110604 556112 110656 556164
rect 110604 555432 110656 555484
rect 116584 555432 116636 555484
rect 37188 554752 37240 554804
rect 67640 554752 67692 554804
rect 141516 554004 141568 554056
rect 159364 554004 159416 554056
rect 108856 553460 108908 553512
rect 118976 553460 119028 553512
rect 50896 553392 50948 553444
rect 67640 553392 67692 553444
rect 108948 553392 109000 553444
rect 141516 553392 141568 553444
rect 142068 553392 142120 553444
rect 53748 552032 53800 552084
rect 67640 552032 67692 552084
rect 108948 552032 109000 552084
rect 124588 552032 124640 552084
rect 107844 551488 107896 551540
rect 110604 551488 110656 551540
rect 38568 550604 38620 550656
rect 67640 550604 67692 550656
rect 108948 550604 109000 550656
rect 138112 550604 138164 550656
rect 108948 549312 109000 549364
rect 132500 549312 132552 549364
rect 35716 549244 35768 549296
rect 67640 549244 67692 549296
rect 108856 549244 108908 549296
rect 142252 549244 142304 549296
rect 52276 547952 52328 548004
rect 67640 547952 67692 548004
rect 39856 547884 39908 547936
rect 67732 547884 67784 547936
rect 61936 546524 61988 546576
rect 67732 546524 67784 546576
rect 60648 546456 60700 546508
rect 67640 546456 67692 546508
rect 108948 546456 109000 546508
rect 135260 546456 135312 546508
rect 108948 545708 109000 545760
rect 113088 545708 113140 545760
rect 125784 545708 125836 545760
rect 110420 545164 110472 545216
rect 111708 545164 111760 545216
rect 133972 545164 134024 545216
rect 35808 545096 35860 545148
rect 68560 545096 68612 545148
rect 108948 545096 109000 545148
rect 139492 545096 139544 545148
rect 108856 545028 108908 545080
rect 110420 545028 110472 545080
rect 25504 544348 25556 544400
rect 68008 544348 68060 544400
rect 63408 542444 63460 542496
rect 67640 542444 67692 542496
rect 46848 542376 46900 542428
rect 67732 542376 67784 542428
rect 108948 542376 109000 542428
rect 136732 542376 136784 542428
rect 129740 541628 129792 541680
rect 299480 541628 299532 541680
rect 109776 541016 109828 541068
rect 129740 541016 129792 541068
rect 63316 540948 63368 541000
rect 67640 540948 67692 541000
rect 108948 540948 109000 541000
rect 142344 540948 142396 541000
rect 107476 540880 107528 540932
rect 109684 540880 109736 540932
rect 62028 539588 62080 539640
rect 67640 539588 67692 539640
rect 4804 539520 4856 539572
rect 99012 539520 99064 539572
rect 95148 539112 95200 539164
rect 118792 539112 118844 539164
rect 97908 539044 97960 539096
rect 113364 539044 113416 539096
rect 59084 538976 59136 539028
rect 73160 538976 73212 539028
rect 88064 538976 88116 539028
rect 118792 538976 118844 539028
rect 126244 538976 126296 539028
rect 57704 538908 57756 538960
rect 90364 538908 90416 538960
rect 98644 538908 98696 538960
rect 120172 538908 120224 538960
rect 54484 538840 54536 538892
rect 57888 538840 57940 538892
rect 91284 538840 91336 538892
rect 99012 538840 99064 538892
rect 124496 538840 124548 538892
rect 15844 538160 15896 538212
rect 98368 538160 98420 538212
rect 103520 538160 103572 538212
rect 109776 538160 109828 538212
rect 155224 538160 155276 538212
rect 580172 538160 580224 538212
rect 102232 537752 102284 537804
rect 110788 537752 110840 537804
rect 70308 537684 70360 537736
rect 81532 537684 81584 537736
rect 102876 537684 102928 537736
rect 127624 537684 127676 537736
rect 45376 537616 45428 537668
rect 56416 537616 56468 537668
rect 57704 537616 57756 537668
rect 81624 537616 81676 537668
rect 83464 537616 83516 537668
rect 90640 537616 90692 537668
rect 98368 537616 98420 537668
rect 122932 537616 122984 537668
rect 44088 537548 44140 537600
rect 73252 537548 73304 537600
rect 79692 537548 79744 537600
rect 87052 537548 87104 537600
rect 95792 537548 95844 537600
rect 121552 537548 121604 537600
rect 52092 537480 52144 537532
rect 82912 537480 82964 537532
rect 84200 537480 84252 537532
rect 98552 537480 98604 537532
rect 100300 537480 100352 537532
rect 132592 537480 132644 537532
rect 94504 537412 94556 537464
rect 100760 537412 100812 537464
rect 70216 536800 70268 536852
rect 75092 536800 75144 536852
rect 84108 536800 84160 536852
rect 84844 536800 84896 536852
rect 102048 536800 102100 536852
rect 104164 536800 104216 536852
rect 35164 536732 35216 536784
rect 106280 536732 106332 536784
rect 100760 536664 100812 536716
rect 118884 536664 118936 536716
rect 97816 536120 97868 536172
rect 110512 536120 110564 536172
rect 118884 536120 118936 536172
rect 128544 536120 128596 536172
rect 106280 536052 106332 536104
rect 131212 536052 131264 536104
rect 71044 535372 71096 535424
rect 77116 535372 77168 535424
rect 48136 534828 48188 534880
rect 75184 534828 75236 534880
rect 99288 534828 99340 534880
rect 114652 534828 114704 534880
rect 115204 534828 115256 534880
rect 128360 534828 128412 534880
rect 53564 534760 53616 534812
rect 83556 534760 83608 534812
rect 93860 534760 93912 534812
rect 120172 534760 120224 534812
rect 46572 534692 46624 534744
rect 78404 534692 78456 534744
rect 89996 534692 90048 534744
rect 118884 534692 118936 534744
rect 46756 533332 46808 533384
rect 76564 533332 76616 533384
rect 49516 532108 49568 532160
rect 76472 532108 76524 532160
rect 97080 532108 97132 532160
rect 121736 532108 121788 532160
rect 52368 532040 52420 532092
rect 79324 532040 79376 532092
rect 87420 532040 87472 532092
rect 109224 532040 109276 532092
rect 54944 531972 54996 532024
rect 86132 531972 86184 532024
rect 95056 531972 95108 532024
rect 121644 531972 121696 532024
rect 56416 529320 56468 529372
rect 72608 529320 72660 529372
rect 46664 529252 46716 529304
rect 70492 529252 70544 529304
rect 40960 529184 41012 529236
rect 74540 529184 74592 529236
rect 110420 529184 110472 529236
rect 110604 529184 110656 529236
rect 128360 529184 128412 529236
rect 3148 528504 3200 528556
rect 110420 528572 110472 528624
rect 39672 526396 39724 526448
rect 71964 526396 72016 526448
rect 34244 525784 34296 525836
rect 69020 525716 69072 525768
rect 579804 525716 579856 525768
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 431224 510620 431276 510672
rect 580172 510620 580224 510672
rect 88248 500284 88300 500336
rect 117412 500284 117464 500336
rect 125600 500284 125652 500336
rect 95240 500216 95292 500268
rect 136824 500216 136876 500268
rect 137100 500216 137152 500268
rect 89352 498788 89404 498840
rect 111800 498788 111852 498840
rect 85488 497564 85540 497616
rect 109316 497564 109368 497616
rect 84108 497496 84160 497548
rect 110420 497496 110472 497548
rect 38476 497428 38528 497480
rect 70400 497428 70452 497480
rect 81624 497428 81676 497480
rect 88248 497428 88300 497480
rect 96436 497428 96488 497480
rect 131304 497428 131356 497480
rect 88064 496272 88116 496324
rect 123116 496272 123168 496324
rect 89628 496204 89680 496256
rect 125692 496204 125744 496256
rect 127072 496204 127124 496256
rect 76472 496136 76524 496188
rect 81532 496136 81584 496188
rect 123300 496136 123352 496188
rect 4804 496068 4856 496120
rect 91100 496068 91152 496120
rect 135352 496068 135404 496120
rect 91100 495456 91152 495508
rect 116032 495456 116084 495508
rect 116400 495456 116452 495508
rect 93216 494980 93268 495032
rect 112168 494980 112220 495032
rect 58992 494844 59044 494896
rect 80980 494844 81032 494896
rect 82268 494844 82320 494896
rect 111984 494844 112036 494896
rect 119068 494844 119120 494896
rect 43904 494776 43956 494828
rect 49608 494776 49660 494828
rect 75460 494776 75512 494828
rect 82912 494776 82964 494828
rect 123024 494776 123076 494828
rect 127256 494776 127308 494828
rect 3516 494708 3568 494760
rect 82820 494708 82872 494760
rect 90640 494708 90692 494760
rect 118700 494708 118752 494760
rect 134064 494708 134116 494760
rect 47860 494504 47912 494556
rect 48044 494504 48096 494556
rect 47860 494028 47912 494080
rect 77392 494028 77444 494080
rect 82820 493960 82872 494012
rect 83556 493960 83608 494012
rect 121460 493960 121512 494012
rect 120080 493892 120132 493944
rect 121828 493892 121880 493944
rect 88708 493824 88760 493876
rect 89536 493824 89588 493876
rect 110512 493552 110564 493604
rect 110696 493552 110748 493604
rect 124404 493552 124456 493604
rect 97724 493484 97776 493536
rect 114744 493484 114796 493536
rect 95148 493416 95200 493468
rect 113272 493416 113324 493468
rect 93216 493348 93268 493400
rect 54760 493280 54812 493332
rect 59176 493280 59228 493332
rect 70032 493280 70084 493332
rect 80980 493280 81032 493332
rect 110512 493280 110564 493332
rect 121460 493348 121512 493400
rect 128452 493348 128504 493400
rect 137284 493280 137336 493332
rect 120080 493212 120132 493264
rect 85488 493144 85540 493196
rect 89628 493144 89680 493196
rect 47952 492668 48004 492720
rect 71136 492668 71188 492720
rect 88708 492668 88760 492720
rect 102140 492668 102192 492720
rect 75184 492600 75236 492652
rect 78404 492600 78456 492652
rect 39948 492056 40000 492108
rect 45468 492056 45520 492108
rect 72240 492056 72292 492108
rect 49608 491988 49660 492040
rect 53104 491988 53156 492040
rect 80060 491988 80112 492040
rect 91928 491988 91980 492040
rect 97908 491988 97960 492040
rect 101404 491988 101456 492040
rect 56232 491920 56284 491972
rect 83464 491920 83516 491972
rect 86132 491920 86184 491972
rect 96988 491920 97040 491972
rect 98368 491920 98420 491972
rect 126980 491920 127032 491972
rect 139400 491920 139452 491972
rect 78404 491648 78456 491700
rect 103612 491648 103664 491700
rect 76656 491580 76708 491632
rect 113272 491580 113324 491632
rect 99656 491512 99708 491564
rect 114560 491512 114612 491564
rect 90364 491444 90416 491496
rect 110604 491444 110656 491496
rect 58624 491376 58676 491428
rect 70400 491376 70452 491428
rect 86776 491376 86828 491428
rect 92480 491376 92532 491428
rect 41236 491308 41288 491360
rect 71780 491308 71832 491360
rect 50804 491240 50856 491292
rect 58624 491240 58676 491292
rect 107568 491240 107620 491292
rect 109040 491240 109092 491292
rect 116400 491240 116452 491292
rect 120080 491240 120132 491292
rect 120356 491172 120408 491224
rect 87420 490696 87472 490748
rect 95056 490696 95108 490748
rect 100024 490696 100076 490748
rect 92848 490628 92900 490680
rect 107568 490628 107620 490680
rect 50804 490560 50856 490612
rect 79048 490560 79100 490612
rect 92020 490560 92072 490612
rect 109408 490560 109460 490612
rect 42616 489948 42668 490000
rect 74356 489948 74408 490000
rect 45284 489880 45336 489932
rect 73436 489880 73488 489932
rect 43812 489812 43864 489864
rect 69020 489812 69072 489864
rect 98000 489812 98052 489864
rect 98644 489812 98696 489864
rect 99196 489812 99248 489864
rect 101220 489812 101272 489864
rect 117320 489812 117372 489864
rect 102232 489268 102284 489320
rect 115204 489268 115256 489320
rect 99196 489200 99248 489252
rect 113824 489200 113876 489252
rect 106188 489132 106240 489184
rect 134156 489132 134208 489184
rect 151820 489132 151872 489184
rect 53656 488452 53708 488504
rect 67640 488452 67692 488504
rect 102324 488452 102376 488504
rect 109132 488452 109184 488504
rect 102232 488044 102284 488096
rect 106188 488044 106240 488096
rect 48228 487772 48280 487824
rect 67640 487772 67692 487824
rect 109132 487772 109184 487824
rect 116032 487772 116084 487824
rect 55128 487092 55180 487144
rect 68008 487092 68060 487144
rect 102232 487092 102284 487144
rect 129924 487160 129976 487212
rect 99472 485800 99524 485852
rect 141056 485800 141108 485852
rect 103428 485052 103480 485104
rect 111984 485052 112036 485104
rect 67640 484372 67692 484424
rect 286324 484372 286376 484424
rect 580172 484372 580224 484424
rect 50988 484304 51040 484356
rect 53104 484304 53156 484356
rect 37004 483624 37056 483676
rect 65892 483624 65944 483676
rect 67640 483624 67692 483676
rect 103428 483624 103480 483676
rect 122840 483624 122892 483676
rect 123392 483624 123444 483676
rect 39764 482944 39816 482996
rect 68100 482944 68152 482996
rect 115204 482944 115256 482996
rect 117412 482944 117464 482996
rect 67364 482400 67416 482452
rect 69848 482400 69900 482452
rect 36912 482264 36964 482316
rect 66904 482264 66956 482316
rect 67456 482264 67508 482316
rect 103428 482264 103480 482316
rect 114560 482264 114612 482316
rect 106280 481788 106332 481840
rect 107016 481788 107068 481840
rect 103336 481720 103388 481772
rect 110328 481720 110380 481772
rect 129832 481720 129884 481772
rect 130384 481720 130436 481772
rect 143724 481720 143776 481772
rect 146300 481652 146352 481704
rect 52184 481584 52236 481636
rect 69112 481584 69164 481636
rect 103428 481584 103480 481636
rect 129832 481584 129884 481636
rect 103336 481516 103388 481568
rect 106280 481516 106332 481568
rect 110328 481516 110380 481568
rect 124220 481516 124272 481568
rect 54852 480224 54904 480276
rect 57244 480224 57296 480276
rect 67640 480156 67692 480208
rect 103336 479544 103388 479596
rect 107660 479544 107712 479596
rect 115204 479544 115256 479596
rect 103428 479476 103480 479528
rect 133880 479476 133932 479528
rect 64420 478864 64472 478916
rect 65800 478864 65852 478916
rect 105636 478864 105688 478916
rect 109224 478864 109276 478916
rect 129004 478864 129056 478916
rect 129832 478864 129884 478916
rect 60556 478796 60608 478848
rect 67272 478796 67324 478848
rect 103428 477504 103480 477556
rect 108948 477436 109000 477488
rect 142160 477436 142212 477488
rect 103336 476824 103388 476876
rect 125876 476824 125928 476876
rect 105176 476756 105228 476808
rect 129832 476756 129884 476808
rect 34336 476076 34388 476128
rect 67640 476076 67692 476128
rect 117964 476076 118016 476128
rect 124312 476076 124364 476128
rect 103244 476008 103296 476060
rect 120264 476008 120316 476060
rect 102232 475940 102284 475992
rect 117964 475940 118016 475992
rect 102324 475872 102376 475924
rect 111892 475872 111944 475924
rect 112628 475872 112680 475924
rect 59084 475396 59136 475448
rect 67640 475396 67692 475448
rect 35624 475328 35676 475380
rect 65984 475328 66036 475380
rect 67732 475328 67784 475380
rect 112628 475328 112680 475380
rect 122840 475328 122892 475380
rect 3424 474716 3476 474768
rect 11704 474716 11756 474768
rect 102232 474648 102284 474700
rect 113180 474648 113232 474700
rect 115480 474648 115532 474700
rect 61844 474308 61896 474360
rect 65984 474308 66036 474360
rect 67640 474308 67692 474360
rect 42616 473356 42668 473408
rect 53840 473356 53892 473408
rect 64696 473288 64748 473340
rect 67640 473288 67692 473340
rect 102232 473288 102284 473340
rect 133144 473288 133196 473340
rect 133788 473288 133840 473340
rect 52184 472608 52236 472660
rect 64696 472608 64748 472660
rect 102232 472608 102284 472660
rect 123208 472608 123260 472660
rect 124128 472608 124180 472660
rect 133788 472608 133840 472660
rect 142160 472608 142212 472660
rect 102324 471996 102376 472048
rect 103428 471996 103480 472048
rect 146392 471996 146444 472048
rect 124128 471248 124180 471300
rect 145012 471248 145064 471300
rect 41328 470500 41380 470552
rect 61384 470568 61436 470620
rect 67640 470568 67692 470620
rect 102232 470568 102284 470620
rect 64604 470500 64656 470552
rect 65984 470500 66036 470552
rect 67732 470500 67784 470552
rect 145012 470568 145064 470620
rect 579988 470568 580040 470620
rect 138020 470500 138072 470552
rect 102232 469888 102284 469940
rect 105544 469888 105596 469940
rect 140964 469888 141016 469940
rect 103612 469820 103664 469872
rect 140780 469820 140832 469872
rect 147864 469820 147916 469872
rect 61752 469548 61804 469600
rect 67640 469548 67692 469600
rect 102232 469208 102284 469260
rect 138020 469208 138072 469260
rect 138204 469208 138256 469260
rect 106188 469140 106240 469192
rect 116124 469140 116176 469192
rect 103612 468460 103664 468512
rect 135444 468460 135496 468512
rect 149152 468460 149204 468512
rect 56324 468324 56376 468376
rect 64144 468324 64196 468376
rect 59268 467848 59320 467900
rect 63224 467848 63276 467900
rect 67640 467848 67692 467900
rect 64788 467780 64840 467832
rect 67456 467780 67508 467832
rect 104164 467100 104216 467152
rect 114836 467100 114888 467152
rect 102232 466488 102284 466540
rect 133788 466488 133840 466540
rect 144920 466420 144972 466472
rect 102324 466352 102376 466404
rect 108304 466352 108356 466404
rect 133788 466352 133840 466404
rect 136640 466352 136692 466404
rect 41052 465672 41104 465724
rect 67640 465672 67692 465724
rect 102232 465672 102284 465724
rect 115940 465672 115992 465724
rect 116860 465672 116912 465724
rect 66076 465332 66128 465384
rect 67548 465332 67600 465384
rect 67916 465332 67968 465384
rect 102232 464992 102284 465044
rect 113916 465060 113968 465112
rect 150624 465060 150676 465112
rect 116860 464992 116912 465044
rect 121644 464992 121696 465044
rect 49424 464312 49476 464364
rect 67640 464312 67692 464364
rect 108304 464312 108356 464364
rect 110788 464312 110840 464364
rect 49424 463632 49476 463684
rect 50344 463632 50396 463684
rect 102232 463632 102284 463684
rect 116584 463632 116636 463684
rect 128636 463700 128688 463752
rect 56508 462952 56560 463004
rect 67640 462952 67692 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 102232 462272 102284 462324
rect 140780 462272 140832 462324
rect 60464 461592 60516 461644
rect 67640 461592 67692 461644
rect 102324 460980 102376 461032
rect 115940 460980 115992 461032
rect 102232 460844 102284 460896
rect 108396 460844 108448 460896
rect 147772 460912 147824 460964
rect 115940 460844 115992 460896
rect 118976 460844 119028 460896
rect 108396 460232 108448 460284
rect 124588 460232 124640 460284
rect 42708 460164 42760 460216
rect 52460 460164 52512 460216
rect 57796 460164 57848 460216
rect 67640 460164 67692 460216
rect 102324 460164 102376 460216
rect 138112 460164 138164 460216
rect 151912 460164 151964 460216
rect 52460 459552 52512 459604
rect 53656 459552 53708 459604
rect 67640 459552 67692 459604
rect 102416 459552 102468 459604
rect 108396 459552 108448 459604
rect 108856 459552 108908 459604
rect 125140 459552 125192 459604
rect 128360 459552 128412 459604
rect 66168 459484 66220 459536
rect 67732 459484 67784 459536
rect 43996 458872 44048 458924
rect 57796 458872 57848 458924
rect 64144 458872 64196 458924
rect 64788 458872 64840 458924
rect 67640 458872 67692 458924
rect 102232 458872 102284 458924
rect 124220 458872 124272 458924
rect 125140 458872 125192 458924
rect 45468 458804 45520 458856
rect 66168 458804 66220 458856
rect 103612 458804 103664 458856
rect 142252 458804 142304 458856
rect 152004 458804 152056 458856
rect 108488 458192 108540 458244
rect 138112 458192 138164 458244
rect 39764 458124 39816 458176
rect 43720 458124 43772 458176
rect 67732 458124 67784 458176
rect 37004 457444 37056 457496
rect 67640 457444 67692 457496
rect 102232 456696 102284 456748
rect 106924 456696 106976 456748
rect 143632 456764 143684 456816
rect 446404 456764 446456 456816
rect 580172 456764 580224 456816
rect 100208 456152 100260 456204
rect 109316 456152 109368 456204
rect 102324 456084 102376 456136
rect 132500 456084 132552 456136
rect 106096 456016 106148 456068
rect 135260 456016 135312 456068
rect 142252 456016 142304 456068
rect 37188 455336 37240 455388
rect 64144 455336 64196 455388
rect 67640 455404 67692 455456
rect 102324 455336 102376 455388
rect 108488 455336 108540 455388
rect 55036 455268 55088 455320
rect 57336 455268 57388 455320
rect 102232 455268 102284 455320
rect 106096 455268 106148 455320
rect 107384 454656 107436 454708
rect 139492 454656 139544 454708
rect 150532 454656 150584 454708
rect 57336 454044 57388 454096
rect 67640 454044 67692 454096
rect 102232 453976 102284 454028
rect 125784 453976 125836 454028
rect 102324 453908 102376 453960
rect 107384 453908 107436 453960
rect 53748 452684 53800 452736
rect 57796 452684 57848 452736
rect 67640 452684 67692 452736
rect 67732 452616 67784 452668
rect 50896 452548 50948 452600
rect 51724 452548 51776 452600
rect 102232 452548 102284 452600
rect 133972 452548 134024 452600
rect 135168 452548 135220 452600
rect 136732 452480 136784 452532
rect 137376 452480 137428 452532
rect 135168 451868 135220 451920
rect 147680 451868 147732 451920
rect 62488 451460 62540 451512
rect 67640 451460 67692 451512
rect 102784 451256 102836 451308
rect 137376 451256 137428 451308
rect 35716 451188 35768 451240
rect 67640 451188 67692 451240
rect 38568 451120 38620 451172
rect 62488 451120 62540 451172
rect 102232 450236 102284 450288
rect 104992 450236 105044 450288
rect 105912 450236 105964 450288
rect 33048 449896 33100 449948
rect 35716 449896 35768 449948
rect 102232 448672 102284 448724
rect 106832 448672 106884 448724
rect 107384 448604 107436 448656
rect 119344 448604 119396 448656
rect 60464 448536 60516 448588
rect 61752 448536 61804 448588
rect 39856 448468 39908 448520
rect 67824 448468 67876 448520
rect 102232 448468 102284 448520
rect 131120 448536 131172 448588
rect 139492 448468 139544 448520
rect 140688 448468 140740 448520
rect 142344 448468 142396 448520
rect 61936 448400 61988 448452
rect 62120 448400 62172 448452
rect 102324 448400 102376 448452
rect 107384 448400 107436 448452
rect 106832 447788 106884 447840
rect 139492 447788 139544 447840
rect 62120 447176 62172 447228
rect 67640 447176 67692 447228
rect 104716 447108 104768 447160
rect 110604 447108 110656 447160
rect 60740 445816 60792 445868
rect 61936 445816 61988 445868
rect 67732 445816 67784 445868
rect 102048 445816 102100 445868
rect 102416 445816 102468 445868
rect 135260 445816 135312 445868
rect 35808 445680 35860 445732
rect 65524 445748 65576 445800
rect 67640 445748 67692 445800
rect 102324 445748 102376 445800
rect 143540 445748 143592 445800
rect 102232 445680 102284 445732
rect 104900 445680 104952 445732
rect 105544 445680 105596 445732
rect 127624 444456 127676 444508
rect 140872 444456 140924 444508
rect 104808 444388 104860 444440
rect 129740 444388 129792 444440
rect 102232 443980 102284 444032
rect 104808 443980 104860 444032
rect 46848 443640 46900 443692
rect 67640 443640 67692 443692
rect 62764 442416 62816 442468
rect 63408 442416 63460 442468
rect 67640 442416 67692 442468
rect 34244 442212 34296 442264
rect 67640 442212 67692 442264
rect 102232 442212 102284 442264
rect 108304 442212 108356 442264
rect 62028 441532 62080 441584
rect 64512 441532 64564 441584
rect 102232 441532 102284 441584
rect 132592 441532 132644 441584
rect 61752 441464 61804 441516
rect 63316 441464 63368 441516
rect 67640 441464 67692 441516
rect 64512 440920 64564 440972
rect 67640 440920 67692 440972
rect 38476 440852 38528 440904
rect 71044 440648 71096 440700
rect 94136 440648 94188 440700
rect 112168 440920 112220 440972
rect 91744 440580 91796 440632
rect 111800 440580 111852 440632
rect 132592 440308 132644 440360
rect 133972 440308 134024 440360
rect 37096 440240 37148 440292
rect 38476 440240 38528 440292
rect 100668 440240 100720 440292
rect 136732 440240 136784 440292
rect 66996 439560 67048 439612
rect 76564 439560 76616 439612
rect 53748 439492 53800 439544
rect 57704 439492 57756 439544
rect 73160 439492 73212 439544
rect 91652 439152 91704 439204
rect 91928 439152 91980 439204
rect 67364 439084 67416 439136
rect 73344 439084 73396 439136
rect 43720 439016 43772 439068
rect 45376 439016 45428 439068
rect 73896 439016 73948 439068
rect 84844 439016 84896 439068
rect 110420 439084 110472 439136
rect 57888 438948 57940 439000
rect 91652 438948 91704 439000
rect 11704 438880 11756 438932
rect 95240 439016 95292 439068
rect 96436 439016 96488 439068
rect 103612 439016 103664 439068
rect 106924 439016 106976 439068
rect 94044 438948 94096 439000
rect 95148 438948 95200 439000
rect 128544 438948 128596 439000
rect 91928 438880 91980 438932
rect 95884 438880 95936 438932
rect 96436 438880 96488 438932
rect 121552 438880 121604 438932
rect 50988 438812 51040 438864
rect 53564 438812 53616 438864
rect 83556 438812 83608 438864
rect 88984 438812 89036 438864
rect 118792 438812 118844 438864
rect 73160 438744 73212 438796
rect 82268 438744 82320 438796
rect 89996 438744 90048 438796
rect 91008 438744 91060 438796
rect 118884 438744 118936 438796
rect 48136 438676 48188 438728
rect 75828 438676 75880 438728
rect 99012 438676 99064 438728
rect 99288 438676 99340 438728
rect 122932 438676 122984 438728
rect 80704 438608 80756 438660
rect 104164 438608 104216 438660
rect 98368 438540 98420 438592
rect 99196 438540 99248 438592
rect 114744 438540 114796 438592
rect 65892 438268 65944 438320
rect 75184 438268 75236 438320
rect 56416 438200 56468 438252
rect 73252 438200 73304 438252
rect 4804 438132 4856 438184
rect 50988 438132 51040 438184
rect 57244 438132 57296 438184
rect 91284 438132 91336 438184
rect 99656 438132 99708 438184
rect 102048 438132 102100 438184
rect 124496 438132 124548 438184
rect 83556 437928 83608 437980
rect 84844 437928 84896 437980
rect 89352 437724 89404 437776
rect 91744 437724 91796 437776
rect 56232 437452 56284 437504
rect 57244 437452 57296 437504
rect 54944 437384 54996 437436
rect 85580 437384 85632 437436
rect 86776 437384 86828 437436
rect 46572 437316 46624 437368
rect 78404 437316 78456 437368
rect 86224 437316 86276 437368
rect 100208 437384 100260 437436
rect 94872 437316 94924 437368
rect 120172 437316 120224 437368
rect 52092 437248 52144 437300
rect 82912 437248 82964 437300
rect 97080 437248 97132 437300
rect 44088 437180 44140 437232
rect 55864 437180 55916 437232
rect 56416 437180 56468 437232
rect 58992 437180 59044 437232
rect 81624 437180 81676 437232
rect 87696 437180 87748 437232
rect 105636 437180 105688 437232
rect 131304 437180 131356 437232
rect 69204 436908 69256 436960
rect 72424 436908 72476 436960
rect 39672 436704 39724 436756
rect 46756 436704 46808 436756
rect 71688 436704 71740 436756
rect 78404 436432 78456 436484
rect 83464 436432 83516 436484
rect 97080 436364 97132 436416
rect 97908 436364 97960 436416
rect 50804 436024 50856 436076
rect 78772 436024 78824 436076
rect 92572 436024 92624 436076
rect 93676 436024 93728 436076
rect 109408 436024 109460 436076
rect 40960 434664 41012 434716
rect 74540 434664 74592 434716
rect 56324 434596 56376 434648
rect 71872 434596 71924 434648
rect 72608 434596 72660 434648
rect 59084 433984 59136 434036
rect 69664 433984 69716 434036
rect 49516 433236 49568 433288
rect 76472 433236 76524 433288
rect 42708 432556 42760 432608
rect 49516 432556 49568 432608
rect 69020 432556 69072 432608
rect 80796 432556 80848 432608
rect 100760 431264 100812 431316
rect 104992 431264 105044 431316
rect 83464 431196 83516 431248
rect 580172 431196 580224 431248
rect 69112 431060 69164 431112
rect 71964 431060 72016 431112
rect 104992 430584 105044 430636
rect 111156 430584 111208 430636
rect 3424 429836 3476 429888
rect 100760 429836 100812 429888
rect 3516 422288 3568 422340
rect 113180 422288 113232 422340
rect 113180 421540 113232 421592
rect 119436 421540 119488 421592
rect 120356 421540 120408 421592
rect 370504 418140 370556 418192
rect 580172 418140 580224 418192
rect 99380 406784 99432 406836
rect 100116 406784 100168 406836
rect 75920 406240 75972 406292
rect 76564 406240 76616 406292
rect 76564 405764 76616 405816
rect 173164 405764 173216 405816
rect 99380 405696 99432 405748
rect 342260 405696 342312 405748
rect 95884 405016 95936 405068
rect 128544 405016 128596 405068
rect 97908 404948 97960 405000
rect 132592 404948 132644 405000
rect 544384 404336 544436 404388
rect 580172 404336 580224 404388
rect 89812 403588 89864 403640
rect 113272 403588 113324 403640
rect 353300 403588 353352 403640
rect 74540 402976 74592 403028
rect 75184 402976 75236 403028
rect 153844 402976 153896 403028
rect 106188 402296 106240 402348
rect 117596 402296 117648 402348
rect 45284 402228 45336 402280
rect 85488 402228 85540 402280
rect 94044 402228 94096 402280
rect 120264 402228 120316 402280
rect 80796 401616 80848 401668
rect 327080 401616 327132 401668
rect 99196 401004 99248 401056
rect 131304 401004 131356 401056
rect 92664 400936 92716 400988
rect 111708 400936 111760 400988
rect 166264 400936 166316 400988
rect 98000 400868 98052 400920
rect 117504 400868 117556 400920
rect 351920 400868 351972 400920
rect 69204 400188 69256 400240
rect 226984 400188 227036 400240
rect 56416 399576 56468 399628
rect 84844 399576 84896 399628
rect 54944 399508 54996 399560
rect 85580 399508 85632 399560
rect 43904 399440 43956 399492
rect 87512 399440 87564 399492
rect 88248 399440 88300 399492
rect 95148 399440 95200 399492
rect 127348 399440 127400 399492
rect 88248 398896 88300 398948
rect 159364 398896 159416 398948
rect 72424 398828 72476 398880
rect 149244 398828 149296 398880
rect 204904 398828 204956 398880
rect 117228 398216 117280 398268
rect 125876 398216 125928 398268
rect 98552 398148 98604 398200
rect 127072 398148 127124 398200
rect 157984 398148 158036 398200
rect 53656 398080 53708 398132
rect 69296 398080 69348 398132
rect 88340 398080 88392 398132
rect 123300 398080 123352 398132
rect 162124 398080 162176 398132
rect 3424 397468 3476 397520
rect 50988 397468 51040 397520
rect 116584 397536 116636 397588
rect 117228 397536 117280 397588
rect 69296 397468 69348 397520
rect 268384 397468 268436 397520
rect 108856 396856 108908 396908
rect 117504 396856 117556 396908
rect 43812 396788 43864 396840
rect 71872 396788 71924 396840
rect 99288 396788 99340 396840
rect 131212 396788 131264 396840
rect 53472 396720 53524 396772
rect 83556 396720 83608 396772
rect 93768 396720 93820 396772
rect 127164 396720 127216 396772
rect 102140 396584 102192 396636
rect 102784 396584 102836 396636
rect 41144 396040 41196 396092
rect 102140 396040 102192 396092
rect 69112 395972 69164 396024
rect 69664 395972 69716 396024
rect 106924 395972 106976 396024
rect 134708 395972 134760 396024
rect 276020 395972 276072 396024
rect 276664 395972 276716 396024
rect 45284 395360 45336 395412
rect 78680 395360 78732 395412
rect 95976 395360 96028 395412
rect 127256 395428 127308 395480
rect 142344 395428 142396 395480
rect 48044 395292 48096 395344
rect 82820 395292 82872 395344
rect 96712 395292 96764 395344
rect 128452 395292 128504 395344
rect 150440 395360 150492 395412
rect 134708 395292 134760 395344
rect 276020 395292 276072 395344
rect 292488 395292 292540 395344
rect 385684 395292 385736 395344
rect 82820 394748 82872 394800
rect 83004 394748 83056 394800
rect 126336 394748 126388 394800
rect 69112 394680 69164 394732
rect 231860 394680 231912 394732
rect 68744 394612 68796 394664
rect 68928 394612 68980 394664
rect 53104 394068 53156 394120
rect 75368 394068 75420 394120
rect 52368 394000 52420 394052
rect 82912 394000 82964 394052
rect 101404 394000 101456 394052
rect 106280 394000 106332 394052
rect 108304 394000 108356 394052
rect 135444 394000 135496 394052
rect 49516 393932 49568 393984
rect 80704 393932 80756 393984
rect 95240 393932 95292 393984
rect 129004 393932 129056 393984
rect 82820 393456 82872 393508
rect 83096 393456 83148 393508
rect 138020 393456 138072 393508
rect 75368 393388 75420 393440
rect 134156 393388 134208 393440
rect 135444 393388 135496 393440
rect 316684 393388 316736 393440
rect 68928 393320 68980 393372
rect 278044 393320 278096 393372
rect 41236 393252 41288 393304
rect 82820 393252 82872 393304
rect 110880 392776 110932 392828
rect 125692 392776 125744 392828
rect 114284 392708 114336 392760
rect 139400 392708 139452 392760
rect 146944 392708 146996 392760
rect 57704 392640 57756 392692
rect 87604 392640 87656 392692
rect 104532 392640 104584 392692
rect 134064 392640 134116 392692
rect 36912 392572 36964 392624
rect 70400 392572 70452 392624
rect 94136 392572 94188 392624
rect 124404 392572 124456 392624
rect 152096 392572 152148 392624
rect 47860 392096 47912 392148
rect 110880 392096 110932 392148
rect 134064 392096 134116 392148
rect 136824 392096 136876 392148
rect 106280 392028 106332 392080
rect 360200 392028 360252 392080
rect 53564 391892 53616 391944
rect 57336 391892 57388 391944
rect 324320 391960 324372 392012
rect 91008 391892 91060 391944
rect 92572 391892 92624 391944
rect 47952 391280 48004 391332
rect 76012 391280 76064 391332
rect 103336 391280 103388 391332
rect 116124 391280 116176 391332
rect 55128 391212 55180 391264
rect 88984 391212 89036 391264
rect 102048 391212 102100 391264
rect 132684 391212 132736 391264
rect 133696 391212 133748 391264
rect 113916 390668 113968 390720
rect 167644 390668 167696 390720
rect 67548 390600 67600 390652
rect 136640 390600 136692 390652
rect 137284 390600 137336 390652
rect 140780 390600 140832 390652
rect 52276 390532 52328 390584
rect 79324 390532 79376 390584
rect 133696 390532 133748 390584
rect 313280 390532 313332 390584
rect 56508 390464 56560 390516
rect 67548 390464 67600 390516
rect 111064 390056 111116 390108
rect 114928 390056 114980 390108
rect 92572 389920 92624 389972
rect 121460 389920 121512 389972
rect 39948 389852 40000 389904
rect 69572 389852 69624 389904
rect 102600 389852 102652 389904
rect 135352 389852 135404 389904
rect 136548 389852 136600 389904
rect 38476 389784 38528 389836
rect 109040 389784 109092 389836
rect 119436 389784 119488 389836
rect 143816 389784 143868 389836
rect 115848 389444 115900 389496
rect 119436 389444 119488 389496
rect 69572 389376 69624 389428
rect 84476 389376 84528 389428
rect 120724 389376 120776 389428
rect 121644 389376 121696 389428
rect 54760 389308 54812 389360
rect 57888 389308 57940 389360
rect 80612 389308 80664 389360
rect 89720 389308 89772 389360
rect 90364 389308 90416 389360
rect 110328 389308 110380 389360
rect 137284 389308 137336 389360
rect 48964 389240 49016 389292
rect 120724 389240 120776 389292
rect 121460 389240 121512 389292
rect 122104 389240 122156 389292
rect 222844 389240 222896 389292
rect 56324 389172 56376 389224
rect 56508 389172 56560 389224
rect 63224 389172 63276 389224
rect 253204 389172 253256 389224
rect 102784 389104 102836 389156
rect 103612 389104 103664 389156
rect 104808 389104 104860 389156
rect 77300 388832 77352 388884
rect 77576 388832 77628 388884
rect 100024 388764 100076 388816
rect 101404 388764 101456 388816
rect 50804 388560 50856 388612
rect 54852 388560 54904 388612
rect 69756 388560 69808 388612
rect 58624 388492 58676 388544
rect 81440 388492 81492 388544
rect 48228 388424 48280 388476
rect 78220 388424 78272 388476
rect 95884 388220 95936 388272
rect 102140 388220 102192 388272
rect 104808 388220 104860 388272
rect 267004 388220 267056 388272
rect 109132 388152 109184 388204
rect 117964 388152 118016 388204
rect 94872 388084 94924 388136
rect 109040 388084 109092 388136
rect 112168 388084 112220 388136
rect 4804 388016 4856 388068
rect 72424 388016 72476 388068
rect 81440 388016 81492 388068
rect 82360 388016 82412 388068
rect 119436 388016 119488 388068
rect 143908 388016 143960 388068
rect 159456 388016 159508 388068
rect 53656 387948 53708 388000
rect 77576 387948 77628 388000
rect 93308 387948 93360 388000
rect 119528 387948 119580 388000
rect 39948 387880 40000 387932
rect 73344 387880 73396 387932
rect 108948 387880 109000 387932
rect 115756 387880 115808 387932
rect 117964 387880 118016 387932
rect 178684 387880 178736 387932
rect 70400 387812 70452 387864
rect 80060 387812 80112 387864
rect 91560 387812 91612 387864
rect 103520 387812 103572 387864
rect 104808 387812 104860 387864
rect 106188 387812 106240 387864
rect 111800 387812 111852 387864
rect 114928 387812 114980 387864
rect 184204 387812 184256 387864
rect 54852 387132 54904 387184
rect 83464 387132 83516 387184
rect 104808 387132 104860 387184
rect 118700 387132 118752 387184
rect 46664 387064 46716 387116
rect 78772 387064 78824 387116
rect 111156 387064 111208 387116
rect 130016 387064 130068 387116
rect 107568 386588 107620 386640
rect 126244 386588 126296 386640
rect 56508 386520 56560 386572
rect 87052 386520 87104 386572
rect 104440 386520 104492 386572
rect 104624 386520 104676 386572
rect 124404 386520 124456 386572
rect 34244 386452 34296 386504
rect 80520 386452 80572 386504
rect 118700 386452 118752 386504
rect 264244 386452 264296 386504
rect 78220 386384 78272 386436
rect 126980 386384 127032 386436
rect 301504 386384 301556 386436
rect 38568 386316 38620 386368
rect 58624 386316 58676 386368
rect 109040 386316 109092 386368
rect 125600 386316 125652 386368
rect 126888 386316 126940 386368
rect 45376 385840 45428 385892
rect 49608 385840 49660 385892
rect 49332 385704 49384 385756
rect 81532 385704 81584 385756
rect 126888 385704 126940 385756
rect 155224 385704 155276 385756
rect 52092 385636 52144 385688
rect 86316 385636 86368 385688
rect 91744 385636 91796 385688
rect 125692 385636 125744 385688
rect 35716 385092 35768 385144
rect 71780 385296 71832 385348
rect 49608 385024 49660 385076
rect 92940 385296 92992 385348
rect 101312 385296 101364 385348
rect 122288 385092 122340 385144
rect 123760 385092 123812 385144
rect 135904 385024 135956 385076
rect 60556 384276 60608 384328
rect 67640 384276 67692 384328
rect 118516 384276 118568 384328
rect 147588 384276 147640 384328
rect 118056 383664 118108 383716
rect 139400 383664 139452 383716
rect 119528 382916 119580 382968
rect 297364 382916 297416 382968
rect 126060 382304 126112 382356
rect 129924 382304 129976 382356
rect 39856 382236 39908 382288
rect 67640 382236 67692 382288
rect 118148 382236 118200 382288
rect 127624 382236 127676 382288
rect 118608 382168 118660 382220
rect 141056 382168 141108 382220
rect 141056 381556 141108 381608
rect 181444 381556 181496 381608
rect 118608 381488 118660 381540
rect 125600 381488 125652 381540
rect 126060 381488 126112 381540
rect 147588 381488 147640 381540
rect 349804 381488 349856 381540
rect 118608 380332 118660 380384
rect 122472 380332 122524 380384
rect 115296 380264 115348 380316
rect 117320 380264 117372 380316
rect 117688 380128 117740 380180
rect 118332 380128 118384 380180
rect 192484 380128 192536 380180
rect 65984 379652 66036 379704
rect 67732 379652 67784 379704
rect 60648 379584 60700 379636
rect 66168 379584 66220 379636
rect 67640 379584 67692 379636
rect 48044 379516 48096 379568
rect 69664 379516 69716 379568
rect 263600 379516 263652 379568
rect 264244 379516 264296 379568
rect 483664 379516 483716 379568
rect 35624 379448 35676 379500
rect 65616 379448 65668 379500
rect 65984 379448 66036 379500
rect 42616 379380 42668 379432
rect 69848 379380 69900 379432
rect 37188 378768 37240 378820
rect 69204 378768 69256 378820
rect 118608 378700 118660 378752
rect 124128 378700 124180 378752
rect 233884 378292 233936 378344
rect 357440 378292 357492 378344
rect 118056 378224 118108 378276
rect 244280 378224 244332 378276
rect 253204 378224 253256 378276
rect 347780 378224 347832 378276
rect 174544 378156 174596 378208
rect 323124 378156 323176 378208
rect 353944 378156 353996 378208
rect 580172 378156 580224 378208
rect 57888 378088 57940 378140
rect 61476 378088 61528 378140
rect 67640 378088 67692 378140
rect 244280 377408 244332 377460
rect 265256 377408 265308 377460
rect 267004 377408 267056 377460
rect 308404 377408 308456 377460
rect 249708 376796 249760 376848
rect 358820 376796 358872 376848
rect 117872 376728 117924 376780
rect 121460 376728 121512 376780
rect 197268 376728 197320 376780
rect 512000 376728 512052 376780
rect 52184 376660 52236 376712
rect 66904 376660 66956 376712
rect 67548 376660 67600 376712
rect 118608 376660 118660 376712
rect 146300 376660 146352 376712
rect 149060 376660 149112 376712
rect 119436 376048 119488 376100
rect 154580 376048 154632 376100
rect 120172 375980 120224 376032
rect 143724 375980 143776 376032
rect 319536 375980 319588 376032
rect 61384 375368 61436 375420
rect 64696 375368 64748 375420
rect 67640 375368 67692 375420
rect 118516 375368 118568 375420
rect 120172 375368 120224 375420
rect 265256 375368 265308 375420
rect 403624 375368 403676 375420
rect 61844 375300 61896 375352
rect 63408 375300 63460 375352
rect 118608 375300 118660 375352
rect 133880 375300 133932 375352
rect 135168 375300 135220 375352
rect 62028 374620 62080 374672
rect 65892 374620 65944 374672
rect 67640 374620 67692 374672
rect 121460 374620 121512 374672
rect 155960 374620 156012 374672
rect 140044 374280 140096 374332
rect 140688 374280 140740 374332
rect 224224 374212 224276 374264
rect 340880 374212 340932 374264
rect 155960 374144 156012 374196
rect 320088 374144 320140 374196
rect 63408 374008 63460 374060
rect 67640 374008 67692 374060
rect 140688 374008 140740 374060
rect 327172 374076 327224 374128
rect 204904 374008 204956 374060
rect 209780 374008 209832 374060
rect 471980 374008 472032 374060
rect 137376 373668 137428 373720
rect 138296 373668 138348 373720
rect 59268 373260 59320 373312
rect 67640 373260 67692 373312
rect 117320 373260 117372 373312
rect 185584 373260 185636 373312
rect 193956 372784 194008 372836
rect 282920 372784 282972 372836
rect 177396 372716 177448 372768
rect 333980 372716 334032 372768
rect 334624 372716 334676 372768
rect 123484 372648 123536 372700
rect 321744 372648 321796 372700
rect 118056 372580 118108 372632
rect 121460 372580 121512 372632
rect 138296 372580 138348 372632
rect 339500 372580 339552 372632
rect 3240 372512 3292 372564
rect 48964 372512 49016 372564
rect 61936 371832 61988 371884
rect 67640 371832 67692 371884
rect 142804 371832 142856 371884
rect 150624 371832 150676 371884
rect 212540 371832 212592 371884
rect 213828 371832 213880 371884
rect 276664 371424 276716 371476
rect 354680 371424 354732 371476
rect 200764 371356 200816 371408
rect 324504 371356 324556 371408
rect 213828 371288 213880 371340
rect 417424 371288 417476 371340
rect 117872 371220 117924 371272
rect 338764 371220 338816 371272
rect 41052 371152 41104 371204
rect 69296 371152 69348 371204
rect 118608 370540 118660 370592
rect 129832 370540 129884 370592
rect 121460 370472 121512 370524
rect 337384 370472 337436 370524
rect 177488 369996 177540 370048
rect 305092 369996 305144 370048
rect 118240 369928 118292 369980
rect 121460 369928 121512 369980
rect 162216 369928 162268 369980
rect 323216 369928 323268 369980
rect 166356 369860 166408 369912
rect 242164 369860 242216 369912
rect 244648 369860 244700 369912
rect 244924 369860 244976 369912
rect 517520 369860 517572 369912
rect 118608 369792 118660 369844
rect 122656 369792 122708 369844
rect 124312 369792 124364 369844
rect 66076 369452 66128 369504
rect 68376 369452 68428 369504
rect 121460 369112 121512 369164
rect 255320 369112 255372 369164
rect 119436 368772 119488 368824
rect 269856 368772 269908 368824
rect 352012 368772 352064 368824
rect 124956 368704 125008 368756
rect 312544 368704 312596 368756
rect 255320 368636 255372 368688
rect 464344 368636 464396 368688
rect 119344 368568 119396 368620
rect 335360 368568 335412 368620
rect 50344 368500 50396 368552
rect 55036 368500 55088 368552
rect 67640 368500 67692 368552
rect 223488 368500 223540 368552
rect 468484 368500 468536 368552
rect 127624 368432 127676 368484
rect 151820 368432 151872 368484
rect 197268 368432 197320 368484
rect 198004 368432 198056 368484
rect 118608 367888 118660 367940
rect 122840 367888 122892 367940
rect 209044 367344 209096 367396
rect 345020 367344 345072 367396
rect 180248 367276 180300 367328
rect 325792 367276 325844 367328
rect 222844 367208 222896 367260
rect 385684 367208 385736 367260
rect 160744 367140 160796 367192
rect 238208 367140 238260 367192
rect 297364 367140 297416 367192
rect 471244 367140 471296 367192
rect 123576 367072 123628 367124
rect 321652 367072 321704 367124
rect 56324 367004 56376 367056
rect 67640 367004 67692 367056
rect 118608 367004 118660 367056
rect 142160 367004 142212 367056
rect 146300 367004 146352 367056
rect 261852 366052 261904 366104
rect 320180 366052 320232 366104
rect 199384 365984 199436 366036
rect 227720 365984 227772 366036
rect 259368 365984 259420 366036
rect 349160 365984 349212 366036
rect 171784 365916 171836 365968
rect 295340 365916 295392 365968
rect 305000 365916 305052 365968
rect 350540 365916 350592 365968
rect 189724 365848 189776 365900
rect 331312 365848 331364 365900
rect 125048 365780 125100 365832
rect 293408 365780 293460 365832
rect 295340 365780 295392 365832
rect 295984 365780 296036 365832
rect 346400 365780 346452 365832
rect 148416 365712 148468 365764
rect 209044 365712 209096 365764
rect 216588 365712 216640 365764
rect 510620 365712 510672 365764
rect 60372 365644 60424 365696
rect 66076 365644 66128 365696
rect 117872 365644 117924 365696
rect 138204 365644 138256 365696
rect 117412 364964 117464 365016
rect 145012 364964 145064 365016
rect 163596 364760 163648 364812
rect 258264 364760 258316 364812
rect 259368 364760 259420 364812
rect 176016 364692 176068 364744
rect 224224 364692 224276 364744
rect 188436 364624 188488 364676
rect 303528 364624 303580 364676
rect 305092 364624 305144 364676
rect 305644 364624 305696 364676
rect 342352 364624 342404 364676
rect 123668 364556 123720 364608
rect 214840 364556 214892 364608
rect 343640 364556 343692 364608
rect 146944 364488 146996 364540
rect 324412 364488 324464 364540
rect 257344 364420 257396 364472
rect 447784 364420 447836 364472
rect 41236 364352 41288 364404
rect 69020 364352 69072 364404
rect 198648 364352 198700 364404
rect 118148 364284 118200 364336
rect 146392 364284 146444 364336
rect 508504 364284 508556 364336
rect 579804 364352 579856 364404
rect 579620 364284 579672 364336
rect 56324 363672 56376 363724
rect 69388 363672 69440 363724
rect 43996 363604 44048 363656
rect 67640 363604 67692 363656
rect 579620 363604 579672 363656
rect 195244 363264 195296 363316
rect 206468 363264 206520 363316
rect 187056 363196 187108 363248
rect 233884 363196 233936 363248
rect 242164 363196 242216 363248
rect 242532 363196 242584 363248
rect 323308 363196 323360 363248
rect 195336 363128 195388 363180
rect 285036 363128 285088 363180
rect 301504 363128 301556 363180
rect 413284 363128 413336 363180
rect 178868 363060 178920 363112
rect 236092 363060 236144 363112
rect 356060 363060 356112 363112
rect 196624 362992 196676 363044
rect 322112 362992 322164 363044
rect 164884 362924 164936 362976
rect 247040 362924 247092 362976
rect 118608 362856 118660 362908
rect 140964 362856 141016 362908
rect 268384 362924 268436 362976
rect 466460 362924 466512 362976
rect 305000 362856 305052 362908
rect 226984 362448 227036 362500
rect 229652 362448 229704 362500
rect 199568 362244 199620 362296
rect 223488 362244 223540 362296
rect 140964 362176 141016 362228
rect 180156 362176 180208 362228
rect 196716 362176 196768 362228
rect 249708 362176 249760 362228
rect 250904 362176 250956 362228
rect 313280 362176 313332 362228
rect 406384 362176 406436 362228
rect 310796 361972 310848 362024
rect 313280 361972 313332 362024
rect 258264 361904 258316 361956
rect 259920 361904 259972 361956
rect 274732 361904 274784 361956
rect 275928 361904 275980 361956
rect 514760 361904 514812 361956
rect 118608 361768 118660 361820
rect 120080 361768 120132 361820
rect 240600 361836 240652 361888
rect 289544 361836 289596 361888
rect 300768 361836 300820 361888
rect 193496 361768 193548 361820
rect 204536 361768 204588 361820
rect 221280 361768 221332 361820
rect 222844 361768 222896 361820
rect 224224 361768 224276 361820
rect 225788 361768 225840 361820
rect 278136 361768 278188 361820
rect 278596 361768 278648 361820
rect 320824 361768 320876 361820
rect 160836 361700 160888 361752
rect 202604 361700 202656 361752
rect 249708 361700 249760 361752
rect 316868 361700 316920 361752
rect 196808 361632 196860 361684
rect 276664 361632 276716 361684
rect 252468 361564 252520 361616
rect 281172 361632 281224 361684
rect 485044 361632 485096 361684
rect 303528 361564 303580 361616
rect 304356 361564 304408 361616
rect 37004 361496 37056 361548
rect 68008 361496 68060 361548
rect 130016 361496 130068 361548
rect 289544 361496 289596 361548
rect 45468 361428 45520 361480
rect 66996 361428 67048 361480
rect 67548 361428 67600 361480
rect 118056 361428 118108 361480
rect 147864 361428 147916 361480
rect 252468 361428 252520 361480
rect 146484 361360 146536 361412
rect 200764 361360 200816 361412
rect 119528 360952 119580 361004
rect 120264 360952 120316 361004
rect 64788 360816 64840 360868
rect 67640 360816 67692 360868
rect 198188 360884 198240 360936
rect 216588 360884 216640 360936
rect 217140 360884 217192 360936
rect 300768 360884 300820 360936
rect 452660 360884 452712 360936
rect 314660 360816 314712 360868
rect 312544 360408 312596 360460
rect 323032 360408 323084 360460
rect 285036 360340 285088 360392
rect 319444 360340 319496 360392
rect 145564 360272 145616 360324
rect 146484 360272 146536 360324
rect 308220 360272 308272 360324
rect 308404 360272 308456 360324
rect 359464 360272 359516 360324
rect 129096 360204 129148 360256
rect 130016 360204 130068 360256
rect 196900 360204 196952 360256
rect 257344 360204 257396 360256
rect 272156 360204 272208 360256
rect 389824 360204 389876 360256
rect 118516 360136 118568 360188
rect 149152 360136 149204 360188
rect 149704 360136 149756 360188
rect 118608 360068 118660 360120
rect 133788 360068 133840 360120
rect 39764 359456 39816 359508
rect 67640 359456 67692 359508
rect 68560 359456 68612 359508
rect 68928 359456 68980 359508
rect 133788 359456 133840 359508
rect 143724 359456 143776 359508
rect 317512 359456 317564 359508
rect 319628 359456 319680 359508
rect 193864 358912 193916 358964
rect 321560 358912 321612 358964
rect 169116 358844 169168 358896
rect 324596 358844 324648 358896
rect 158168 358776 158220 358828
rect 320364 358776 320416 358828
rect 64144 358708 64196 358760
rect 67456 358708 67508 358760
rect 67640 358708 67692 358760
rect 122656 358096 122708 358148
rect 146392 358096 146444 358148
rect 53564 358028 53616 358080
rect 67640 358028 67692 358080
rect 118608 358028 118660 358080
rect 120724 358028 120776 358080
rect 148324 358028 148376 358080
rect 193496 358028 193548 358080
rect 3424 357824 3476 357876
rect 7564 357824 7616 357876
rect 146392 357416 146444 357468
rect 198096 357416 198148 357468
rect 118608 357348 118660 357400
rect 144920 357348 144972 357400
rect 146208 357348 146260 357400
rect 198740 356940 198792 356992
rect 199660 356940 199712 356992
rect 118608 356668 118660 356720
rect 142436 356668 142488 356720
rect 142804 356668 142856 356720
rect 151084 356668 151136 356720
rect 193956 356668 194008 356720
rect 191104 356192 191156 356244
rect 197360 356192 197412 356244
rect 42616 356056 42668 356108
rect 67916 356056 67968 356108
rect 57796 355376 57848 355428
rect 67640 355376 67692 355428
rect 52184 355308 52236 355360
rect 54208 355308 54260 355360
rect 67732 355308 67784 355360
rect 118148 354696 118200 354748
rect 182824 354696 182876 354748
rect 117780 354628 117832 354680
rect 128636 354628 128688 354680
rect 128636 354016 128688 354068
rect 115940 353948 115992 354000
rect 137284 353948 137336 354000
rect 142160 353948 142212 354000
rect 198188 353948 198240 354000
rect 49608 352588 49660 352640
rect 68560 352588 68612 352640
rect 33048 352520 33100 352572
rect 63500 352520 63552 352572
rect 118608 352520 118660 352572
rect 144920 352452 144972 352504
rect 145564 352452 145616 352504
rect 15844 351908 15896 351960
rect 49424 351908 49476 351960
rect 49608 351908 49660 351960
rect 63500 351908 63552 351960
rect 64420 351908 64472 351960
rect 67640 351908 67692 351960
rect 118056 351840 118108 351892
rect 147772 351840 147824 351892
rect 118608 351160 118660 351212
rect 170404 351160 170456 351212
rect 177304 351160 177356 351212
rect 198740 351160 198792 351212
rect 322112 351160 322164 351212
rect 360844 351160 360896 351212
rect 504364 351160 504416 351212
rect 580172 351160 580224 351212
rect 60464 350548 60516 350600
rect 61844 350548 61896 350600
rect 67640 350548 67692 350600
rect 118608 350276 118660 350328
rect 124220 350276 124272 350328
rect 117964 349800 118016 349852
rect 118700 349800 118752 349852
rect 322756 349800 322808 349852
rect 323216 349800 323268 349852
rect 489184 349800 489236 349852
rect 46572 349188 46624 349240
rect 68008 349188 68060 349240
rect 35808 349120 35860 349172
rect 62120 349120 62172 349172
rect 67640 349052 67692 349104
rect 118608 349052 118660 349104
rect 151820 349052 151872 349104
rect 153108 349052 153160 349104
rect 117688 348984 117740 349036
rect 152004 348984 152056 349036
rect 153016 348984 153068 349036
rect 153108 348372 153160 348424
rect 188344 348372 188396 348424
rect 320824 348372 320876 348424
rect 448520 348372 448572 348424
rect 65524 347692 65576 347744
rect 66076 347692 66128 347744
rect 117412 347692 117464 347744
rect 132500 347692 132552 347744
rect 133788 347692 133840 347744
rect 133788 347012 133840 347064
rect 180064 347012 180116 347064
rect 319628 347012 319680 347064
rect 469220 347012 469272 347064
rect 66076 346944 66128 346996
rect 67640 346944 67692 346996
rect 183008 346400 183060 346452
rect 197360 346400 197412 346452
rect 7564 346332 7616 346384
rect 68560 346332 68612 346384
rect 68836 346332 68888 346384
rect 118608 346332 118660 346384
rect 142252 346332 142304 346384
rect 143448 346332 143500 346384
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 118516 345584 118568 345636
rect 119712 345584 119764 345636
rect 143632 345652 143684 345704
rect 144276 345652 144328 345704
rect 322480 345652 322532 345704
rect 327080 345652 327132 345704
rect 461584 345652 461636 345704
rect 43904 345040 43956 345092
rect 68652 345040 68704 345092
rect 118608 344972 118660 345024
rect 138112 344972 138164 345024
rect 46848 344292 46900 344344
rect 58992 344292 59044 344344
rect 138112 344292 138164 344344
rect 186964 344292 187016 344344
rect 321652 344292 321704 344344
rect 328460 344292 328512 344344
rect 58992 343680 59044 343732
rect 67640 343680 67692 343732
rect 41328 343612 41380 343664
rect 62764 343612 62816 343664
rect 67640 343544 67692 343596
rect 117872 343544 117924 343596
rect 150532 343544 150584 343596
rect 117504 342932 117556 342984
rect 126796 342932 126848 342984
rect 117688 342864 117740 342916
rect 127164 342864 127216 342916
rect 322480 342864 322532 342916
rect 327172 342864 327224 342916
rect 465080 342864 465132 342916
rect 34152 342184 34204 342236
rect 68652 342184 68704 342236
rect 118608 342184 118660 342236
rect 147680 342184 147732 342236
rect 328552 342184 328604 342236
rect 370504 342184 370556 342236
rect 147680 341504 147732 341556
rect 178776 341504 178828 341556
rect 322572 341504 322624 341556
rect 322848 341504 322900 341556
rect 328552 341504 328604 341556
rect 61752 340892 61804 340944
rect 63316 340892 63368 340944
rect 67640 340892 67692 340944
rect 117412 340824 117464 340876
rect 138296 340824 138348 340876
rect 117320 340756 117372 340808
rect 129096 340756 129148 340808
rect 43812 340212 43864 340264
rect 122748 340212 122800 340264
rect 150532 340212 150584 340264
rect 69204 340144 69256 340196
rect 132960 340144 133012 340196
rect 427820 340144 427872 340196
rect 497464 340144 497516 340196
rect 73068 339872 73120 339924
rect 73206 339872 73258 339924
rect 37096 339600 37148 339652
rect 70400 339600 70452 339652
rect 71320 339600 71372 339652
rect 59084 339532 59136 339584
rect 70492 339532 70544 339584
rect 70676 339532 70728 339584
rect 64512 339464 64564 339516
rect 67180 339464 67232 339516
rect 67640 339464 67692 339516
rect 106924 339464 106976 339516
rect 117320 339464 117372 339516
rect 132500 339464 132552 339516
rect 132960 339464 133012 339516
rect 169668 339464 169720 339516
rect 197360 339464 197412 339516
rect 322388 339464 322440 339516
rect 332876 339464 332928 339516
rect 113180 339396 113232 339448
rect 113916 339396 113968 339448
rect 119344 339396 119396 339448
rect 55864 339328 55916 339380
rect 73896 339328 73948 339380
rect 87420 339328 87472 339380
rect 87604 339328 87656 339380
rect 191104 339328 191156 339380
rect 54852 339260 54904 339312
rect 79692 339260 79744 339312
rect 104808 339260 104860 339312
rect 132684 339260 132736 339312
rect 97724 339124 97776 339176
rect 97908 339124 97960 339176
rect 117688 339124 117740 339176
rect 135260 339192 135312 339244
rect 84844 339056 84896 339108
rect 110604 338988 110656 339040
rect 111708 338988 111760 339040
rect 199568 339056 199620 339108
rect 68560 338852 68612 338904
rect 98644 338852 98696 338904
rect 55128 338784 55180 338836
rect 91008 338784 91060 338836
rect 91928 338784 91980 338836
rect 54852 338716 54904 338768
rect 104808 338716 104860 338768
rect 79692 338172 79744 338224
rect 83464 338172 83516 338224
rect 49516 338036 49568 338088
rect 53380 338036 53432 338088
rect 103520 338036 103572 338088
rect 131212 338036 131264 338088
rect 57704 337968 57756 338020
rect 91284 337968 91336 338020
rect 91744 337968 91796 338020
rect 115756 337968 115808 338020
rect 142252 337968 142304 338020
rect 143448 337968 143500 338020
rect 43720 337900 43772 337952
rect 74540 337900 74592 337952
rect 75276 337900 75328 337952
rect 115204 337900 115256 337952
rect 140044 337900 140096 337952
rect 50896 337832 50948 337884
rect 86132 337832 86184 337884
rect 86868 337832 86920 337884
rect 99656 337696 99708 337748
rect 100668 337696 100720 337748
rect 119528 337832 119580 337884
rect 109960 337764 110012 337816
rect 126336 337764 126388 337816
rect 115204 337696 115256 337748
rect 115388 337696 115440 337748
rect 45468 337492 45520 337544
rect 70032 337492 70084 337544
rect 101404 337492 101456 337544
rect 53380 337424 53432 337476
rect 82268 337424 82320 337476
rect 101956 337424 102008 337476
rect 102876 337424 102928 337476
rect 115112 337424 115164 337476
rect 150532 337424 150584 337476
rect 151728 337424 151780 337476
rect 197360 337424 197412 337476
rect 53748 337356 53800 337408
rect 55128 337356 55180 337408
rect 84200 337356 84252 337408
rect 86868 337356 86920 337408
rect 131212 337356 131264 337408
rect 133880 337356 133932 337408
rect 196900 337356 196952 337408
rect 107568 337288 107620 337340
rect 122196 337288 122248 337340
rect 91100 336812 91152 336864
rect 94504 336812 94556 336864
rect 126336 336812 126388 336864
rect 129740 336812 129792 336864
rect 75828 336744 75880 336796
rect 97264 336744 97316 336796
rect 49608 336676 49660 336728
rect 57244 336676 57296 336728
rect 91100 336676 91152 336728
rect 100300 336676 100352 336728
rect 129004 336744 129056 336796
rect 138112 336744 138164 336796
rect 143448 336744 143500 336796
rect 175924 336744 175976 336796
rect 54944 336608 54996 336660
rect 89076 336608 89128 336660
rect 106188 336608 106240 336660
rect 133972 336608 134024 336660
rect 56416 336540 56468 336592
rect 86408 336540 86460 336592
rect 113824 336540 113876 336592
rect 131120 336540 131172 336592
rect 48136 336472 48188 336524
rect 76564 336472 76616 336524
rect 46756 336404 46808 336456
rect 71964 336404 72016 336456
rect 72424 336404 72476 336456
rect 86224 336064 86276 336116
rect 117964 336064 118016 336116
rect 66996 335996 67048 336048
rect 121460 335996 121512 336048
rect 322480 335996 322532 336048
rect 333980 335996 334032 336048
rect 195428 335588 195480 335640
rect 197728 335588 197780 335640
rect 52092 335248 52144 335300
rect 88708 335248 88760 335300
rect 92572 335248 92624 335300
rect 93768 335248 93820 335300
rect 125692 335248 125744 335300
rect 46664 335180 46716 335232
rect 80704 335180 80756 335232
rect 98368 335180 98420 335232
rect 127348 335180 127400 335232
rect 42708 335112 42760 335164
rect 75920 335112 75972 335164
rect 108028 335112 108080 335164
rect 135444 335112 135496 335164
rect 52368 335044 52420 335096
rect 84844 335044 84896 335096
rect 97816 335044 97868 335096
rect 120264 335044 120316 335096
rect 121460 334568 121512 334620
rect 131212 334568 131264 334620
rect 188436 334568 188488 334620
rect 322480 334568 322532 334620
rect 325792 334568 325844 334620
rect 329840 334568 329892 334620
rect 97080 334500 97132 334552
rect 97816 334500 97868 334552
rect 75920 334364 75972 334416
rect 77116 334364 77168 334416
rect 50712 333956 50764 334008
rect 52368 333956 52420 334008
rect 88708 333956 88760 334008
rect 89168 333956 89220 334008
rect 127348 333956 127400 334008
rect 128360 333956 128412 334008
rect 45284 333888 45336 333940
rect 81624 333888 81676 333940
rect 95148 333888 95200 333940
rect 128544 333888 128596 333940
rect 189724 333888 189776 333940
rect 53472 333820 53524 333872
rect 87604 333820 87656 333872
rect 100944 333820 100996 333872
rect 102048 333820 102100 333872
rect 132592 333820 132644 333872
rect 49332 333752 49384 333804
rect 83556 333752 83608 333804
rect 189080 333208 189132 333260
rect 190368 333208 190420 333260
rect 199476 333208 199528 333260
rect 333980 333208 334032 333260
rect 371884 333208 371936 333260
rect 81624 332664 81676 332716
rect 82084 332664 82136 332716
rect 48136 332596 48188 332648
rect 53472 332596 53524 332648
rect 74632 332596 74684 332648
rect 189080 332596 189132 332648
rect 47952 332528 48004 332580
rect 78404 332528 78456 332580
rect 107384 332528 107436 332580
rect 125508 332528 125560 332580
rect 104900 331984 104952 332036
rect 127624 331984 127676 332036
rect 56416 331916 56468 331968
rect 124312 331916 124364 331968
rect 159548 331916 159600 331968
rect 37096 331848 37148 331900
rect 108028 331848 108080 331900
rect 122196 331848 122248 331900
rect 124404 331848 124456 331900
rect 175188 331848 175240 331900
rect 322204 331712 322256 331764
rect 327448 331712 327500 331764
rect 4804 331236 4856 331288
rect 37096 331236 37148 331288
rect 77944 331236 77996 331288
rect 78404 331236 78456 331288
rect 175188 331236 175240 331288
rect 197360 331236 197412 331288
rect 93216 331168 93268 331220
rect 122104 331168 122156 331220
rect 124312 331168 124364 331220
rect 322756 331032 322808 331084
rect 324320 331032 324372 331084
rect 52092 330556 52144 330608
rect 95056 330556 95108 330608
rect 95148 330556 95200 330608
rect 113824 330556 113876 330608
rect 57796 330488 57848 330540
rect 131120 330488 131172 330540
rect 160744 330488 160796 330540
rect 84292 329196 84344 329248
rect 116032 329196 116084 329248
rect 103520 329128 103572 329180
rect 151084 329128 151136 329180
rect 68744 329060 68796 329112
rect 177396 329060 177448 329112
rect 123760 328448 123812 328500
rect 124128 328448 124180 328500
rect 165528 328448 165580 328500
rect 197360 328448 197412 328500
rect 86316 327904 86368 327956
rect 124128 327904 124180 327956
rect 111800 327836 111852 327888
rect 174544 327836 174596 327888
rect 70492 327768 70544 327820
rect 141424 327768 141476 327820
rect 88340 327700 88392 327752
rect 178868 327700 178920 327752
rect 322756 327700 322808 327752
rect 324320 327700 324372 327752
rect 482284 327700 482336 327752
rect 107476 327088 107528 327140
rect 115296 327088 115348 327140
rect 185676 327088 185728 327140
rect 197360 327088 197412 327140
rect 108672 327020 108724 327072
rect 140872 327020 140924 327072
rect 93124 326544 93176 326596
rect 115388 326544 115440 326596
rect 54944 326476 54996 326528
rect 106924 326476 106976 326528
rect 115296 326476 115348 326528
rect 162216 326476 162268 326528
rect 57704 326408 57756 326460
rect 120172 326408 120224 326460
rect 140872 326408 140924 326460
rect 152648 326408 152700 326460
rect 88984 326340 89036 326392
rect 176016 326340 176068 326392
rect 322848 326340 322900 326392
rect 494152 326340 494204 326392
rect 106188 325048 106240 325100
rect 113824 325048 113876 325100
rect 71780 324980 71832 325032
rect 166356 324980 166408 325032
rect 96620 324912 96672 324964
rect 196808 324912 196860 324964
rect 360844 324912 360896 324964
rect 380900 324912 380952 324964
rect 320364 324300 320416 324352
rect 322848 324300 322900 324352
rect 380900 324300 380952 324352
rect 382188 324300 382240 324352
rect 580172 324300 580224 324352
rect 49424 323688 49476 323740
rect 117964 323688 118016 323740
rect 89168 323620 89220 323672
rect 160744 323620 160796 323672
rect 73160 323552 73212 323604
rect 164884 323552 164936 323604
rect 322480 322940 322532 322992
rect 331220 322940 331272 322992
rect 128268 322872 128320 322924
rect 134156 322872 134208 322924
rect 197360 322872 197412 322924
rect 70400 322192 70452 322244
rect 170496 322192 170548 322244
rect 77944 320900 77996 320952
rect 134524 320900 134576 320952
rect 49516 320832 49568 320884
rect 148416 320832 148468 320884
rect 167828 320832 167880 320884
rect 198188 320832 198240 320884
rect 172336 320152 172388 320204
rect 197360 320152 197412 320204
rect 322848 320152 322900 320204
rect 324320 320152 324372 320204
rect 499672 320152 499724 320204
rect 67456 319608 67508 319660
rect 122104 319608 122156 319660
rect 117320 319540 117372 319592
rect 180248 319540 180300 319592
rect 75184 319472 75236 319524
rect 108672 319472 108724 319524
rect 111064 319472 111116 319524
rect 177488 319472 177540 319524
rect 95332 319404 95384 319456
rect 171784 319404 171836 319456
rect 3424 319064 3476 319116
rect 7564 319064 7616 319116
rect 112536 318724 112588 318776
rect 143540 318724 143592 318776
rect 144828 318724 144880 318776
rect 84384 318112 84436 318164
rect 113916 318112 113968 318164
rect 65616 318044 65668 318096
rect 115204 318044 115256 318096
rect 144828 318044 144880 318096
rect 171784 318044 171836 318096
rect 115848 317500 115900 317552
rect 128636 317500 128688 317552
rect 155316 317500 155368 317552
rect 116676 317432 116728 317484
rect 193128 317432 193180 317484
rect 197360 317432 197412 317484
rect 101956 317364 102008 317416
rect 131304 317364 131356 317416
rect 131488 317364 131540 317416
rect 322480 317364 322532 317416
rect 335452 317364 335504 317416
rect 336648 317364 336700 317416
rect 93952 316820 94004 316872
rect 115848 316820 115900 316872
rect 131488 316820 131540 316872
rect 151084 316820 151136 316872
rect 69480 316752 69532 316804
rect 107108 316752 107160 316804
rect 111616 316752 111668 316804
rect 177488 316752 177540 316804
rect 80704 316684 80756 316736
rect 191104 316684 191156 316736
rect 336648 316684 336700 316736
rect 454684 316684 454736 316736
rect 75276 315936 75328 315988
rect 114652 315936 114704 315988
rect 114652 315324 114704 315376
rect 115296 315324 115348 315376
rect 79416 315256 79468 315308
rect 136824 315256 136876 315308
rect 166540 315256 166592 315308
rect 102784 314644 102836 314696
rect 184848 314644 184900 314696
rect 197360 314644 197412 314696
rect 7564 314576 7616 314628
rect 48044 314576 48096 314628
rect 105452 314576 105504 314628
rect 136732 314576 136784 314628
rect 322480 314576 322532 314628
rect 331312 314576 331364 314628
rect 82084 314032 82136 314084
rect 144184 314032 144236 314084
rect 90916 313964 90968 314016
rect 153936 313964 153988 314016
rect 48044 313896 48096 313948
rect 116584 313896 116636 313948
rect 136732 313896 136784 313948
rect 163504 313896 163556 313948
rect 331312 313896 331364 313948
rect 500960 313896 501012 313948
rect 129096 313284 129148 313336
rect 197360 313284 197412 313336
rect 60464 312672 60516 312724
rect 122196 312672 122248 312724
rect 97264 312604 97316 312656
rect 164884 312604 164936 312656
rect 81440 312536 81492 312588
rect 163596 312536 163648 312588
rect 181536 312536 181588 312588
rect 195428 312536 195480 312588
rect 322848 312536 322900 312588
rect 324504 312536 324556 312588
rect 395344 312536 395396 312588
rect 97816 311176 97868 311228
rect 156604 311176 156656 311228
rect 72424 311108 72476 311160
rect 148416 311108 148468 311160
rect 186320 311108 186372 311160
rect 187608 311108 187660 311160
rect 198096 311108 198148 311160
rect 89720 310564 89772 310616
rect 188988 310564 189040 310616
rect 197360 310564 197412 310616
rect 66168 310496 66220 310548
rect 186320 310496 186372 310548
rect 107108 310428 107160 310480
rect 125784 310428 125836 310480
rect 172336 310428 172388 310480
rect 173348 310428 173400 310480
rect 89076 309748 89128 309800
rect 152464 309748 152516 309800
rect 322480 309748 322532 309800
rect 325700 309748 325752 309800
rect 377404 309748 377456 309800
rect 178868 309204 178920 309256
rect 197360 309204 197412 309256
rect 73896 309136 73948 309188
rect 185676 309136 185728 309188
rect 126888 309068 126940 309120
rect 131304 309068 131356 309120
rect 96528 308524 96580 308576
rect 138664 308524 138716 308576
rect 73804 308456 73856 308508
rect 119896 308456 119948 308508
rect 83556 308388 83608 308440
rect 146944 308388 146996 308440
rect 165436 308388 165488 308440
rect 198280 308388 198332 308440
rect 73068 307096 73120 307148
rect 135996 307096 136048 307148
rect 85580 307028 85632 307080
rect 196716 307028 196768 307080
rect 321744 307028 321796 307080
rect 475384 307028 475436 307080
rect 70400 306484 70452 306536
rect 87604 306416 87656 306468
rect 162216 306416 162268 306468
rect 3424 306280 3476 306332
rect 15844 306280 15896 306332
rect 197452 306280 197504 306332
rect 199384 306280 199436 306332
rect 91008 305736 91060 305788
rect 136732 305736 136784 305788
rect 79324 305668 79376 305720
rect 142804 305668 142856 305720
rect 102048 305600 102100 305652
rect 166356 305600 166408 305652
rect 111156 304988 111208 305040
rect 167828 304988 167880 305040
rect 322480 304988 322532 305040
rect 327172 304988 327224 305040
rect 91744 304308 91796 304360
rect 149704 304308 149756 304360
rect 55036 304240 55088 304292
rect 134616 304240 134668 304292
rect 119896 303968 119948 304020
rect 123760 303968 123812 304020
rect 69204 303628 69256 303680
rect 197728 303628 197780 303680
rect 198648 303628 198700 303680
rect 99288 303016 99340 303068
rect 140044 303016 140096 303068
rect 66076 302948 66128 303000
rect 130568 302948 130620 303000
rect 79324 302880 79376 302932
rect 147036 302880 147088 302932
rect 186228 302880 186280 302932
rect 198004 302880 198056 302932
rect 113272 302336 113324 302388
rect 116676 302336 116728 302388
rect 48044 302268 48096 302320
rect 69112 302268 69164 302320
rect 69480 302268 69532 302320
rect 86960 302268 87012 302320
rect 163596 302268 163648 302320
rect 64512 302200 64564 302252
rect 193036 302200 193088 302252
rect 197360 302200 197412 302252
rect 322480 302200 322532 302252
rect 325700 302200 325752 302252
rect 58992 301656 59044 301708
rect 101404 301656 101456 301708
rect 93768 301588 93820 301640
rect 137284 301588 137336 301640
rect 87696 301520 87748 301572
rect 143816 301520 143868 301572
rect 162308 301520 162360 301572
rect 69480 301452 69532 301504
rect 184756 301452 184808 301504
rect 66904 301316 66956 301368
rect 68836 301316 68888 301368
rect 102140 300908 102192 300960
rect 133236 300908 133288 300960
rect 68836 300840 68888 300892
rect 162400 300840 162452 300892
rect 98552 300636 98604 300688
rect 102784 300636 102836 300688
rect 117872 300228 117924 300280
rect 125600 300228 125652 300280
rect 148508 300228 148560 300280
rect 104992 300160 105044 300212
rect 139400 300160 139452 300212
rect 170588 300160 170640 300212
rect 184756 300160 184808 300212
rect 197360 300160 197412 300212
rect 100760 300024 100812 300076
rect 101220 300024 101272 300076
rect 146392 300092 146444 300144
rect 176568 300092 176620 300144
rect 197268 300092 197320 300144
rect 322572 300092 322624 300144
rect 322756 300092 322808 300144
rect 356704 300092 356756 300144
rect 361488 300092 361540 300144
rect 580264 300092 580316 300144
rect 82820 299684 82872 299736
rect 136088 299684 136140 299736
rect 52368 299616 52420 299668
rect 100760 299616 100812 299668
rect 109684 299616 109736 299668
rect 115572 299616 115624 299668
rect 176568 299616 176620 299668
rect 81900 299548 81952 299600
rect 169024 299548 169076 299600
rect 11704 299480 11756 299532
rect 117872 299480 117924 299532
rect 94504 299072 94556 299124
rect 95148 299072 95200 299124
rect 111708 298800 111760 298852
rect 133144 298800 133196 298852
rect 83464 298732 83516 298784
rect 129740 298732 129792 298784
rect 94504 298324 94556 298376
rect 152740 298324 152792 298376
rect 99656 298256 99708 298308
rect 189724 298256 189776 298308
rect 53656 298052 53708 298104
rect 65524 298188 65576 298240
rect 167920 298188 167972 298240
rect 75276 298120 75328 298172
rect 182916 298120 182968 298172
rect 50804 297508 50856 297560
rect 56232 297508 56284 297560
rect 67548 297508 67600 297560
rect 25504 297372 25556 297424
rect 56324 297372 56376 297424
rect 97080 297372 97132 297424
rect 97908 297372 97960 297424
rect 145564 297372 145616 297424
rect 319536 297372 319588 297424
rect 353944 297372 353996 297424
rect 388444 297372 388496 297424
rect 194508 297236 194560 297288
rect 197360 297236 197412 297288
rect 112536 296964 112588 297016
rect 124864 296964 124916 297016
rect 100668 296896 100720 296948
rect 104808 296896 104860 296948
rect 116584 296896 116636 296948
rect 144276 296896 144328 296948
rect 83556 296828 83608 296880
rect 129004 296828 129056 296880
rect 90640 296760 90692 296812
rect 147036 296760 147088 296812
rect 76472 296692 76524 296744
rect 174636 296692 174688 296744
rect 59084 295944 59136 295996
rect 73896 295944 73948 295996
rect 149796 295944 149848 295996
rect 183008 295944 183060 295996
rect 107568 295672 107620 295724
rect 140136 295672 140188 295724
rect 100944 295604 100996 295656
rect 141516 295604 141568 295656
rect 113180 295536 113232 295588
rect 113824 295536 113876 295588
rect 158076 295536 158128 295588
rect 115204 295468 115256 295520
rect 115756 295468 115808 295520
rect 159640 295468 159692 295520
rect 68928 295400 68980 295452
rect 134800 295400 134852 295452
rect 69112 295332 69164 295384
rect 195704 295332 195756 295384
rect 197452 295332 197504 295384
rect 322480 295332 322532 295384
rect 331312 295332 331364 295384
rect 71320 295264 71372 295316
rect 75184 295264 75236 295316
rect 80336 295264 80388 295316
rect 86224 295264 86276 295316
rect 117044 295264 117096 295316
rect 123576 295264 123628 295316
rect 109316 294856 109368 294908
rect 111064 294856 111116 294908
rect 111248 294856 111300 294908
rect 124956 294856 125008 294908
rect 106740 294788 106792 294840
rect 125048 294788 125100 294840
rect 72608 294720 72660 294772
rect 87696 294720 87748 294772
rect 88708 294720 88760 294772
rect 119436 294720 119488 294772
rect 56508 294652 56560 294704
rect 111156 294652 111208 294704
rect 119620 294652 119672 294704
rect 149244 294652 149296 294704
rect 88064 294584 88116 294636
rect 107568 294584 107620 294636
rect 108028 294584 108080 294636
rect 196624 294584 196676 294636
rect 322756 294584 322808 294636
rect 420920 294584 420972 294636
rect 74632 294312 74684 294364
rect 75460 294312 75512 294364
rect 77300 294312 77352 294364
rect 78036 294312 78088 294364
rect 104900 294312 104952 294364
rect 105820 294312 105872 294364
rect 77116 294244 77168 294296
rect 79324 294244 79376 294296
rect 86132 294244 86184 294296
rect 87604 294244 87656 294296
rect 55036 294108 55088 294160
rect 74540 294108 74592 294160
rect 46756 294040 46808 294092
rect 79692 294040 79744 294092
rect 110604 294040 110656 294092
rect 117228 294040 117280 294092
rect 33784 293972 33836 294024
rect 79416 293972 79468 294024
rect 84200 293972 84252 294024
rect 180248 293972 180300 294024
rect 44088 293224 44140 293276
rect 75920 293224 75972 293276
rect 322848 293224 322900 293276
rect 324412 293224 324464 293276
rect 370504 293224 370556 293276
rect 2780 293156 2832 293208
rect 4804 293156 4856 293208
rect 93216 292884 93268 292936
rect 127624 292884 127676 292936
rect 53104 292816 53156 292868
rect 92572 292816 92624 292868
rect 92940 292816 92992 292868
rect 93860 292816 93912 292868
rect 130476 292816 130528 292868
rect 80980 292748 81032 292800
rect 123484 292748 123536 292800
rect 73896 292680 73948 292732
rect 124128 292680 124180 292732
rect 5448 292612 5500 292664
rect 96436 292612 96488 292664
rect 98368 292612 98420 292664
rect 98736 292612 98788 292664
rect 195336 292612 195388 292664
rect 68744 292544 68796 292596
rect 196624 292544 196676 292596
rect 71688 292476 71740 292528
rect 86408 292476 86460 292528
rect 121460 292476 121512 292528
rect 152096 292476 152148 292528
rect 155408 292476 155460 292528
rect 118056 292408 118108 292460
rect 124220 292408 124272 292460
rect 124128 292340 124180 292392
rect 129832 292340 129884 292392
rect 66076 291796 66128 291848
rect 89076 292068 89128 292120
rect 92296 291864 92348 291916
rect 117228 291864 117280 291916
rect 171876 291796 171928 291848
rect 156696 291184 156748 291236
rect 322480 291184 322532 291236
rect 340144 291184 340196 291236
rect 38568 291116 38620 291168
rect 67640 291116 67692 291168
rect 15844 290436 15896 290488
rect 38568 290436 38620 290488
rect 129280 290436 129332 290488
rect 142436 290436 142488 290488
rect 121552 289960 121604 290012
rect 152556 289960 152608 290012
rect 121460 289892 121512 289944
rect 173256 289892 173308 289944
rect 181628 289892 181680 289944
rect 197452 289892 197504 289944
rect 42708 289824 42760 289876
rect 67640 289824 67692 289876
rect 124036 289824 124088 289876
rect 198004 289824 198056 289876
rect 121552 289756 121604 289808
rect 195244 289756 195296 289808
rect 121460 289688 121512 289740
rect 123760 289688 123812 289740
rect 124036 289688 124088 289740
rect 69020 289144 69072 289196
rect 69756 289144 69808 289196
rect 123576 289076 123628 289128
rect 128360 289076 128412 289128
rect 187700 289076 187752 289128
rect 187700 288396 187752 288448
rect 188896 288396 188948 288448
rect 197452 288396 197504 288448
rect 340144 288396 340196 288448
rect 495440 288396 495492 288448
rect 121460 288328 121512 288380
rect 169116 288328 169168 288380
rect 121552 288260 121604 288312
rect 142344 288260 142396 288312
rect 143448 288260 143500 288312
rect 143448 287648 143500 287700
rect 163688 287648 163740 287700
rect 322756 287648 322808 287700
rect 358728 287648 358780 287700
rect 506480 287648 506532 287700
rect 49424 287036 49476 287088
rect 67640 287036 67692 287088
rect 52092 286968 52144 287020
rect 67732 286968 67784 287020
rect 121552 286968 121604 287020
rect 124220 286968 124272 287020
rect 121644 286900 121696 286952
rect 124312 286900 124364 286952
rect 121460 286832 121512 286884
rect 143724 286832 143776 286884
rect 66076 286288 66128 286340
rect 68192 286288 68244 286340
rect 143724 286288 143776 286340
rect 196808 286288 196860 286340
rect 52184 285676 52236 285728
rect 67824 285676 67876 285728
rect 191196 285676 191248 285728
rect 197452 285676 197504 285728
rect 322480 285676 322532 285728
rect 329932 285676 329984 285728
rect 58992 285608 59044 285660
rect 67640 285608 67692 285660
rect 121460 285608 121512 285660
rect 193864 285608 193916 285660
rect 121552 285540 121604 285592
rect 145012 285540 145064 285592
rect 121644 284996 121696 285048
rect 158168 284996 158220 285048
rect 145012 284928 145064 284980
rect 195980 284928 196032 284980
rect 38568 284316 38620 284368
rect 67640 284316 67692 284368
rect 65524 284248 65576 284300
rect 67732 284248 67784 284300
rect 121460 284248 121512 284300
rect 131304 284248 131356 284300
rect 126244 284180 126296 284232
rect 133604 284180 133656 284232
rect 121460 282888 121512 282940
rect 124956 282888 125008 282940
rect 132592 282888 132644 282940
rect 133604 282888 133656 282940
rect 190276 282888 190328 282940
rect 197452 282888 197504 282940
rect 322480 282888 322532 282940
rect 328552 282888 328604 282940
rect 41144 282820 41196 282872
rect 67640 282820 67692 282872
rect 121460 281528 121512 281580
rect 166448 281528 166500 281580
rect 180340 281528 180392 281580
rect 197452 281528 197504 281580
rect 121552 281460 121604 281512
rect 187056 281460 187108 281512
rect 178776 280780 178828 280832
rect 186136 280780 186188 280832
rect 50896 280168 50948 280220
rect 67640 280168 67692 280220
rect 121460 280168 121512 280220
rect 129188 280168 129240 280220
rect 186136 280168 186188 280220
rect 197452 280168 197504 280220
rect 322480 280168 322532 280220
rect 336004 280168 336056 280220
rect 41420 280100 41472 280152
rect 42616 280100 42668 280152
rect 67732 280100 67784 280152
rect 56232 280032 56284 280084
rect 67640 280032 67692 280084
rect 29644 279420 29696 279472
rect 41420 279420 41472 279472
rect 121460 278740 121512 278792
rect 192576 278740 192628 278792
rect 59084 278672 59136 278724
rect 67640 278672 67692 278724
rect 152648 277992 152700 278044
rect 183468 277992 183520 278044
rect 57796 277380 57848 277432
rect 67640 277380 67692 277432
rect 121460 277380 121512 277432
rect 142896 277380 142948 277432
rect 183468 277380 183520 277432
rect 197452 277380 197504 277432
rect 122748 277312 122800 277364
rect 160836 277312 160888 277364
rect 121460 277244 121512 277296
rect 132500 277244 132552 277296
rect 321836 276632 321888 276684
rect 493324 276632 493376 276684
rect 56140 276020 56192 276072
rect 67732 276020 67784 276072
rect 121460 276020 121512 276072
rect 160928 276020 160980 276072
rect 320824 276020 320876 276072
rect 321836 276020 321888 276072
rect 56508 275952 56560 276004
rect 67640 275952 67692 276004
rect 121552 274728 121604 274780
rect 122104 274728 122156 274780
rect 144368 274728 144420 274780
rect 175096 274728 175148 274780
rect 197452 274728 197504 274780
rect 53656 274660 53708 274712
rect 67640 274660 67692 274712
rect 121460 274660 121512 274712
rect 187056 274660 187108 274712
rect 60464 274592 60516 274644
rect 67732 274592 67784 274644
rect 322388 274592 322440 274644
rect 339500 274592 339552 274644
rect 133236 273912 133288 273964
rect 195244 273912 195296 273964
rect 339500 273912 339552 273964
rect 382924 273912 382976 273964
rect 121460 273300 121512 273352
rect 169116 273300 169168 273352
rect 43812 273232 43864 273284
rect 67640 273232 67692 273284
rect 123760 273232 123812 273284
rect 177948 273232 178000 273284
rect 197452 273232 197504 273284
rect 336004 273232 336056 273284
rect 457444 273232 457496 273284
rect 121460 273164 121512 273216
rect 133880 273164 133932 273216
rect 52092 271872 52144 271924
rect 67640 271872 67692 271924
rect 417424 271872 417476 271924
rect 419540 271872 419592 271924
rect 580172 271872 580224 271924
rect 53564 271804 53616 271856
rect 67732 271804 67784 271856
rect 124956 271124 125008 271176
rect 197452 271124 197504 271176
rect 65984 270512 66036 270564
rect 68100 270512 68152 270564
rect 121460 270512 121512 270564
rect 174544 270512 174596 270564
rect 121460 269628 121512 269680
rect 124956 269628 125008 269680
rect 176016 269288 176068 269340
rect 180340 269288 180392 269340
rect 59084 269084 59136 269136
rect 67640 269084 67692 269136
rect 121460 269084 121512 269136
rect 133236 269084 133288 269136
rect 322848 269084 322900 269136
rect 327264 269084 327316 269136
rect 47860 269016 47912 269068
rect 48228 269016 48280 269068
rect 121552 269016 121604 269068
rect 150440 269016 150492 269068
rect 43904 268404 43956 268456
rect 55220 268404 55272 268456
rect 48228 268336 48280 268388
rect 67640 268336 67692 268388
rect 134800 268336 134852 268388
rect 194324 268200 194376 268252
rect 197452 268200 197504 268252
rect 121460 267724 121512 267776
rect 134708 267724 134760 267776
rect 150440 267724 150492 267776
rect 154028 267724 154080 267776
rect 45376 267656 45428 267708
rect 67732 267656 67784 267708
rect 322480 267656 322532 267708
rect 335360 267656 335412 267708
rect 336648 267656 336700 267708
rect 55220 266976 55272 267028
rect 56324 266976 56376 267028
rect 67640 266976 67692 267028
rect 336648 266976 336700 267028
rect 499764 266976 499816 267028
rect 121460 266432 121512 266484
rect 144460 266432 144512 266484
rect 3056 266364 3108 266416
rect 50344 266364 50396 266416
rect 121552 266364 121604 266416
rect 158168 266364 158220 266416
rect 179420 266364 179472 266416
rect 180708 266364 180760 266416
rect 197360 266364 197412 266416
rect 54852 266296 54904 266348
rect 67640 266296 67692 266348
rect 121460 265004 121512 265056
rect 145656 265004 145708 265056
rect 121552 264936 121604 264988
rect 151360 264936 151412 264988
rect 322480 264936 322532 264988
rect 330024 264936 330076 264988
rect 121460 264868 121512 264920
rect 125600 264868 125652 264920
rect 21364 264188 21416 264240
rect 43996 264188 44048 264240
rect 53840 264188 53892 264240
rect 124128 264188 124180 264240
rect 183376 264188 183428 264240
rect 60464 263644 60516 263696
rect 67640 263644 67692 263696
rect 53840 263576 53892 263628
rect 54852 263576 54904 263628
rect 67732 263576 67784 263628
rect 121460 263576 121512 263628
rect 138756 263576 138808 263628
rect 175096 263576 175148 263628
rect 178776 263576 178828 263628
rect 183376 263576 183428 263628
rect 197360 263576 197412 263628
rect 360292 263576 360344 263628
rect 361488 263576 361540 263628
rect 490564 263576 490616 263628
rect 57704 263508 57756 263560
rect 67640 263508 67692 263560
rect 121552 263508 121604 263560
rect 121460 263440 121512 263492
rect 138112 263440 138164 263492
rect 138112 263032 138164 263084
rect 141608 263032 141660 263084
rect 334348 262828 334400 262880
rect 360292 262828 360344 262880
rect 60372 262216 60424 262268
rect 67640 262216 67692 262268
rect 64512 262148 64564 262200
rect 67824 262148 67876 262200
rect 121552 262148 121604 262200
rect 128268 262216 128320 262268
rect 152648 262216 152700 262268
rect 322480 262216 322532 262268
rect 334072 262216 334124 262268
rect 334348 262216 334400 262268
rect 121460 262012 121512 262064
rect 123760 262012 123812 262064
rect 123668 261468 123720 261520
rect 138020 261468 138072 261520
rect 186320 261468 186372 261520
rect 56508 260856 56560 260908
rect 67732 260856 67784 260908
rect 186320 260856 186372 260908
rect 187516 260856 187568 260908
rect 197360 260856 197412 260908
rect 56416 260788 56468 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 150440 260788 150492 260840
rect 150440 260108 150492 260160
rect 151728 260108 151780 260160
rect 160836 260108 160888 260160
rect 370504 260108 370556 260160
rect 520924 260108 520976 260160
rect 121460 259428 121512 259480
rect 131764 259428 131816 259480
rect 194416 259428 194468 259480
rect 197360 259428 197412 259480
rect 322480 259428 322532 259480
rect 327356 259428 327408 259480
rect 121552 259360 121604 259412
rect 136640 259360 136692 259412
rect 137100 259360 137152 259412
rect 137100 258680 137152 258732
rect 161020 258680 161072 258732
rect 188804 258680 188856 258732
rect 194416 258680 194468 258732
rect 520924 258680 520976 258732
rect 579988 258680 580040 258732
rect 66076 258136 66128 258188
rect 67640 258136 67692 258188
rect 322848 258136 322900 258188
rect 324504 258136 324556 258188
rect 57704 258068 57756 258120
rect 67732 258068 67784 258120
rect 121644 258068 121696 258120
rect 137468 258068 137520 258120
rect 393964 258068 394016 258120
rect 34244 258000 34296 258052
rect 67640 258000 67692 258052
rect 121460 258000 121512 258052
rect 154580 258000 154632 258052
rect 14464 257320 14516 257372
rect 34244 257320 34296 257372
rect 53564 256708 53616 256760
rect 67640 256708 67692 256760
rect 121552 256708 121604 256760
rect 126244 256708 126296 256760
rect 133880 256708 133932 256760
rect 197360 256708 197412 256760
rect 121460 256640 121512 256692
rect 136732 256640 136784 256692
rect 136732 256028 136784 256080
rect 169208 256028 169260 256080
rect 141608 255960 141660 256012
rect 181812 255960 181864 256012
rect 63132 255280 63184 255332
rect 67640 255280 67692 255332
rect 181812 255280 181864 255332
rect 182088 255280 182140 255332
rect 197360 255280 197412 255332
rect 50712 255212 50764 255264
rect 67732 255212 67784 255264
rect 52276 255144 52328 255196
rect 67640 255144 67692 255196
rect 122104 254600 122156 254652
rect 130384 254600 130436 254652
rect 122472 254532 122524 254584
rect 167736 254532 167788 254584
rect 121460 253920 121512 253972
rect 142988 253920 143040 253972
rect 47676 253852 47728 253904
rect 48044 253852 48096 253904
rect 67640 253852 67692 253904
rect 63224 253784 63276 253836
rect 67732 253784 67784 253836
rect 32404 253172 32456 253224
rect 47676 253172 47728 253224
rect 121460 252628 121512 252680
rect 155500 252628 155552 252680
rect 120816 252560 120868 252612
rect 191748 252560 191800 252612
rect 197360 252560 197412 252612
rect 322848 252560 322900 252612
rect 324412 252560 324464 252612
rect 121460 252492 121512 252544
rect 155960 252492 156012 252544
rect 192852 251608 192904 251660
rect 196716 251608 196768 251660
rect 121460 251200 121512 251252
rect 184296 251200 184348 251252
rect 66168 251132 66220 251184
rect 67640 251132 67692 251184
rect 167920 250452 167972 250504
rect 194416 250452 194468 250504
rect 194416 249908 194468 249960
rect 197360 249908 197412 249960
rect 121460 249772 121512 249824
rect 133328 249772 133380 249824
rect 121552 249704 121604 249756
rect 140228 249772 140280 249824
rect 156788 249772 156840 249824
rect 121460 249636 121512 249688
rect 129096 249636 129148 249688
rect 35716 249024 35768 249076
rect 56232 249024 56284 249076
rect 195336 248956 195388 249008
rect 197360 248956 197412 249008
rect 56232 248412 56284 248464
rect 67640 248412 67692 248464
rect 322480 248412 322532 248464
rect 335452 248412 335504 248464
rect 434720 248412 434772 248464
rect 121460 247120 121512 247172
rect 137376 247120 137428 247172
rect 66168 247052 66220 247104
rect 67640 247052 67692 247104
rect 121552 247052 121604 247104
rect 178960 247052 179012 247104
rect 135904 246508 135956 246560
rect 136640 246508 136692 246560
rect 121460 246168 121512 246220
rect 125048 246168 125100 246220
rect 121552 245692 121604 245744
rect 151268 245692 151320 245744
rect 136640 245624 136692 245676
rect 195888 245624 195940 245676
rect 198096 245624 198148 245676
rect 322480 245624 322532 245676
rect 332692 245624 332744 245676
rect 374644 245624 374696 245676
rect 54944 245556 54996 245608
rect 67640 245556 67692 245608
rect 53380 245488 53432 245540
rect 67364 245488 67416 245540
rect 195336 245012 195388 245064
rect 196716 245012 196768 245064
rect 137468 244876 137520 244928
rect 189816 244876 189868 244928
rect 121552 244264 121604 244316
rect 123760 244264 123812 244316
rect 321744 244264 321796 244316
rect 378784 244264 378836 244316
rect 37096 244196 37148 244248
rect 67732 244196 67784 244248
rect 121460 244196 121512 244248
rect 131212 244196 131264 244248
rect 49516 244128 49568 244180
rect 67640 244128 67692 244180
rect 194232 243788 194284 243840
rect 195980 243788 196032 243840
rect 198280 243788 198332 243840
rect 194324 243652 194376 243704
rect 195980 243652 196032 243704
rect 68560 243516 68612 243568
rect 68928 243516 68980 243568
rect 145656 243516 145708 243568
rect 195336 243516 195388 243568
rect 135168 242972 135220 243024
rect 176108 242972 176160 243024
rect 121552 242904 121604 242956
rect 191656 242904 191708 242956
rect 321468 242904 321520 242956
rect 443644 242904 443696 242956
rect 121460 242836 121512 242888
rect 134616 242836 134668 242888
rect 135168 242836 135220 242888
rect 155500 242156 155552 242208
rect 193864 242156 193916 242208
rect 121460 241476 121512 241528
rect 140688 241476 140740 241528
rect 3424 241408 3476 241460
rect 40868 241408 40920 241460
rect 41236 241408 41288 241460
rect 322204 241408 322256 241460
rect 324596 241408 324648 241460
rect 162400 240796 162452 240848
rect 195796 240796 195848 240848
rect 40868 240728 40920 240780
rect 58716 240728 58768 240780
rect 144460 240728 144512 240780
rect 196532 240728 196584 240780
rect 121460 240252 121512 240304
rect 155500 240252 155552 240304
rect 120632 240184 120684 240236
rect 191196 240184 191248 240236
rect 119988 240116 120040 240168
rect 199660 240116 199712 240168
rect 324596 240116 324648 240168
rect 502340 240116 502392 240168
rect 3516 240048 3568 240100
rect 37188 240048 37240 240100
rect 194508 240048 194560 240100
rect 196808 240048 196860 240100
rect 70400 239776 70452 239828
rect 71308 239776 71360 239828
rect 76012 239776 76064 239828
rect 77104 239776 77156 239828
rect 84292 239776 84344 239828
rect 85476 239776 85528 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 89720 239776 89772 239828
rect 90628 239776 90680 239828
rect 95240 239776 95292 239828
rect 96424 239776 96476 239828
rect 102140 239776 102192 239828
rect 102864 239776 102916 239828
rect 107660 239776 107712 239828
rect 108660 239776 108712 239828
rect 110420 239776 110472 239828
rect 111236 239776 111288 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 219440 239776 219492 239828
rect 220590 239776 220642 239828
rect 238760 239776 238812 239828
rect 239910 239776 239962 239828
rect 247040 239776 247092 239828
rect 248282 239776 248334 239828
rect 258080 239776 258132 239828
rect 259230 239776 259282 239828
rect 266360 239776 266412 239828
rect 267602 239776 267654 239828
rect 285680 239776 285732 239828
rect 286922 239776 286974 239828
rect 63132 239572 63184 239624
rect 73804 239572 73856 239624
rect 60372 239504 60424 239556
rect 76380 239504 76432 239556
rect 65984 239436 66036 239488
rect 195060 239436 195112 239488
rect 204168 239436 204220 239488
rect 319536 239436 319588 239488
rect 69848 239368 69900 239420
rect 83464 239368 83516 239420
rect 191656 239368 191708 239420
rect 320088 239368 320140 239420
rect 321744 239368 321796 239420
rect 535460 239368 535512 239420
rect 580172 239368 580224 239420
rect 200948 239164 201000 239216
rect 204904 239164 204956 239216
rect 199844 239096 199896 239148
rect 202236 239096 202288 239148
rect 77760 239028 77812 239080
rect 200120 239028 200172 239080
rect 104164 238960 104216 239012
rect 120816 238960 120868 239012
rect 121460 238960 121512 239012
rect 155592 238960 155644 239012
rect 195980 238960 196032 239012
rect 202144 238960 202196 239012
rect 85580 238892 85632 238944
rect 86776 238892 86828 238944
rect 123576 238892 123628 238944
rect 37188 238824 37240 238876
rect 111892 238824 111944 238876
rect 112536 238824 112588 238876
rect 114468 238824 114520 238876
rect 124404 238824 124456 238876
rect 152740 238824 152792 238876
rect 237380 238824 237432 238876
rect 238024 238824 238076 238876
rect 201592 238756 201644 238808
rect 252836 238756 252888 238808
rect 535460 238756 535512 238808
rect 50988 238688 51040 238740
rect 82268 238688 82320 238740
rect 118976 238688 119028 238740
rect 130568 238688 130620 238740
rect 48136 238620 48188 238672
rect 72608 238620 72660 238672
rect 83556 238620 83608 238672
rect 149060 238620 149112 238672
rect 316592 238620 316644 238672
rect 88708 238552 88760 238604
rect 241888 238552 241940 238604
rect 118332 238484 118384 238536
rect 144920 238484 144972 238536
rect 195336 238484 195388 238536
rect 331588 238484 331640 238536
rect 115112 238416 115164 238468
rect 146300 238416 146352 238468
rect 200120 238416 200172 238468
rect 216772 238416 216824 238468
rect 105452 238348 105504 238400
rect 282184 238348 282236 238400
rect 69940 238280 69992 238332
rect 119988 238280 120040 238332
rect 71964 238144 72016 238196
rect 79232 238144 79284 238196
rect 80980 238144 81032 238196
rect 88984 238144 89036 238196
rect 73252 238076 73304 238128
rect 86224 238076 86276 238128
rect 196624 238076 196676 238128
rect 204076 238076 204128 238128
rect 315948 238076 316000 238128
rect 320180 238076 320232 238128
rect 67548 238008 67600 238060
rect 105544 238008 105596 238060
rect 184296 238008 184348 238060
rect 200672 238008 200724 238060
rect 316592 238008 316644 238060
rect 438860 238008 438912 238060
rect 204076 237668 204128 237720
rect 205824 237668 205876 237720
rect 244280 237464 244332 237516
rect 246396 237464 246448 237516
rect 216772 237396 216824 237448
rect 217324 237396 217376 237448
rect 221464 237396 221516 237448
rect 223212 237396 223264 237448
rect 229744 237396 229796 237448
rect 231584 237396 231636 237448
rect 235356 237396 235408 237448
rect 236092 237396 236144 237448
rect 246304 237396 246356 237448
rect 250904 237396 250956 237448
rect 251824 237396 251876 237448
rect 254768 237396 254820 237448
rect 291844 237396 291896 237448
rect 297272 237396 297324 237448
rect 300124 237396 300176 237448
rect 301780 237396 301832 237448
rect 307116 237396 307168 237448
rect 308220 237396 308272 237448
rect 312636 237396 312688 237448
rect 314016 237396 314068 237448
rect 318064 237396 318116 237448
rect 318524 237396 318576 237448
rect 498292 237396 498344 237448
rect 58716 237328 58768 237380
rect 103520 237328 103572 237380
rect 113180 237328 113232 237380
rect 114468 237328 114520 237380
rect 149796 237328 149848 237380
rect 198004 237328 198056 237380
rect 204168 237328 204220 237380
rect 55128 237260 55180 237312
rect 86132 237260 86184 237312
rect 95792 237260 95844 237312
rect 126980 237260 127032 237312
rect 142896 237260 142948 237312
rect 331312 237260 331364 237312
rect 49608 237192 49660 237244
rect 76656 237192 76708 237244
rect 113824 237192 113876 237244
rect 133880 237192 133932 237244
rect 151360 237192 151412 237244
rect 328552 237192 328604 237244
rect 195888 237124 195940 237176
rect 303712 237124 303764 237176
rect 148600 237056 148652 237108
rect 195980 237056 196032 237108
rect 183376 236988 183428 237040
rect 504364 236988 504416 237040
rect 160928 236716 160980 236768
rect 195336 236716 195388 236768
rect 68652 236648 68704 236700
rect 249800 236648 249852 236700
rect 316684 235968 316736 236020
rect 320272 235968 320324 236020
rect 503720 235968 503772 236020
rect 504364 235968 504416 236020
rect 89352 235900 89404 235952
rect 142160 235900 142212 235952
rect 158168 235900 158220 235952
rect 329932 235900 329984 235952
rect 91284 235832 91336 235884
rect 129280 235832 129332 235884
rect 174636 235832 174688 235884
rect 244280 235832 244332 235884
rect 244924 235832 244976 235884
rect 73896 235764 73948 235816
rect 120632 235764 120684 235816
rect 39764 235696 39816 235748
rect 91744 235696 91796 235748
rect 118608 235696 118660 235748
rect 131120 235696 131172 235748
rect 194232 235492 194284 235544
rect 213184 235492 213236 235544
rect 163596 235424 163648 235476
rect 196624 235424 196676 235476
rect 187056 235356 187108 235408
rect 222844 235356 222896 235408
rect 106096 235288 106148 235340
rect 175096 235288 175148 235340
rect 198832 235288 198884 235340
rect 324688 235288 324740 235340
rect 67364 235220 67416 235272
rect 280252 235220 280304 235272
rect 303712 235220 303764 235272
rect 498384 235220 498436 235272
rect 175096 235084 175148 235136
rect 176016 235084 176068 235136
rect 117688 234948 117740 235000
rect 118608 234948 118660 235000
rect 288900 234608 288952 234660
rect 289452 234608 289504 234660
rect 432604 234608 432656 234660
rect 46572 234540 46624 234592
rect 109040 234540 109092 234592
rect 134708 234540 134760 234592
rect 327264 234540 327316 234592
rect 328368 234540 328420 234592
rect 48228 234472 48280 234524
rect 195152 234472 195204 234524
rect 196532 234472 196584 234524
rect 321468 234472 321520 234524
rect 322204 234472 322256 234524
rect 50344 234404 50396 234456
rect 85580 234404 85632 234456
rect 200672 234404 200724 234456
rect 321560 234404 321612 234456
rect 321836 234404 321888 234456
rect 159640 234336 159692 234388
rect 218704 234336 218756 234388
rect 109040 234132 109092 234184
rect 109960 234132 110012 234184
rect 47584 234064 47636 234116
rect 48228 234064 48280 234116
rect 74540 233860 74592 233912
rect 75184 233860 75236 233912
rect 79232 233860 79284 233912
rect 84292 233928 84344 233980
rect 84200 233724 84252 233776
rect 171876 233928 171928 233980
rect 270500 233928 270552 233980
rect 328368 233928 328420 233980
rect 335360 233928 335412 233980
rect 202788 233860 202840 233912
rect 203892 233860 203944 233912
rect 321560 233860 321612 233912
rect 333980 233860 334032 233912
rect 60464 233180 60516 233232
rect 327080 233180 327132 233232
rect 328368 233180 328420 233232
rect 56508 233112 56560 233164
rect 178868 233112 178920 233164
rect 81624 233044 81676 233096
rect 132592 233044 132644 233096
rect 156788 233044 156840 233096
rect 265624 233044 265676 233096
rect 166540 232976 166592 233028
rect 262956 232976 263008 233028
rect 189816 232568 189868 232620
rect 222936 232568 222988 232620
rect 328368 232568 328420 232620
rect 345112 232568 345164 232620
rect 169668 232500 169720 232552
rect 418160 232500 418212 232552
rect 418160 231820 418212 231872
rect 419448 231820 419500 231872
rect 580172 231820 580224 231872
rect 54852 231752 54904 231804
rect 319260 231752 319312 231804
rect 82820 231684 82872 231736
rect 136640 231684 136692 231736
rect 144368 231684 144420 231736
rect 334072 231684 334124 231736
rect 87052 231616 87104 231668
rect 235356 231616 235408 231668
rect 147128 231548 147180 231600
rect 292580 231548 292632 231600
rect 193036 231140 193088 231192
rect 209136 231140 209188 231192
rect 182088 231072 182140 231124
rect 496820 231072 496872 231124
rect 292580 230936 292632 230988
rect 293224 230936 293276 230988
rect 38568 230392 38620 230444
rect 327356 230392 327408 230444
rect 328368 230392 328420 230444
rect 76656 230324 76708 230376
rect 280160 230324 280212 230376
rect 281448 230324 281500 230376
rect 73804 230256 73856 230308
rect 187700 230256 187752 230308
rect 195336 230256 195388 230308
rect 325700 230256 325752 230308
rect 100208 229848 100260 229900
rect 249064 229848 249116 229900
rect 255964 229848 256016 229900
rect 315948 229848 316000 229900
rect 328368 229848 328420 229900
rect 336740 229848 336792 229900
rect 111892 229780 111944 229832
rect 262864 229780 262916 229832
rect 281448 229780 281500 229832
rect 340236 229780 340288 229832
rect 17224 229712 17276 229764
rect 83556 229712 83608 229764
rect 187700 229712 187752 229764
rect 188804 229712 188856 229764
rect 350632 229712 350684 229764
rect 315948 229100 316000 229152
rect 316776 229100 316828 229152
rect 56324 229032 56376 229084
rect 318064 229032 318116 229084
rect 155592 228964 155644 229016
rect 311900 228964 311952 229016
rect 97632 228896 97684 228948
rect 251824 228896 251876 228948
rect 162308 228828 162360 228880
rect 277400 228828 277452 228880
rect 59084 228352 59136 228404
rect 145656 228352 145708 228404
rect 190276 228352 190328 228404
rect 521660 228352 521712 228404
rect 277400 227740 277452 227792
rect 278044 227740 278096 227792
rect 311900 227740 311952 227792
rect 312544 227740 312596 227792
rect 91744 227672 91796 227724
rect 298744 227672 298796 227724
rect 178960 227604 179012 227656
rect 340144 227604 340196 227656
rect 84384 227536 84436 227588
rect 229744 227536 229796 227588
rect 95056 227468 95108 227520
rect 181536 227468 181588 227520
rect 187608 227060 187660 227112
rect 307024 227060 307076 227112
rect 52092 226992 52144 227044
rect 245016 226992 245068 227044
rect 305644 226992 305696 227044
rect 342904 226992 342956 227044
rect 202696 226312 202748 226364
rect 318064 226312 318116 226364
rect 123760 226244 123812 226296
rect 309140 226244 309192 226296
rect 56232 226176 56284 226228
rect 233240 226176 233292 226228
rect 193864 226108 193916 226160
rect 330024 226108 330076 226160
rect 70492 226040 70544 226092
rect 201500 226040 201552 226092
rect 202696 226040 202748 226092
rect 185676 225700 185728 225752
rect 211804 225700 211856 225752
rect 42708 225632 42760 225684
rect 266452 225632 266504 225684
rect 210240 225564 210292 225616
rect 485136 225564 485188 225616
rect 233240 224952 233292 225004
rect 233884 224952 233936 225004
rect 309140 224952 309192 225004
rect 309876 224952 309928 225004
rect 95240 224884 95292 224936
rect 260840 224884 260892 224936
rect 261484 224884 261536 224936
rect 76012 224816 76064 224868
rect 213920 224816 213972 224868
rect 222936 224816 222988 224868
rect 321652 224816 321704 224868
rect 159548 224748 159600 224800
rect 289820 224748 289872 224800
rect 290464 224748 290516 224800
rect 154028 224680 154080 224732
rect 276020 224680 276072 224732
rect 276664 224680 276716 224732
rect 213920 224408 213972 224460
rect 214564 224408 214616 224460
rect 66076 224272 66128 224324
rect 220084 224272 220136 224324
rect 67456 224204 67508 224256
rect 251180 224204 251232 224256
rect 276664 224204 276716 224256
rect 478880 224204 478932 224256
rect 247040 223592 247092 223644
rect 318156 223592 318208 223644
rect 102232 223524 102284 223576
rect 273260 223524 273312 223576
rect 273996 223524 274048 223576
rect 93952 223456 94004 223508
rect 247040 223456 247092 223508
rect 170588 223388 170640 223440
rect 238760 223388 238812 223440
rect 239496 223388 239548 223440
rect 68744 222912 68796 222964
rect 253940 222912 253992 222964
rect 183468 222844 183520 222896
rect 475476 222844 475528 222896
rect 195980 222164 196032 222216
rect 196808 222164 196860 222216
rect 347872 222164 347924 222216
rect 69204 222096 69256 222148
rect 256700 222096 256752 222148
rect 163688 222028 163740 222080
rect 300124 222028 300176 222080
rect 74632 221960 74684 222012
rect 195980 221960 196032 222012
rect 256700 221960 256752 222012
rect 257344 221960 257396 222012
rect 195244 221552 195296 221604
rect 278780 221552 278832 221604
rect 49424 221484 49476 221536
rect 232596 221484 232648 221536
rect 175188 221416 175240 221468
rect 510712 221416 510764 221468
rect 142988 220736 143040 220788
rect 323584 220804 323636 220856
rect 347964 220804 348016 220856
rect 158076 220668 158128 220720
rect 332692 220668 332744 220720
rect 177488 220260 177540 220312
rect 232504 220260 232556 220312
rect 101496 220192 101548 220244
rect 255320 220192 255372 220244
rect 57704 220124 57756 220176
rect 277400 220124 277452 220176
rect 181628 220056 181680 220108
rect 417424 220056 417476 220108
rect 148508 219376 148560 219428
rect 335452 219376 335504 219428
rect 84292 219308 84344 219360
rect 229100 219308 229152 219360
rect 230388 219308 230440 219360
rect 86224 219240 86276 219292
rect 208400 219240 208452 219292
rect 475384 218900 475436 218952
rect 480260 218900 480312 218952
rect 230388 218832 230440 218884
rect 291936 218832 291988 218884
rect 156696 218764 156748 218816
rect 238024 218764 238076 218816
rect 140136 218696 140188 218748
rect 258172 218696 258224 218748
rect 483664 218696 483716 218748
rect 514852 218696 514904 218748
rect 208400 218016 208452 218068
rect 209228 218016 209280 218068
rect 220728 218016 220780 218068
rect 346492 218016 346544 218068
rect 514852 218016 514904 218068
rect 580172 218016 580224 218068
rect 110512 217948 110564 218000
rect 140780 217948 140832 218000
rect 336004 217948 336056 218000
rect 78772 217880 78824 217932
rect 219440 217880 219492 217932
rect 220728 217880 220780 217932
rect 198924 217404 198976 217456
rect 324504 217404 324556 217456
rect 130476 217336 130528 217388
rect 263600 217336 263652 217388
rect 170496 217268 170548 217320
rect 367100 217268 367152 217320
rect 53564 216588 53616 216640
rect 312636 216588 312688 216640
rect 92572 216520 92624 216572
rect 246304 216520 246356 216572
rect 152556 216044 152608 216096
rect 240784 216044 240836 216096
rect 145656 215976 145708 216028
rect 274732 215976 274784 216028
rect 184756 215908 184808 215960
rect 446496 215908 446548 215960
rect 3332 215228 3384 215280
rect 21364 215228 21416 215280
rect 118700 215228 118752 215280
rect 307116 215228 307168 215280
rect 186136 214820 186188 214872
rect 240876 214820 240928 214872
rect 93860 214752 93912 214804
rect 246396 214752 246448 214804
rect 53656 214684 53708 214736
rect 235264 214684 235316 214736
rect 233884 214616 233936 214668
rect 486424 214616 486476 214668
rect 176568 214548 176620 214600
rect 502984 214548 503036 214600
rect 72424 213868 72476 213920
rect 258080 213868 258132 213920
rect 259368 213868 259420 213920
rect 103704 213800 103756 213852
rect 271880 213800 271932 213852
rect 272524 213800 272576 213852
rect 80060 213732 80112 213784
rect 221464 213732 221516 213784
rect 182916 213324 182968 213376
rect 267740 213324 267792 213376
rect 127624 213256 127676 213308
rect 236644 213256 236696 213308
rect 187516 213188 187568 213240
rect 407764 213188 407816 213240
rect 114560 212440 114612 212492
rect 295340 212440 295392 212492
rect 88984 212372 89036 212424
rect 224960 212372 225012 212424
rect 225604 212372 225656 212424
rect 295340 212032 295392 212084
rect 295984 212032 296036 212084
rect 153844 211964 153896 212016
rect 286324 211964 286376 212016
rect 102140 211896 102192 211948
rect 249984 211896 250036 211948
rect 259368 211896 259420 211948
rect 341524 211896 341576 211948
rect 126428 211828 126480 211880
rect 277492 211828 277544 211880
rect 173348 211760 173400 211812
rect 507860 211760 507912 211812
rect 107752 211080 107804 211132
rect 285680 211080 285732 211132
rect 319536 211148 319588 211200
rect 432604 211080 432656 211132
rect 446404 211080 446456 211132
rect 431960 210672 432012 210724
rect 432604 210672 432656 210724
rect 136088 210536 136140 210588
rect 262220 210536 262272 210588
rect 43812 210468 43864 210520
rect 239404 210468 239456 210520
rect 7564 210400 7616 210452
rect 110512 210400 110564 210452
rect 167644 210400 167696 210452
rect 231124 210400 231176 210452
rect 237380 210400 237432 210452
rect 483020 210400 483072 210452
rect 422300 209992 422352 210044
rect 425704 209992 425756 210044
rect 105544 209720 105596 209772
rect 266360 209720 266412 209772
rect 162216 209176 162268 209228
rect 226984 209176 227036 209228
rect 159456 209108 159508 209160
rect 273904 209108 273956 209160
rect 56140 209040 56192 209092
rect 222936 209040 222988 209092
rect 239496 209040 239548 209092
rect 513288 209040 513340 209092
rect 266360 208360 266412 208412
rect 267004 208360 267056 208412
rect 99380 208292 99432 208344
rect 269120 208292 269172 208344
rect 196624 207816 196676 207868
rect 280160 207816 280212 207868
rect 77300 207748 77352 207800
rect 252836 207748 252888 207800
rect 272524 207748 272576 207800
rect 325700 207748 325752 207800
rect 46756 207680 46808 207732
rect 276020 207680 276072 207732
rect 194416 207612 194468 207664
rect 517612 207612 517664 207664
rect 269120 207000 269172 207052
rect 269764 207000 269816 207052
rect 149704 206456 149756 206508
rect 196624 206456 196676 206508
rect 122196 206388 122248 206440
rect 252744 206388 252796 206440
rect 74540 206320 74592 206372
rect 254032 206320 254084 206372
rect 262956 206320 263008 206372
rect 505192 206320 505244 206372
rect 180708 206252 180760 206304
rect 436100 206252 436152 206304
rect 512644 206252 512696 206304
rect 513288 206252 513340 206304
rect 580172 206252 580224 206304
rect 107660 205572 107712 205624
rect 284300 205572 284352 205624
rect 140044 205096 140096 205148
rect 195244 205096 195296 205148
rect 284300 205096 284352 205148
rect 284944 205096 284996 205148
rect 89812 205028 89864 205080
rect 228364 205028 228416 205080
rect 76564 204960 76616 205012
rect 263692 204960 263744 205012
rect 188896 204892 188948 204944
rect 400864 204892 400916 204944
rect 98000 204212 98052 204264
rect 147680 204212 147732 204264
rect 148324 204212 148376 204264
rect 429844 204212 429896 204264
rect 431224 204212 431276 204264
rect 147036 203736 147088 203788
rect 233884 203736 233936 203788
rect 96620 203668 96672 203720
rect 259460 203668 259512 203720
rect 111800 203600 111852 203652
rect 276112 203600 276164 203652
rect 293224 203600 293276 203652
rect 429844 203600 429896 203652
rect 147680 203532 147732 203584
rect 399484 203532 399536 203584
rect 3424 202784 3476 202836
rect 120172 202784 120224 202836
rect 198556 202376 198608 202428
rect 321560 202376 321612 202428
rect 115940 202308 115992 202360
rect 245108 202308 245160 202360
rect 137284 202240 137336 202292
rect 349252 202240 349304 202292
rect 55036 202172 55088 202224
rect 269120 202172 269172 202224
rect 144276 202104 144328 202156
rect 396724 202104 396776 202156
rect 157984 201016 158036 201068
rect 213276 201016 213328 201068
rect 211804 200948 211856 201000
rect 313924 200948 313976 201000
rect 191748 200880 191800 200932
rect 296076 200880 296128 200932
rect 141516 200812 141568 200864
rect 273260 200812 273312 200864
rect 166264 200744 166316 200796
rect 199476 200744 199528 200796
rect 204904 200744 204956 200796
rect 513380 200744 513432 200796
rect 155500 199588 155552 199640
rect 238116 199588 238168 199640
rect 133144 199520 133196 199572
rect 216036 199520 216088 199572
rect 177948 199452 178000 199504
rect 338120 199452 338172 199504
rect 86960 199384 87012 199436
rect 267832 199384 267884 199436
rect 300124 199384 300176 199436
rect 509332 199384 509384 199436
rect 144184 198092 144236 198144
rect 289176 198092 289228 198144
rect 83464 198024 83516 198076
rect 232688 198024 232740 198076
rect 172428 197956 172480 198008
rect 200764 197956 200816 198008
rect 218704 197956 218756 198008
rect 516140 197956 516192 198008
rect 189724 196800 189776 196852
rect 281540 196800 281592 196852
rect 151084 196732 151136 196784
rect 291844 196732 291896 196784
rect 295984 196732 296036 196784
rect 327172 196732 327224 196784
rect 138664 196664 138716 196716
rect 351184 196664 351236 196716
rect 124956 196596 125008 196648
rect 265164 196596 265216 196648
rect 278044 196596 278096 196648
rect 506572 196596 506624 196648
rect 235356 195440 235408 195492
rect 309784 195440 309836 195492
rect 178868 195372 178920 195424
rect 314016 195372 314068 195424
rect 89720 195304 89772 195356
rect 254124 195304 254176 195356
rect 257344 195304 257396 195356
rect 325976 195304 326028 195356
rect 145564 195236 145616 195288
rect 199384 195236 199436 195288
rect 213184 195236 213236 195288
rect 503812 195236 503864 195288
rect 217324 194080 217376 194132
rect 321652 194080 321704 194132
rect 126244 194012 126296 194064
rect 240968 194012 241020 194064
rect 100760 193944 100812 193996
rect 252652 193944 252704 193996
rect 142804 193876 142856 193928
rect 354772 193876 354824 193928
rect 152648 193808 152700 193860
rect 410616 193808 410668 193860
rect 151268 192788 151320 192840
rect 242256 192788 242308 192840
rect 141424 192720 141476 192772
rect 211804 192720 211856 192772
rect 225604 192720 225656 192772
rect 328736 192720 328788 192772
rect 92480 192652 92532 192704
rect 256976 192652 257028 192704
rect 175096 192584 175148 192636
rect 343824 192584 343876 192636
rect 70400 192516 70452 192568
rect 254216 192516 254268 192568
rect 165528 192448 165580 192500
rect 411904 192448 411956 192500
rect 249064 191292 249116 191344
rect 271880 191292 271932 191344
rect 202236 191224 202288 191276
rect 335544 191224 335596 191276
rect 69112 191156 69164 191208
rect 251272 191156 251324 191208
rect 273996 191156 274048 191208
rect 331404 191156 331456 191208
rect 118608 191088 118660 191140
rect 503904 191088 503956 191140
rect 153936 190068 153988 190120
rect 195336 190068 195388 190120
rect 192576 190000 192628 190052
rect 243544 190000 243596 190052
rect 169024 189932 169076 189984
rect 264980 189932 265032 189984
rect 135996 189864 136048 189916
rect 198004 189864 198056 189916
rect 221464 189864 221516 189916
rect 335636 189864 335688 189916
rect 138756 189796 138808 189848
rect 256792 189796 256844 189848
rect 181536 189728 181588 189780
rect 345204 189728 345256 189780
rect 3424 188980 3476 189032
rect 53104 188980 53156 189032
rect 155224 188572 155276 188624
rect 204996 188572 205048 188624
rect 220084 188572 220136 188624
rect 273352 188572 273404 188624
rect 124864 188504 124916 188556
rect 271972 188504 272024 188556
rect 84200 188436 84252 188488
rect 250076 188436 250128 188488
rect 114468 188368 114520 188420
rect 334072 188368 334124 188420
rect 57796 188300 57848 188352
rect 259552 188300 259604 188352
rect 265624 188300 265676 188352
rect 494336 188300 494388 188352
rect 137376 187144 137428 187196
rect 255412 187144 255464 187196
rect 110420 187076 110472 187128
rect 249892 187076 249944 187128
rect 146944 187008 146996 187060
rect 352104 187008 352156 187060
rect 50896 186940 50948 186992
rect 266360 186940 266412 186992
rect 228364 185920 228416 185972
rect 262404 185920 262456 185972
rect 134524 185852 134576 185904
rect 213184 185852 213236 185904
rect 229744 185852 229796 185904
rect 342444 185852 342496 185904
rect 122104 185784 122156 185836
rect 249064 185784 249116 185836
rect 131764 185716 131816 185768
rect 263784 185716 263836 185768
rect 191196 185648 191248 185700
rect 339592 185648 339644 185700
rect 393964 185648 394016 185700
rect 425336 185648 425388 185700
rect 125048 185580 125100 185632
rect 258356 185580 258408 185632
rect 290464 185580 290516 185632
rect 498476 185580 498528 185632
rect 102048 184900 102100 184952
rect 205088 184900 205140 184952
rect 244924 184356 244976 184408
rect 290464 184356 290516 184408
rect 485044 184356 485096 184408
rect 501144 184356 501196 184408
rect 173256 184288 173308 184340
rect 251364 184288 251416 184340
rect 251824 184288 251876 184340
rect 340972 184288 341024 184340
rect 471244 184288 471296 184340
rect 488632 184288 488684 184340
rect 152464 184220 152516 184272
rect 202236 184220 202288 184272
rect 214564 184220 214616 184272
rect 330116 184220 330168 184272
rect 457444 184220 457496 184272
rect 510804 184220 510856 184272
rect 160836 184152 160888 184204
rect 506664 184152 506716 184204
rect 107568 183608 107620 183660
rect 173164 183608 173216 183660
rect 125508 183540 125560 183592
rect 214656 183540 214708 183592
rect 169116 183132 169168 183184
rect 260932 183132 260984 183184
rect 160744 183064 160796 183116
rect 215944 183064 215996 183116
rect 242164 183064 242216 183116
rect 341064 183064 341116 183116
rect 133328 182996 133380 183048
rect 248052 182996 248104 183048
rect 202788 182928 202840 182980
rect 352196 182928 352248 182980
rect 184848 182860 184900 182912
rect 345296 182860 345348 182912
rect 414664 182860 414716 182912
rect 505100 182860 505152 182912
rect 22744 182792 22796 182844
rect 109040 182792 109092 182844
rect 178776 182792 178828 182844
rect 343916 182792 343968 182844
rect 419264 182792 419316 182844
rect 580264 182792 580316 182844
rect 132408 182384 132460 182436
rect 164884 182384 164936 182436
rect 110696 182316 110748 182368
rect 170496 182316 170548 182368
rect 112444 182248 112496 182300
rect 171968 182248 172020 182300
rect 119528 182180 119580 182232
rect 196808 182180 196860 182232
rect 489184 182180 489236 182232
rect 490564 182180 490616 182232
rect 454684 182112 454736 182164
rect 455604 182112 455656 182164
rect 461584 182112 461636 182164
rect 462596 182112 462648 182164
rect 475476 182112 475528 182164
rect 476580 182112 476632 182164
rect 485136 182112 485188 182164
rect 485780 182112 485832 182164
rect 242256 181704 242308 181756
rect 260840 181704 260892 181756
rect 486424 181704 486476 181756
rect 492864 181704 492916 181756
rect 240968 181636 241020 181688
rect 262312 181636 262364 181688
rect 410524 181636 410576 181688
rect 444012 181636 444064 181688
rect 446496 181636 446548 181688
rect 460204 181636 460256 181688
rect 464344 181636 464396 181688
rect 474188 181636 474240 181688
rect 482284 181636 482336 181688
rect 502524 181636 502576 181688
rect 159364 181568 159416 181620
rect 198096 181568 198148 181620
rect 222844 181568 222896 181620
rect 269212 181568 269264 181620
rect 284944 181568 284996 181620
rect 338212 181568 338264 181620
rect 403624 181568 403676 181620
rect 441620 181568 441672 181620
rect 443644 181568 443696 181620
rect 505284 181568 505336 181620
rect 166356 181500 166408 181552
rect 209044 181500 209096 181552
rect 232688 181500 232740 181552
rect 259644 181500 259696 181552
rect 262864 181500 262916 181552
rect 446404 181500 446456 181552
rect 447784 181500 447836 181552
rect 507952 181500 508004 181552
rect 196716 181432 196768 181484
rect 451372 181432 451424 181484
rect 468484 181432 468536 181484
rect 501236 181432 501288 181484
rect 129464 180956 129516 181008
rect 166540 180956 166592 181008
rect 124036 180888 124088 180940
rect 167920 180888 167972 180940
rect 118424 180820 118476 180872
rect 169208 180820 169260 180872
rect 238116 180344 238168 180396
rect 261024 180344 261076 180396
rect 222936 180276 222988 180328
rect 249340 180276 249392 180328
rect 165436 180208 165488 180260
rect 239036 180208 239088 180260
rect 309876 180208 309928 180260
rect 325884 180208 325936 180260
rect 167828 180140 167880 180192
rect 335452 180140 335504 180192
rect 493324 180140 493376 180192
rect 512092 180140 512144 180192
rect 156604 180072 156656 180124
rect 210424 180072 210476 180124
rect 216128 180072 216180 180124
rect 509240 180072 509292 180124
rect 385684 180004 385736 180056
rect 386328 180004 386380 180056
rect 490656 179868 490708 179920
rect 495532 179868 495584 179920
rect 134708 179596 134760 179648
rect 165436 179596 165488 179648
rect 126612 179528 126664 179580
rect 170680 179528 170732 179580
rect 115848 179460 115900 179512
rect 166264 179460 166316 179512
rect 414664 179460 414716 179512
rect 492588 179460 492640 179512
rect 97816 179392 97868 179444
rect 171876 179392 171928 179444
rect 386328 179392 386380 179444
rect 580264 179392 580316 179444
rect 236644 178984 236696 179036
rect 255504 178984 255556 179036
rect 240784 178916 240836 178968
rect 265072 178916 265124 178968
rect 231124 178848 231176 178900
rect 274640 178848 274692 178900
rect 312544 178848 312596 178900
rect 327264 178848 327316 178900
rect 180248 178780 180300 178832
rect 247960 178780 248012 178832
rect 261484 178780 261536 178832
rect 321284 178780 321336 178832
rect 246304 178712 246356 178764
rect 349344 178712 349396 178764
rect 195888 178644 195940 178696
rect 417516 178644 417568 178696
rect 502984 178644 503036 178696
rect 580172 178644 580224 178696
rect 98736 178372 98788 178424
rect 196716 178372 196768 178424
rect 148232 178304 148284 178356
rect 170404 178304 170456 178356
rect 110328 178236 110380 178288
rect 178776 178236 178828 178288
rect 113732 178168 113784 178220
rect 196900 178168 196952 178220
rect 127072 178100 127124 178152
rect 214564 178100 214616 178152
rect 159916 178032 159968 178084
rect 169024 178032 169076 178084
rect 308404 178032 308456 178084
rect 316040 178032 316092 178084
rect 316408 178032 316460 178084
rect 246396 177624 246448 177676
rect 255596 177624 255648 177676
rect 314016 177624 314068 177676
rect 332784 177624 332836 177676
rect 238024 177556 238076 177608
rect 258264 177556 258316 177608
rect 312636 177556 312688 177608
rect 339500 177556 339552 177608
rect 174544 177488 174596 177540
rect 258080 177488 258132 177540
rect 307116 177488 307168 177540
rect 334164 177488 334216 177540
rect 239036 177420 239088 177472
rect 334256 177420 334308 177472
rect 209136 177352 209188 177404
rect 332600 177352 332652 177404
rect 198648 177284 198700 177336
rect 323124 177284 323176 177336
rect 133144 177012 133196 177064
rect 165528 177012 165580 177064
rect 108120 176944 108172 176996
rect 169116 176944 169168 176996
rect 103336 176876 103388 176928
rect 167552 176876 167604 176928
rect 136088 176808 136140 176860
rect 202788 176808 202840 176860
rect 104624 176740 104676 176792
rect 174636 176740 174688 176792
rect 128176 176672 128228 176724
rect 214196 176672 214248 176724
rect 340144 176672 340196 176724
rect 416780 176672 416832 176724
rect 202788 176604 202840 176656
rect 213920 176604 213972 176656
rect 243544 176604 243596 176656
rect 249248 176604 249300 176656
rect 319536 176604 319588 176656
rect 327080 176604 327132 176656
rect 163504 176264 163556 176316
rect 206376 176264 206428 176316
rect 120816 176196 120868 176248
rect 166632 176196 166684 176248
rect 121920 176128 121972 176180
rect 173256 176128 173308 176180
rect 102048 176060 102100 176112
rect 167828 176060 167880 176112
rect 318156 176060 318208 176112
rect 328644 176060 328696 176112
rect 130752 175992 130804 176044
rect 214104 175992 214156 176044
rect 245108 175992 245160 176044
rect 261116 175992 261168 176044
rect 318064 175992 318116 176044
rect 331496 175992 331548 176044
rect 116952 175924 117004 175976
rect 166356 175924 166408 175976
rect 166448 175924 166500 175976
rect 251456 175924 251508 175976
rect 269764 175924 269816 175976
rect 324412 175924 324464 175976
rect 495532 175924 495584 175976
rect 502432 175924 502484 175976
rect 248052 175788 248104 175840
rect 249156 175788 249208 175840
rect 165436 175176 165488 175228
rect 213920 175176 213972 175228
rect 165528 175108 165580 175160
rect 214012 175108 214064 175160
rect 338764 174496 338816 174548
rect 348424 174496 348476 174548
rect 296260 174020 296312 174072
rect 307668 174020 307720 174072
rect 285220 173952 285272 174004
rect 307576 173952 307628 174004
rect 265808 173884 265860 173936
rect 307116 173884 307168 173936
rect 358084 173884 358136 173936
rect 416780 173884 416832 173936
rect 164884 173816 164936 173868
rect 213920 173816 213972 173868
rect 252468 173816 252520 173868
rect 263600 173816 263652 173868
rect 280804 172660 280856 172712
rect 307576 172660 307628 172712
rect 263048 172592 263100 172644
rect 307116 172592 307168 172644
rect 260380 172524 260432 172576
rect 307668 172524 307720 172576
rect 496912 172524 496964 172576
rect 501052 172524 501104 172576
rect 166540 172456 166592 172508
rect 213920 172456 213972 172508
rect 252468 172456 252520 172508
rect 260932 172456 260984 172508
rect 324320 172456 324372 172508
rect 358820 172456 358872 172508
rect 252100 172388 252152 172440
rect 255412 172388 255464 172440
rect 261668 171776 261720 171828
rect 307300 171776 307352 171828
rect 252468 171504 252520 171556
rect 258080 171504 258132 171556
rect 167644 171300 167696 171352
rect 170588 171300 170640 171352
rect 283656 171164 283708 171216
rect 306932 171164 306984 171216
rect 267188 171096 267240 171148
rect 307668 171096 307720 171148
rect 170680 171028 170732 171080
rect 213920 171028 213972 171080
rect 324320 171028 324372 171080
rect 354680 171028 354732 171080
rect 252376 170552 252428 170604
rect 256884 170552 256936 170604
rect 252468 170144 252520 170196
rect 259644 170144 259696 170196
rect 285128 169872 285180 169924
rect 307300 169872 307352 169924
rect 268476 169804 268528 169856
rect 307668 169804 307720 169856
rect 260288 169736 260340 169788
rect 307484 169736 307536 169788
rect 324964 169736 325016 169788
rect 327080 169736 327132 169788
rect 167920 169668 167972 169720
rect 213920 169668 213972 169720
rect 324320 169668 324372 169720
rect 335636 169668 335688 169720
rect 324504 169600 324556 169652
rect 332600 169600 332652 169652
rect 252376 169464 252428 169516
rect 258172 169464 258224 169516
rect 252468 169124 252520 169176
rect 259460 169124 259512 169176
rect 174636 168988 174688 169040
rect 214472 168988 214524 169040
rect 297364 168988 297416 169040
rect 306564 168988 306616 169040
rect 264428 168444 264480 168496
rect 307116 168444 307168 168496
rect 264244 168376 264296 168428
rect 307668 168376 307720 168428
rect 338764 168376 338816 168428
rect 416780 168376 416832 168428
rect 166632 168308 166684 168360
rect 214012 168308 214064 168360
rect 252468 168308 252520 168360
rect 262220 168308 262272 168360
rect 324320 168308 324372 168360
rect 347780 168308 347832 168360
rect 496912 168308 496964 168360
rect 502340 168308 502392 168360
rect 503628 168308 503680 168360
rect 173256 168240 173308 168292
rect 213920 168240 213972 168292
rect 324504 168240 324556 168292
rect 345020 168240 345072 168292
rect 300216 167696 300268 167748
rect 306748 167696 306800 167748
rect 259368 167628 259420 167680
rect 307024 167628 307076 167680
rect 503628 167628 503680 167680
rect 543004 167628 543056 167680
rect 252468 167560 252520 167612
rect 258264 167560 258316 167612
rect 269856 167016 269908 167068
rect 307484 167016 307536 167068
rect 166356 166948 166408 167000
rect 214104 166948 214156 167000
rect 252376 166948 252428 167000
rect 263692 166948 263744 167000
rect 324320 166948 324372 167000
rect 334256 166948 334308 167000
rect 496912 166948 496964 167000
rect 503904 166948 503956 167000
rect 504180 166948 504232 167000
rect 169208 166880 169260 166932
rect 214012 166880 214064 166932
rect 252468 166880 252520 166932
rect 261024 166880 261076 166932
rect 196808 166812 196860 166864
rect 213920 166812 213972 166864
rect 252284 166812 252336 166864
rect 256976 166812 257028 166864
rect 287796 166268 287848 166320
rect 307300 166268 307352 166320
rect 504180 166268 504232 166320
rect 555424 166268 555476 166320
rect 271328 165656 271380 165708
rect 307668 165656 307720 165708
rect 257436 165588 257488 165640
rect 306748 165588 306800 165640
rect 353944 165588 353996 165640
rect 416780 165588 416832 165640
rect 556160 165588 556212 165640
rect 580172 165588 580224 165640
rect 166264 165520 166316 165572
rect 213920 165520 213972 165572
rect 252468 165520 252520 165572
rect 270500 165520 270552 165572
rect 324320 165520 324372 165572
rect 335544 165520 335596 165572
rect 497004 165520 497056 165572
rect 509332 165520 509384 165572
rect 510528 165520 510580 165572
rect 252284 165452 252336 165504
rect 262404 165452 262456 165504
rect 324504 165452 324556 165504
rect 331404 165452 331456 165504
rect 257528 164840 257580 164892
rect 306564 164840 306616 164892
rect 496912 164840 496964 164892
rect 501236 164840 501288 164892
rect 504364 164840 504416 164892
rect 510528 164840 510580 164892
rect 525064 164840 525116 164892
rect 276664 164296 276716 164348
rect 307116 164296 307168 164348
rect 252376 164228 252428 164280
rect 259552 164228 259604 164280
rect 269764 164228 269816 164280
rect 307668 164228 307720 164280
rect 334624 164228 334676 164280
rect 416780 164228 416832 164280
rect 3240 164160 3292 164212
rect 33784 164160 33836 164212
rect 171968 164160 172020 164212
rect 214012 164160 214064 164212
rect 252468 164160 252520 164212
rect 269120 164160 269172 164212
rect 324320 164160 324372 164212
rect 332784 164160 332836 164212
rect 496912 164160 496964 164212
rect 506664 164160 506716 164212
rect 556160 164160 556212 164212
rect 196900 164092 196952 164144
rect 213920 164092 213972 164144
rect 252376 164092 252428 164144
rect 256792 164092 256844 164144
rect 268568 163548 268620 163600
rect 307484 163548 307536 163600
rect 261484 163480 261536 163532
rect 307392 163480 307444 163532
rect 286416 162868 286468 162920
rect 307668 162868 307720 162920
rect 170496 162800 170548 162852
rect 213920 162800 213972 162852
rect 252376 162800 252428 162852
rect 266360 162800 266412 162852
rect 324320 162800 324372 162852
rect 342352 162800 342404 162852
rect 496912 162800 496964 162852
rect 512644 162800 512696 162852
rect 178776 162732 178828 162784
rect 214012 162732 214064 162784
rect 252468 162732 252520 162784
rect 265164 162732 265216 162784
rect 274088 162120 274140 162172
rect 306748 162120 306800 162172
rect 304264 161576 304316 161628
rect 307484 161576 307536 161628
rect 278136 161508 278188 161560
rect 307576 161508 307628 161560
rect 262956 161440 263008 161492
rect 307668 161440 307720 161492
rect 345664 161440 345716 161492
rect 416780 161440 416832 161492
rect 169116 161372 169168 161424
rect 213920 161372 213972 161424
rect 252468 161372 252520 161424
rect 261116 161372 261168 161424
rect 496912 161372 496964 161424
rect 535460 161372 535512 161424
rect 173164 161304 173216 161356
rect 214012 161304 214064 161356
rect 301504 160216 301556 160268
rect 307576 160216 307628 160268
rect 324320 160216 324372 160268
rect 327448 160216 327500 160268
rect 264336 160148 264388 160200
rect 307668 160148 307720 160200
rect 253480 160080 253532 160132
rect 307484 160080 307536 160132
rect 324320 160012 324372 160064
rect 331496 160012 331548 160064
rect 496912 160012 496964 160064
rect 529940 160012 529992 160064
rect 497004 159944 497056 159996
rect 503720 159944 503772 159996
rect 167644 159332 167696 159384
rect 214012 159332 214064 159384
rect 293408 158856 293460 158908
rect 306564 158856 306616 158908
rect 260472 158788 260524 158840
rect 307668 158788 307720 158840
rect 258816 158720 258868 158772
rect 307576 158720 307628 158772
rect 167828 158652 167880 158704
rect 213920 158652 213972 158704
rect 251364 158652 251416 158704
rect 253940 158652 253992 158704
rect 324320 158652 324372 158704
rect 336924 158652 336976 158704
rect 496912 158652 496964 158704
rect 517612 158652 517664 158704
rect 544384 158652 544436 158704
rect 252192 158584 252244 158636
rect 255504 158584 255556 158636
rect 251916 157972 251968 158024
rect 264244 157972 264296 158024
rect 287888 157496 287940 157548
rect 306564 157496 306616 157548
rect 267004 157428 267056 157480
rect 307668 157428 307720 157480
rect 263600 157360 263652 157412
rect 307484 157360 307536 157412
rect 331864 157360 331916 157412
rect 416780 157360 416832 157412
rect 205088 157292 205140 157344
rect 213920 157292 213972 157344
rect 252468 157292 252520 157344
rect 273260 157292 273312 157344
rect 324320 157292 324372 157344
rect 338304 157292 338356 157344
rect 496912 157292 496964 157344
rect 582380 157292 582432 157344
rect 252376 157224 252428 157276
rect 263784 157224 263836 157276
rect 285036 156068 285088 156120
rect 307668 156068 307720 156120
rect 272708 156000 272760 156052
rect 306564 156000 306616 156052
rect 260196 155932 260248 155984
rect 307576 155932 307628 155984
rect 336004 155932 336056 155984
rect 416780 155932 416832 155984
rect 171876 155864 171928 155916
rect 214012 155864 214064 155916
rect 324320 155864 324372 155916
rect 331312 155864 331364 155916
rect 496912 155864 496964 155916
rect 519544 155864 519596 155916
rect 196716 155796 196768 155848
rect 213920 155796 213972 155848
rect 170588 155184 170640 155236
rect 214564 155184 214616 155236
rect 272800 155184 272852 155236
rect 307392 155184 307444 155236
rect 262864 154640 262916 154692
rect 307576 154640 307628 154692
rect 261760 154572 261812 154624
rect 307668 154572 307720 154624
rect 356796 154572 356848 154624
rect 416780 154572 416832 154624
rect 251548 154504 251600 154556
rect 254216 154504 254268 154556
rect 324320 154504 324372 154556
rect 341064 154504 341116 154556
rect 497004 154504 497056 154556
rect 505284 154504 505336 154556
rect 252468 154436 252520 154488
rect 267832 154436 267884 154488
rect 324412 154436 324464 154488
rect 328736 154436 328788 154488
rect 496912 154436 496964 154488
rect 502524 154436 502576 154488
rect 252376 154368 252428 154420
rect 274732 154368 274784 154420
rect 251824 153824 251876 153876
rect 263600 153824 263652 153876
rect 267096 153824 267148 153876
rect 307484 153824 307536 153876
rect 174544 153280 174596 153332
rect 214012 153280 214064 153332
rect 302976 153280 303028 153332
rect 307668 153280 307720 153332
rect 166264 153212 166316 153264
rect 213920 153212 213972 153264
rect 298744 153212 298796 153264
rect 306564 153212 306616 153264
rect 360844 153212 360896 153264
rect 416780 153212 416832 153264
rect 252376 153144 252428 153196
rect 271972 153144 272024 153196
rect 324320 153144 324372 153196
rect 330024 153144 330076 153196
rect 252284 153076 252336 153128
rect 269212 153076 269264 153128
rect 252468 153008 252520 153060
rect 266452 153008 266504 153060
rect 496912 152600 496964 152652
rect 498476 152600 498528 152652
rect 276848 152464 276900 152516
rect 307668 152464 307720 152516
rect 189724 151784 189776 151836
rect 213920 151784 213972 151836
rect 258724 151784 258776 151836
rect 307668 151784 307720 151836
rect 324320 151716 324372 151768
rect 339592 151716 339644 151768
rect 252376 151648 252428 151700
rect 271880 151648 271932 151700
rect 252468 151580 252520 151632
rect 276112 151580 276164 151632
rect 252284 151444 252336 151496
rect 254124 151444 254176 151496
rect 256148 151036 256200 151088
rect 306656 151036 306708 151088
rect 303068 150560 303120 150612
rect 307668 150560 307720 150612
rect 209136 150492 209188 150544
rect 214012 150492 214064 150544
rect 289268 150492 289320 150544
rect 307300 150492 307352 150544
rect 196716 150424 196768 150476
rect 213920 150424 213972 150476
rect 264244 150424 264296 150476
rect 306932 150424 306984 150476
rect 359556 150424 359608 150476
rect 416780 150424 416832 150476
rect 3424 150356 3476 150408
rect 15844 150356 15896 150408
rect 170404 150356 170456 150408
rect 214012 150356 214064 150408
rect 252468 150356 252520 150408
rect 264980 150356 265032 150408
rect 324320 150356 324372 150408
rect 335452 150356 335504 150408
rect 496820 150356 496872 150408
rect 506572 150356 506624 150408
rect 252284 150288 252336 150340
rect 255596 150288 255648 150340
rect 324412 150288 324464 150340
rect 333980 150288 334032 150340
rect 287980 149200 288032 149252
rect 306932 149200 306984 149252
rect 279516 149132 279568 149184
rect 306564 149132 306616 149184
rect 265716 149064 265768 149116
rect 307300 149064 307352 149116
rect 363604 149064 363656 149116
rect 416780 149064 416832 149116
rect 169024 148996 169076 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 278780 148996 278832 149048
rect 324412 148996 324464 149048
rect 342444 148996 342496 149048
rect 496820 148996 496872 149048
rect 505192 148996 505244 149048
rect 252376 148928 252428 148980
rect 254032 148928 254084 148980
rect 324320 148928 324372 148980
rect 329932 148928 329984 148980
rect 286600 147772 286652 147824
rect 307484 147772 307536 147824
rect 257344 147704 257396 147756
rect 307576 147704 307628 147756
rect 256240 147636 256292 147688
rect 307668 147636 307720 147688
rect 369860 147636 369912 147688
rect 416780 147636 416832 147688
rect 252468 147568 252520 147620
rect 280160 147568 280212 147620
rect 324320 147568 324372 147620
rect 352012 147568 352064 147620
rect 496820 147568 496872 147620
rect 510804 147568 510856 147620
rect 252100 147500 252152 147552
rect 255320 147500 255372 147552
rect 249892 147296 249944 147348
rect 249800 147092 249852 147144
rect 300308 146412 300360 146464
rect 307576 146412 307628 146464
rect 209228 146344 209280 146396
rect 214012 146344 214064 146396
rect 269948 146344 270000 146396
rect 307668 146344 307720 146396
rect 176016 146276 176068 146328
rect 213920 146276 213972 146328
rect 254768 146276 254820 146328
rect 307484 146276 307536 146328
rect 356704 146276 356756 146328
rect 416780 146276 416832 146328
rect 252468 146208 252520 146260
rect 273352 146208 273404 146260
rect 324412 146208 324464 146260
rect 350632 146208 350684 146260
rect 252376 146140 252428 146192
rect 270592 146140 270644 146192
rect 324320 146140 324372 146192
rect 328460 146140 328512 146192
rect 496820 145664 496872 145716
rect 499672 145664 499724 145716
rect 255964 145596 256016 145648
rect 306932 145596 306984 145648
rect 254952 145528 255004 145580
rect 307208 145528 307260 145580
rect 171876 144916 171928 144968
rect 213920 144916 213972 144968
rect 296168 144916 296220 144968
rect 306932 144916 306984 144968
rect 252376 144848 252428 144900
rect 262312 144848 262364 144900
rect 252468 144780 252520 144832
rect 260840 144780 260892 144832
rect 169024 144168 169076 144220
rect 214656 144168 214708 144220
rect 264520 144168 264572 144220
rect 307484 144168 307536 144220
rect 507768 144168 507820 144220
rect 512000 144168 512052 144220
rect 280896 143624 280948 143676
rect 306564 143624 306616 143676
rect 187148 143556 187200 143608
rect 213920 143556 213972 143608
rect 253388 143556 253440 143608
rect 307668 143556 307720 143608
rect 342352 143556 342404 143608
rect 416872 143556 416924 143608
rect 496820 143556 496872 143608
rect 507768 143556 507820 143608
rect 252468 143488 252520 143540
rect 265072 143488 265124 143540
rect 324320 143488 324372 143540
rect 332692 143488 332744 143540
rect 342260 143488 342312 143540
rect 416780 143488 416832 143540
rect 252376 143420 252428 143472
rect 258356 143420 258408 143472
rect 257620 142808 257672 142860
rect 307116 142808 307168 142860
rect 333244 142808 333296 142860
rect 342260 142808 342312 142860
rect 211896 142264 211948 142316
rect 214472 142264 214524 142316
rect 283748 142196 283800 142248
rect 307668 142196 307720 142248
rect 181536 142128 181588 142180
rect 213920 142128 213972 142180
rect 253204 142128 253256 142180
rect 307576 142128 307628 142180
rect 496912 142128 496964 142180
rect 513288 142128 513340 142180
rect 324412 142060 324464 142112
rect 349160 142060 349212 142112
rect 353300 142060 353352 142112
rect 416780 142060 416832 142112
rect 496820 142060 496872 142112
rect 512092 142060 512144 142112
rect 519544 142060 519596 142112
rect 324320 141992 324372 142044
rect 328552 141992 328604 142044
rect 253664 141380 253716 141432
rect 307024 141380 307076 141432
rect 496820 141380 496872 141432
rect 516140 141380 516192 141432
rect 174636 140836 174688 140888
rect 214012 140836 214064 140888
rect 290648 140836 290700 140888
rect 307576 140836 307628 140888
rect 170404 140768 170456 140820
rect 213920 140768 213972 140820
rect 254860 140768 254912 140820
rect 307668 140768 307720 140820
rect 352656 140768 352708 140820
rect 353300 140768 353352 140820
rect 252376 140700 252428 140752
rect 277492 140700 277544 140752
rect 496820 140700 496872 140752
rect 502984 140700 503036 140752
rect 252468 140632 252520 140684
rect 276020 140632 276072 140684
rect 167920 140020 167972 140072
rect 209136 140020 209188 140072
rect 516140 140020 516192 140072
rect 580172 140020 580224 140072
rect 252008 139748 252060 139800
rect 260472 139748 260524 139800
rect 294788 139544 294840 139596
rect 307576 139544 307628 139596
rect 210516 139476 210568 139528
rect 214012 139476 214064 139528
rect 260104 139476 260156 139528
rect 307668 139476 307720 139528
rect 206468 139408 206520 139460
rect 213920 139408 213972 139460
rect 256056 139408 256108 139460
rect 307484 139408 307536 139460
rect 367744 139408 367796 139460
rect 416780 139408 416832 139460
rect 252468 139340 252520 139392
rect 280252 139340 280304 139392
rect 496820 139340 496872 139392
rect 514852 139340 514904 139392
rect 324320 139068 324372 139120
rect 325976 139068 326028 139120
rect 202328 138048 202380 138100
rect 214012 138048 214064 138100
rect 286508 138048 286560 138100
rect 307668 138048 307720 138100
rect 170496 137980 170548 138032
rect 213920 137980 213972 138032
rect 250628 137980 250680 138032
rect 307576 137980 307628 138032
rect 3240 137912 3292 137964
rect 14464 137912 14516 137964
rect 252376 137912 252428 137964
rect 281540 137912 281592 137964
rect 324412 137912 324464 137964
rect 346492 137912 346544 137964
rect 496820 137912 496872 137964
rect 520924 137912 520976 137964
rect 252468 137844 252520 137896
rect 267740 137844 267792 137896
rect 324320 137844 324372 137896
rect 338120 137844 338172 137896
rect 252100 137232 252152 137284
rect 267188 137232 267240 137284
rect 275284 137232 275336 137284
rect 307392 137232 307444 137284
rect 253296 136892 253348 136944
rect 253664 136892 253716 136944
rect 268384 136688 268436 136740
rect 307668 136688 307720 136740
rect 198188 136620 198240 136672
rect 213920 136620 213972 136672
rect 250536 136620 250588 136672
rect 307116 136620 307168 136672
rect 370504 136620 370556 136672
rect 416780 136620 416832 136672
rect 252192 136552 252244 136604
rect 296260 136552 296312 136604
rect 324320 136552 324372 136604
rect 352196 136552 352248 136604
rect 496912 136552 496964 136604
rect 508504 136552 508556 136604
rect 252376 136484 252428 136536
rect 285220 136484 285272 136536
rect 496820 136484 496872 136536
rect 502432 136484 502484 136536
rect 252468 136416 252520 136468
rect 277400 136416 277452 136468
rect 252284 136348 252336 136400
rect 265808 136348 265860 136400
rect 295984 135464 296036 135516
rect 307116 135464 307168 135516
rect 284944 135396 284996 135448
rect 307668 135396 307720 135448
rect 207756 135328 207808 135380
rect 214012 135328 214064 135380
rect 283564 135328 283616 135380
rect 307576 135328 307628 135380
rect 178776 135260 178828 135312
rect 213920 135260 213972 135312
rect 265624 135260 265676 135312
rect 307484 135260 307536 135312
rect 376024 135260 376076 135312
rect 416780 135260 416832 135312
rect 252468 135192 252520 135244
rect 280804 135192 280856 135244
rect 340236 135192 340288 135244
rect 417332 135192 417384 135244
rect 252376 135124 252428 135176
rect 263048 135124 263100 135176
rect 324320 135124 324372 135176
rect 350540 135124 350592 135176
rect 324412 135056 324464 135108
rect 346584 135056 346636 135108
rect 276940 134512 276992 134564
rect 307300 134512 307352 134564
rect 300124 133968 300176 134020
rect 307576 133968 307628 134020
rect 177488 133900 177540 133952
rect 213920 133900 213972 133952
rect 282276 133900 282328 133952
rect 307668 133900 307720 133952
rect 252376 133832 252428 133884
rect 283656 133832 283708 133884
rect 374644 133832 374696 133884
rect 419356 133832 419408 133884
rect 496820 133832 496872 133884
rect 503812 133832 503864 133884
rect 252468 133764 252520 133816
rect 260380 133764 260432 133816
rect 324320 133560 324372 133612
rect 327264 133560 327316 133612
rect 260472 133152 260524 133204
rect 306840 133152 306892 133204
rect 386328 133152 386380 133204
rect 419632 133152 419684 133204
rect 304356 132608 304408 132660
rect 306932 132608 306984 132660
rect 297456 132540 297508 132592
rect 307668 132540 307720 132592
rect 254676 132472 254728 132524
rect 307576 132472 307628 132524
rect 252468 132404 252520 132456
rect 300216 132404 300268 132456
rect 411904 132404 411956 132456
rect 417332 132404 417384 132456
rect 252376 132336 252428 132388
rect 285128 132336 285180 132388
rect 252468 132268 252520 132320
rect 268476 132268 268528 132320
rect 301596 131248 301648 131300
rect 307668 131248 307720 131300
rect 180248 131180 180300 131232
rect 214012 131180 214064 131232
rect 289084 131180 289136 131232
rect 306564 131180 306616 131232
rect 171968 131112 172020 131164
rect 213920 131112 213972 131164
rect 278044 131112 278096 131164
rect 307576 131112 307628 131164
rect 252468 131044 252520 131096
rect 297364 131044 297416 131096
rect 324320 131044 324372 131096
rect 349344 131044 349396 131096
rect 496820 131044 496872 131096
rect 509240 131044 509292 131096
rect 252376 130976 252428 131028
rect 264428 130976 264480 131028
rect 252468 130432 252520 130484
rect 260288 130432 260340 130484
rect 297548 129888 297600 129940
rect 307668 129888 307720 129940
rect 205088 129820 205140 129872
rect 214012 129820 214064 129872
rect 294604 129820 294656 129872
rect 307576 129820 307628 129872
rect 173256 129752 173308 129804
rect 213920 129752 213972 129804
rect 261576 129752 261628 129804
rect 307300 129752 307352 129804
rect 252468 129684 252520 129736
rect 269856 129684 269908 129736
rect 324320 129684 324372 129736
rect 334164 129684 334216 129736
rect 496820 129684 496872 129736
rect 514760 129684 514812 129736
rect 252376 129616 252428 129668
rect 257528 129616 257580 129668
rect 252192 129412 252244 129464
rect 257436 129412 257488 129464
rect 297364 128392 297416 128444
rect 307576 128392 307628 128444
rect 273996 128324 274048 128376
rect 307668 128324 307720 128376
rect 252376 128256 252428 128308
rect 287796 128256 287848 128308
rect 324320 128256 324372 128308
rect 338212 128256 338264 128308
rect 382924 128256 382976 128308
rect 417608 128256 417660 128308
rect 496820 128256 496872 128308
rect 507860 128256 507912 128308
rect 252284 128188 252336 128240
rect 271328 128188 271380 128240
rect 324412 128188 324464 128240
rect 330116 128188 330168 128240
rect 252468 128120 252520 128172
rect 261484 128120 261536 128172
rect 270040 127576 270092 127628
rect 307208 127576 307260 127628
rect 525064 127576 525116 127628
rect 580172 127576 580224 127628
rect 287704 127032 287756 127084
rect 306564 127032 306616 127084
rect 173164 126964 173216 127016
rect 213920 126964 213972 127016
rect 271236 126964 271288 127016
rect 307668 126964 307720 127016
rect 252468 126896 252520 126948
rect 268568 126896 268620 126948
rect 251916 126828 251968 126880
rect 254952 126828 255004 126880
rect 496820 126488 496872 126540
rect 499856 126488 499908 126540
rect 292028 125740 292080 125792
rect 307576 125740 307628 125792
rect 176108 125672 176160 125724
rect 213920 125672 213972 125724
rect 268476 125672 268528 125724
rect 307668 125672 307720 125724
rect 57796 125604 57848 125656
rect 65156 125604 65208 125656
rect 167644 125604 167696 125656
rect 214012 125604 214064 125656
rect 254584 125604 254636 125656
rect 306564 125604 306616 125656
rect 252284 125536 252336 125588
rect 276664 125536 276716 125588
rect 324320 125536 324372 125588
rect 347964 125536 348016 125588
rect 496820 125536 496872 125588
rect 517520 125536 517572 125588
rect 252468 125468 252520 125520
rect 269764 125468 269816 125520
rect 324412 125468 324464 125520
rect 343640 125468 343692 125520
rect 252376 125400 252428 125452
rect 253296 125400 253348 125452
rect 252376 124856 252428 124908
rect 305644 124856 305696 124908
rect 302884 124312 302936 124364
rect 307668 124312 307720 124364
rect 193864 124244 193916 124296
rect 214012 124244 214064 124296
rect 280804 124244 280856 124296
rect 307576 124244 307628 124296
rect 185676 124176 185728 124228
rect 213920 124176 213972 124228
rect 279424 124176 279476 124228
rect 307300 124176 307352 124228
rect 252468 124108 252520 124160
rect 274088 124108 274140 124160
rect 324320 124108 324372 124160
rect 357440 124108 357492 124160
rect 496912 124108 496964 124160
rect 505100 124108 505152 124160
rect 324412 124040 324464 124092
rect 343916 124040 343968 124092
rect 496820 124040 496872 124092
rect 499764 124040 499816 124092
rect 252100 123156 252152 123208
rect 256240 123156 256292 123208
rect 272616 122952 272668 123004
rect 307576 122952 307628 123004
rect 184296 122884 184348 122936
rect 214012 122884 214064 122936
rect 298836 122884 298888 122936
rect 307668 122884 307720 122936
rect 56508 122816 56560 122868
rect 66076 122816 66128 122868
rect 170588 122816 170640 122868
rect 213920 122816 213972 122868
rect 252468 122748 252520 122800
rect 304264 122748 304316 122800
rect 324412 122748 324464 122800
rect 347872 122748 347924 122800
rect 382188 122748 382240 122800
rect 416780 122748 416832 122800
rect 496820 122748 496872 122800
rect 521660 122748 521712 122800
rect 252376 122680 252428 122732
rect 278136 122680 278188 122732
rect 324320 122680 324372 122732
rect 345296 122680 345348 122732
rect 252284 122612 252336 122664
rect 262956 122612 263008 122664
rect 182916 121524 182968 121576
rect 213920 121524 213972 121576
rect 293316 121524 293368 121576
rect 307576 121524 307628 121576
rect 167828 121456 167880 121508
rect 214012 121456 214064 121508
rect 285128 121456 285180 121508
rect 307668 121456 307720 121508
rect 252468 121388 252520 121440
rect 301504 121388 301556 121440
rect 324412 121388 324464 121440
rect 356060 121388 356112 121440
rect 388444 121388 388496 121440
rect 416780 121388 416832 121440
rect 252376 121320 252428 121372
rect 264336 121320 264388 121372
rect 324320 121320 324372 121372
rect 328644 121320 328696 121372
rect 252284 121252 252336 121304
rect 253480 121252 253532 121304
rect 304448 120232 304500 120284
rect 307576 120232 307628 120284
rect 178868 120164 178920 120216
rect 213920 120164 213972 120216
rect 276664 120164 276716 120216
rect 307668 120164 307720 120216
rect 174728 120096 174780 120148
rect 214012 120096 214064 120148
rect 253296 120096 253348 120148
rect 307484 120096 307536 120148
rect 252468 120028 252520 120080
rect 293408 120028 293460 120080
rect 496820 119620 496872 119672
rect 499580 119620 499632 119672
rect 252376 119552 252428 119604
rect 258816 119552 258868 119604
rect 170680 118804 170732 118856
rect 214012 118804 214064 118856
rect 172060 118736 172112 118788
rect 213920 118736 213972 118788
rect 300400 118736 300452 118788
rect 307668 118736 307720 118788
rect 251916 118668 251968 118720
rect 254860 118668 254912 118720
rect 293224 118668 293276 118720
rect 307576 118668 307628 118720
rect 252468 118600 252520 118652
rect 287888 118600 287940 118652
rect 324412 118600 324464 118652
rect 345204 118600 345256 118652
rect 252376 118532 252428 118584
rect 267004 118532 267056 118584
rect 324320 118532 324372 118584
rect 343824 118532 343876 118584
rect 496820 118396 496872 118448
rect 501144 118396 501196 118448
rect 171784 117920 171836 117972
rect 209136 117920 209188 117972
rect 252008 117920 252060 117972
rect 300308 117920 300360 117972
rect 496820 117648 496872 117700
rect 500960 117648 501012 117700
rect 287796 117512 287848 117564
rect 306748 117512 306800 117564
rect 301688 117444 301740 117496
rect 307576 117444 307628 117496
rect 173440 117376 173492 117428
rect 214012 117376 214064 117428
rect 292120 117376 292172 117428
rect 307484 117376 307536 117428
rect 169116 117308 169168 117360
rect 213920 117308 213972 117360
rect 304264 117308 304316 117360
rect 307668 117308 307720 117360
rect 252284 117240 252336 117292
rect 285036 117240 285088 117292
rect 324412 117240 324464 117292
rect 334072 117240 334124 117292
rect 342904 117240 342956 117292
rect 416780 117240 416832 117292
rect 496912 117240 496964 117292
rect 510712 117240 510764 117292
rect 252468 117172 252520 117224
rect 272800 117172 272852 117224
rect 324320 117172 324372 117224
rect 345112 117172 345164 117224
rect 252376 117104 252428 117156
rect 260196 117104 260248 117156
rect 301504 116084 301556 116136
rect 307484 116084 307536 116136
rect 198280 116016 198332 116068
rect 214012 116016 214064 116068
rect 272524 116016 272576 116068
rect 307576 116016 307628 116068
rect 192576 115948 192628 116000
rect 213920 115948 213972 116000
rect 269856 115948 269908 116000
rect 307668 115948 307720 116000
rect 252468 115880 252520 115932
rect 272708 115880 272760 115932
rect 324320 115880 324372 115932
rect 339500 115880 339552 115932
rect 252376 115812 252428 115864
rect 262864 115812 262916 115864
rect 324412 115812 324464 115864
rect 336740 115812 336792 115864
rect 196808 114588 196860 114640
rect 214012 114588 214064 114640
rect 296260 114588 296312 114640
rect 307576 114588 307628 114640
rect 177580 114520 177632 114572
rect 213920 114520 213972 114572
rect 278136 114520 278188 114572
rect 307668 114520 307720 114572
rect 252284 114452 252336 114504
rect 298744 114452 298796 114504
rect 324320 114452 324372 114504
rect 340972 114452 341024 114504
rect 252468 114384 252520 114436
rect 267096 114384 267148 114436
rect 324412 114384 324464 114436
rect 336832 114384 336884 114436
rect 252376 114316 252428 114368
rect 261760 114316 261812 114368
rect 251824 113772 251876 113824
rect 254768 113772 254820 113824
rect 300308 113296 300360 113348
rect 307668 113296 307720 113348
rect 196900 113228 196952 113280
rect 213920 113228 213972 113280
rect 267004 113228 267056 113280
rect 306748 113228 306800 113280
rect 169300 113160 169352 113212
rect 214012 113160 214064 113212
rect 261484 113160 261536 113212
rect 307576 113160 307628 113212
rect 252468 113092 252520 113144
rect 302976 113092 303028 113144
rect 324320 113092 324372 113144
rect 335360 113092 335412 113144
rect 349252 113092 349304 113144
rect 367744 113092 367796 113144
rect 395344 113092 395396 113144
rect 416780 113092 416832 113144
rect 252376 113024 252428 113076
rect 276848 113024 276900 113076
rect 252468 112888 252520 112940
rect 256148 112888 256200 112940
rect 322940 112412 322992 112464
rect 349252 112412 349304 112464
rect 200948 111868 201000 111920
rect 213920 111868 213972 111920
rect 286416 111868 286468 111920
rect 307576 111868 307628 111920
rect 174820 111800 174872 111852
rect 214012 111800 214064 111852
rect 276756 111800 276808 111852
rect 307668 111800 307720 111852
rect 496912 111800 496964 111852
rect 499580 111800 499632 111852
rect 167920 111732 167972 111784
rect 196716 111732 196768 111784
rect 252468 111732 252520 111784
rect 308496 111732 308548 111784
rect 371884 111732 371936 111784
rect 416780 111732 416832 111784
rect 496820 111732 496872 111784
rect 506480 111732 506532 111784
rect 252376 111664 252428 111716
rect 257620 111664 257672 111716
rect 3424 110984 3476 111036
rect 7564 110984 7616 111036
rect 252468 110644 252520 110696
rect 258724 110644 258776 110696
rect 289360 110576 289412 110628
rect 307484 110576 307536 110628
rect 173348 110508 173400 110560
rect 213920 110508 213972 110560
rect 257436 110508 257488 110560
rect 307576 110508 307628 110560
rect 166356 110440 166408 110492
rect 214012 110440 214064 110492
rect 250444 110440 250496 110492
rect 307668 110440 307720 110492
rect 252284 110372 252336 110424
rect 303068 110372 303120 110424
rect 324320 110372 324372 110424
rect 332876 110372 332928 110424
rect 377404 110372 377456 110424
rect 416780 110372 416832 110424
rect 496820 110372 496872 110424
rect 510620 110372 510672 110424
rect 252468 110304 252520 110356
rect 289268 110304 289320 110356
rect 252376 110236 252428 110288
rect 264244 110236 264296 110288
rect 324412 109692 324464 109744
rect 329840 109692 329892 109744
rect 302976 109148 303028 109200
rect 306748 109148 306800 109200
rect 178960 109080 179012 109132
rect 213920 109080 213972 109132
rect 294696 109080 294748 109132
rect 307576 109080 307628 109132
rect 166448 109012 166500 109064
rect 214012 109012 214064 109064
rect 285036 109012 285088 109064
rect 307668 109012 307720 109064
rect 252284 108944 252336 108996
rect 287980 108944 288032 108996
rect 252468 108876 252520 108928
rect 279516 108876 279568 108928
rect 252376 108808 252428 108860
rect 265716 108808 265768 108860
rect 324320 108740 324372 108792
rect 327172 108740 327224 108792
rect 282368 107856 282420 107908
rect 307484 107856 307536 107908
rect 169208 107720 169260 107772
rect 213920 107720 213972 107772
rect 287888 107720 287940 107772
rect 307668 107720 307720 107772
rect 167920 107652 167972 107704
rect 214012 107652 214064 107704
rect 303068 107652 303120 107704
rect 306932 107652 306984 107704
rect 252468 107584 252520 107636
rect 286600 107584 286652 107636
rect 324320 107584 324372 107636
rect 340880 107584 340932 107636
rect 403716 107584 403768 107636
rect 416780 107584 416832 107636
rect 252376 107516 252428 107568
rect 257344 107516 257396 107568
rect 290556 106428 290608 106480
rect 307576 106428 307628 106480
rect 181628 106360 181680 106412
rect 213920 106360 213972 106412
rect 269764 106360 269816 106412
rect 307484 106360 307536 106412
rect 169024 106292 169076 106344
rect 214012 106292 214064 106344
rect 249064 106292 249116 106344
rect 307668 106292 307720 106344
rect 252468 106224 252520 106276
rect 255964 106224 256016 106276
rect 341524 106224 341576 106276
rect 416780 106224 416832 106276
rect 496820 106224 496872 106276
rect 507952 106224 508004 106276
rect 252192 105612 252244 105664
rect 283748 105612 283800 105664
rect 252284 105544 252336 105596
rect 296168 105544 296220 105596
rect 300216 105000 300268 105052
rect 307484 105000 307536 105052
rect 283656 104932 283708 104984
rect 307576 104932 307628 104984
rect 202420 104864 202472 104916
rect 213920 104864 213972 104916
rect 264336 104864 264388 104916
rect 307668 104864 307720 104916
rect 252468 104796 252520 104848
rect 269948 104796 270000 104848
rect 359464 104796 359516 104848
rect 416780 104796 416832 104848
rect 252376 104728 252428 104780
rect 264520 104728 264572 104780
rect 267096 103640 267148 103692
rect 306748 103640 306800 103692
rect 264244 103572 264296 103624
rect 307576 103572 307628 103624
rect 188436 103504 188488 103556
rect 213920 103504 213972 103556
rect 264428 103504 264480 103556
rect 307668 103504 307720 103556
rect 407764 103436 407816 103488
rect 416780 103436 416832 103488
rect 252468 103368 252520 103420
rect 275284 103368 275336 103420
rect 252376 103300 252428 103352
rect 280896 103300 280948 103352
rect 251180 102892 251232 102944
rect 253388 102892 253440 102944
rect 330484 102756 330536 102808
rect 376024 102756 376076 102808
rect 296168 102280 296220 102332
rect 306748 102280 306800 102332
rect 207848 102212 207900 102264
rect 213920 102212 213972 102264
rect 280988 102212 281040 102264
rect 307668 102212 307720 102264
rect 192668 102144 192720 102196
rect 214012 102144 214064 102196
rect 262864 102144 262916 102196
rect 307576 102144 307628 102196
rect 252468 102076 252520 102128
rect 276940 102076 276992 102128
rect 252192 101396 252244 101448
rect 256056 101396 256108 101448
rect 298744 100852 298796 100904
rect 307576 100852 307628 100904
rect 206560 100784 206612 100836
rect 214012 100784 214064 100836
rect 260196 100784 260248 100836
rect 307668 100784 307720 100836
rect 200856 100716 200908 100768
rect 213920 100716 213972 100768
rect 258724 100716 258776 100768
rect 306932 100716 306984 100768
rect 252376 100648 252428 100700
rect 290648 100648 290700 100700
rect 360200 100648 360252 100700
rect 370504 100648 370556 100700
rect 378784 100648 378836 100700
rect 494060 100648 494112 100700
rect 519544 100648 519596 100700
rect 580172 100648 580224 100700
rect 252468 100580 252520 100632
rect 270040 100580 270092 100632
rect 406384 100580 406436 100632
rect 496820 100580 496872 100632
rect 252284 100512 252336 100564
rect 260472 100512 260524 100564
rect 167736 99968 167788 100020
rect 214564 99968 214616 100020
rect 325700 99968 325752 100020
rect 360200 99968 360252 100020
rect 254768 99492 254820 99544
rect 307576 99492 307628 99544
rect 275284 99424 275336 99476
rect 307668 99424 307720 99476
rect 164884 99356 164936 99408
rect 213920 99356 213972 99408
rect 252468 99288 252520 99340
rect 261668 99288 261720 99340
rect 419632 99288 419684 99340
rect 580264 99288 580316 99340
rect 251916 99220 251968 99272
rect 254952 99220 255004 99272
rect 400864 99220 400916 99272
rect 493968 99220 494020 99272
rect 410616 99152 410668 99204
rect 496912 99152 496964 99204
rect 171784 98608 171836 98660
rect 214012 98608 214064 98660
rect 324412 98608 324464 98660
rect 331588 98608 331640 98660
rect 264520 98064 264572 98116
rect 307668 98064 307720 98116
rect 212448 97996 212500 98048
rect 213920 97996 213972 98048
rect 251916 97996 251968 98048
rect 306748 97996 306800 98048
rect 3424 97928 3476 97980
rect 17224 97928 17276 97980
rect 324320 97928 324372 97980
rect 346400 97928 346452 97980
rect 399484 97928 399536 97980
rect 494336 97928 494388 97980
rect 413284 97860 413336 97912
rect 497004 97860 497056 97912
rect 420184 97316 420236 97368
rect 427728 97316 427780 97368
rect 166540 97248 166592 97300
rect 214656 97248 214708 97300
rect 252008 97248 252060 97300
rect 259368 97248 259420 97300
rect 308404 97248 308456 97300
rect 421564 97248 421616 97300
rect 458916 97248 458968 97300
rect 467104 97248 467156 97300
rect 492496 97248 492548 97300
rect 439504 96908 439556 96960
rect 440884 96908 440936 96960
rect 454040 96908 454092 96960
rect 455052 96908 455104 96960
rect 461584 96908 461636 96960
rect 464896 96908 464948 96960
rect 465724 96908 465776 96960
rect 467288 96908 467340 96960
rect 472624 96908 472676 96960
rect 474556 96908 474608 96960
rect 481640 96908 481692 96960
rect 482652 96908 482704 96960
rect 486424 96908 486476 96960
rect 487712 96908 487764 96960
rect 289268 96772 289320 96824
rect 307668 96772 307720 96824
rect 417424 96772 417476 96824
rect 420552 96772 420604 96824
rect 258816 96704 258868 96756
rect 306932 96704 306984 96756
rect 253388 96636 253440 96688
rect 307576 96636 307628 96688
rect 186228 96568 186280 96620
rect 321468 96568 321520 96620
rect 350540 96568 350592 96620
rect 351184 96568 351236 96620
rect 501052 96568 501104 96620
rect 282184 96500 282236 96552
rect 321560 96500 321612 96552
rect 309784 96432 309836 96484
rect 321652 96432 321704 96484
rect 203616 95208 203668 95260
rect 213920 95208 213972 95260
rect 247684 95208 247736 95260
rect 307668 95208 307720 95260
rect 203524 95140 203576 95192
rect 321376 95140 321428 95192
rect 389824 95140 389876 95192
rect 499580 95140 499632 95192
rect 204168 95072 204220 95124
rect 321836 95072 321888 95124
rect 206284 95004 206336 95056
rect 321744 95004 321796 95056
rect 290464 94936 290516 94988
rect 323032 94936 323084 94988
rect 296076 94868 296128 94920
rect 323216 94868 323268 94920
rect 304908 94800 304960 94852
rect 324504 94800 324556 94852
rect 129556 94460 129608 94512
rect 214012 94460 214064 94512
rect 333980 94460 334032 94512
rect 494244 94460 494296 94512
rect 124496 94052 124548 94104
rect 174636 94052 174688 94104
rect 112352 93984 112404 94036
rect 172060 93984 172112 94036
rect 122840 93916 122892 93968
rect 185676 93916 185728 93968
rect 85580 93848 85632 93900
rect 212448 93848 212500 93900
rect 56508 93780 56560 93832
rect 192668 93780 192720 93832
rect 308404 93780 308456 93832
rect 420920 93780 420972 93832
rect 57796 93712 57848 93764
rect 188436 93712 188488 93764
rect 291936 93712 291988 93764
rect 323124 93712 323176 93764
rect 151728 93304 151780 93356
rect 166264 93304 166316 93356
rect 123208 93236 123260 93288
rect 170404 93236 170456 93288
rect 134708 93168 134760 93220
rect 214748 93168 214800 93220
rect 320824 93168 320876 93220
rect 420184 93168 420236 93220
rect 100576 93100 100628 93152
rect 200948 93100 201000 93152
rect 419172 93100 419224 93152
rect 580264 93100 580316 93152
rect 88064 92420 88116 92472
rect 171784 92420 171836 92472
rect 202144 92420 202196 92472
rect 324596 92420 324648 92472
rect 119344 92352 119396 92404
rect 202328 92352 202380 92404
rect 86776 92284 86828 92336
rect 129556 92284 129608 92336
rect 133144 92284 133196 92336
rect 176016 92284 176068 92336
rect 129464 92216 129516 92268
rect 166540 92216 166592 92268
rect 110696 92148 110748 92200
rect 134708 92148 134760 92200
rect 152096 92148 152148 92200
rect 189724 92148 189776 92200
rect 136088 92080 136140 92132
rect 167736 92080 167788 92132
rect 199476 91740 199528 91792
rect 313280 91740 313332 91792
rect 84844 91128 84896 91180
rect 111156 91128 111208 91180
rect 74816 91060 74868 91112
rect 111064 91060 111116 91112
rect 67640 90992 67692 91044
rect 206560 90992 206612 91044
rect 210424 90992 210476 91044
rect 333980 90992 334032 91044
rect 110052 90924 110104 90976
rect 198280 90924 198332 90976
rect 113824 90856 113876 90908
rect 178776 90856 178828 90908
rect 119896 90788 119948 90840
rect 167828 90788 167880 90840
rect 151544 90720 151596 90772
rect 174544 90720 174596 90772
rect 289176 90312 289228 90364
rect 321560 90312 321612 90364
rect 465080 90312 465132 90364
rect 88984 89632 89036 89684
rect 164884 89632 164936 89684
rect 134892 89564 134944 89616
rect 209228 89564 209280 89616
rect 102048 89496 102100 89548
rect 174820 89496 174872 89548
rect 111616 89428 111668 89480
rect 173440 89428 173492 89480
rect 118056 89360 118108 89412
rect 170496 89360 170548 89412
rect 120908 89292 120960 89344
rect 170588 89292 170640 89344
rect 170404 88952 170456 89004
rect 307300 88952 307352 89004
rect 316040 88952 316092 89004
rect 333244 88952 333296 89004
rect 334716 88952 334768 89004
rect 462320 88952 462372 89004
rect 122104 88272 122156 88324
rect 210516 88272 210568 88324
rect 124128 88204 124180 88256
rect 193864 88204 193916 88256
rect 97448 88136 97500 88188
rect 166448 88136 166500 88188
rect 104440 88068 104492 88120
rect 169300 88068 169352 88120
rect 151636 88000 151688 88052
rect 213368 88000 213420 88052
rect 115296 87932 115348 87984
rect 170680 87932 170732 87984
rect 318800 87660 318852 87712
rect 352656 87660 352708 87712
rect 352564 87592 352616 87644
rect 456800 87592 456852 87644
rect 90640 86912 90692 86964
rect 202420 86912 202472 86964
rect 353300 86912 353352 86964
rect 421564 86912 421616 86964
rect 504364 86912 504416 86964
rect 580172 86912 580224 86964
rect 126060 86844 126112 86896
rect 211896 86844 211948 86896
rect 107936 86776 107988 86828
rect 192576 86776 192628 86828
rect 97080 86708 97132 86760
rect 173164 86708 173216 86760
rect 115756 86640 115808 86692
rect 178868 86640 178920 86692
rect 342260 86300 342312 86352
rect 353300 86300 353352 86352
rect 178684 86232 178736 86284
rect 253204 86232 253256 86284
rect 311900 86232 311952 86284
rect 342352 86232 342404 86284
rect 349804 86232 349856 86284
rect 455420 86232 455472 86284
rect 3148 85484 3200 85536
rect 32404 85484 32456 85536
rect 67732 85484 67784 85536
rect 214840 85484 214892 85536
rect 104624 85416 104676 85468
rect 171968 85416 172020 85468
rect 100116 85348 100168 85400
rect 166356 85348 166408 85400
rect 110144 85280 110196 85332
rect 169116 85280 169168 85332
rect 117136 85212 117188 85264
rect 174728 85212 174780 85264
rect 126704 85144 126756 85196
rect 181536 85144 181588 85196
rect 336096 84804 336148 84856
rect 460940 84804 460992 84856
rect 66076 84124 66128 84176
rect 214564 84124 214616 84176
rect 103336 84056 103388 84108
rect 196900 84056 196952 84108
rect 92388 83988 92440 84040
rect 181628 83988 181680 84040
rect 125508 83920 125560 83972
rect 176108 83920 176160 83972
rect 131028 83852 131080 83904
rect 171876 83852 171928 83904
rect 192484 83444 192536 83496
rect 315304 83444 315356 83496
rect 332048 83444 332100 83496
rect 463700 83444 463752 83496
rect 103428 82764 103480 82816
rect 205088 82764 205140 82816
rect 95056 82696 95108 82748
rect 169208 82696 169260 82748
rect 106188 82628 106240 82680
rect 177580 82628 177632 82680
rect 122748 82560 122800 82612
rect 184296 82560 184348 82612
rect 126888 82492 126940 82544
rect 167644 82492 167696 82544
rect 216036 82220 216088 82272
rect 239404 82220 239456 82272
rect 207664 82152 207716 82204
rect 232504 82152 232556 82204
rect 195336 82084 195388 82136
rect 246304 82084 246356 82136
rect 324320 82084 324372 82136
rect 461584 82084 461636 82136
rect 107476 81336 107528 81388
rect 196808 81336 196860 81388
rect 351920 81336 351972 81388
rect 465724 81336 465776 81388
rect 121368 81268 121420 81320
rect 206468 81268 206520 81320
rect 95148 81200 95200 81252
rect 167920 81200 167972 81252
rect 118608 81132 118660 81184
rect 182916 81132 182968 81184
rect 187056 80656 187108 80708
rect 307116 80656 307168 80708
rect 317420 80656 317472 80708
rect 351920 80656 351972 80708
rect 114376 79976 114428 80028
rect 213460 79976 213512 80028
rect 96528 79908 96580 79960
rect 178960 79908 179012 79960
rect 93768 79840 93820 79892
rect 169024 79840 169076 79892
rect 101956 79772 102008 79824
rect 173256 79772 173308 79824
rect 209044 79432 209096 79484
rect 238024 79432 238076 79484
rect 198096 79364 198148 79416
rect 244924 79364 244976 79416
rect 173164 79296 173216 79348
rect 307208 79296 307260 79348
rect 309784 79296 309836 79348
rect 470600 79296 470652 79348
rect 110328 78616 110380 78668
rect 177488 78616 177540 78668
rect 339408 78616 339460 78668
rect 471980 78616 472032 78668
rect 128268 78548 128320 78600
rect 187148 78548 187200 78600
rect 269948 78072 270000 78124
rect 334624 78072 334676 78124
rect 196624 78004 196676 78056
rect 279516 78004 279568 78056
rect 45560 77936 45612 77988
rect 297548 77936 297600 77988
rect 303620 77256 303672 77308
rect 339408 77256 339460 77308
rect 111156 77188 111208 77240
rect 200856 77188 200908 77240
rect 99288 77120 99340 77172
rect 173348 77120 173400 77172
rect 199384 76644 199436 76696
rect 86960 76576 87012 76628
rect 285128 76576 285180 76628
rect 287060 76576 287112 76628
rect 336004 76576 336056 76628
rect 2780 76508 2832 76560
rect 294788 76508 294840 76560
rect 20 75828 72 75880
rect 1308 75828 1360 75880
rect 249156 75828 249208 75880
rect 111064 75760 111116 75812
rect 203616 75760 203668 75812
rect 69020 75216 69072 75268
rect 300400 75216 300452 75268
rect 63408 75148 63460 75200
rect 309876 75148 309928 75200
rect 312544 75148 312596 75200
rect 469220 75148 469272 75200
rect 343732 74468 343784 74520
rect 459560 74468 459612 74520
rect 110420 73924 110472 73976
rect 257436 73924 257488 73976
rect 80060 73856 80112 73908
rect 304448 73856 304500 73908
rect 61936 73788 61988 73840
rect 338856 73788 338908 73840
rect 339500 73176 339552 73228
rect 343732 73176 343784 73228
rect 419356 73108 419408 73160
rect 579988 73108 580040 73160
rect 352104 73040 352156 73092
rect 426532 73040 426584 73092
rect 114560 72564 114612 72616
rect 289360 72564 289412 72616
rect 44088 72496 44140 72548
rect 240784 72496 240836 72548
rect 59360 72428 59412 72480
rect 301688 72428 301740 72480
rect 345756 71748 345808 71800
rect 352104 71748 352156 71800
rect 3424 71680 3476 71732
rect 52368 71680 52420 71732
rect 495716 71680 495768 71732
rect 41328 71612 41380 71664
rect 332048 71612 332100 71664
rect 186964 71068 187016 71120
rect 333244 71068 333296 71120
rect 84200 71000 84252 71052
rect 253296 71000 253348 71052
rect 331312 70524 331364 70576
rect 332048 70524 332100 70576
rect 333244 70388 333296 70440
rect 334716 70388 334768 70440
rect 204996 69776 205048 69828
rect 289820 69776 289872 69828
rect 63316 69708 63368 69760
rect 292580 69708 292632 69760
rect 40040 69640 40092 69692
rect 280988 69640 281040 69692
rect 297548 69640 297600 69692
rect 472624 69640 472676 69692
rect 60556 68960 60608 69012
rect 335360 68960 335412 69012
rect 336096 68960 336148 69012
rect 292580 68892 292632 68944
rect 474740 68892 474792 68944
rect 93860 68348 93912 68400
rect 293316 68348 293368 68400
rect 20720 68280 20772 68332
rect 254768 68280 254820 68332
rect 2688 67532 2740 67584
rect 5448 67532 5500 67584
rect 251364 67532 251416 67584
rect 289820 67532 289872 67584
rect 476120 67532 476172 67584
rect 180156 66920 180208 66972
rect 257344 66920 257396 66972
rect 262220 66920 262272 66972
rect 338764 66920 338816 66972
rect 62120 66852 62172 66904
rect 292120 66852 292172 66904
rect 61844 66172 61896 66224
rect 269120 66172 269172 66224
rect 269948 66172 270000 66224
rect 285680 66172 285732 66224
rect 286324 66172 286376 66224
rect 477500 66172 477552 66224
rect 121460 65560 121512 65612
rect 305920 65560 305972 65612
rect 31760 65492 31812 65544
rect 273996 65492 274048 65544
rect 60648 64812 60700 64864
rect 273260 64812 273312 64864
rect 279516 64812 279568 64864
rect 480260 64812 480312 64864
rect 273260 64404 273312 64456
rect 274088 64404 274140 64456
rect 73160 64132 73212 64184
rect 293224 64132 293276 64184
rect 278780 63520 278832 63572
rect 279516 63520 279568 63572
rect 98000 62840 98052 62892
rect 298836 62840 298888 62892
rect 278228 62772 278280 62824
rect 481732 62772 481784 62824
rect 274640 62024 274692 62076
rect 481640 62024 481692 62076
rect 104900 61480 104952 61532
rect 272616 61480 272668 61532
rect 59176 61412 59228 61464
rect 285128 61412 285180 61464
rect 17960 61344 18012 61396
rect 300308 61344 300360 61396
rect 271880 60732 271932 60784
rect 274640 60732 274692 60784
rect 513288 60664 513340 60716
rect 580172 60664 580224 60716
rect 118700 60052 118752 60104
rect 279424 60052 279476 60104
rect 15200 59984 15252 60036
rect 258816 59984 258868 60036
rect 268568 59984 268620 60036
rect 483020 59984 483072 60036
rect 3056 59304 3108 59356
rect 25504 59304 25556 59356
rect 211804 58828 211856 58880
rect 264980 58828 265032 58880
rect 74540 58760 74592 58812
rect 254676 58760 254728 58812
rect 484400 58760 484452 58812
rect 56600 58692 56652 58744
rect 278044 58692 278096 58744
rect 57888 58624 57940 58676
rect 332600 58624 332652 58676
rect 261668 57876 261720 57928
rect 485780 57876 485832 57928
rect 332600 57740 332652 57792
rect 414664 57808 414716 57860
rect 260840 57672 260892 57724
rect 261668 57672 261720 57724
rect 102140 57332 102192 57384
rect 305828 57332 305880 57384
rect 52460 57264 52512 57316
rect 261576 57264 261628 57316
rect 6920 57196 6972 57248
rect 264520 57196 264572 57248
rect 209136 56040 209188 56092
rect 253940 56040 253992 56092
rect 51080 55972 51132 56024
rect 264428 55972 264480 56024
rect 67640 55904 67692 55956
rect 297456 55904 297508 55956
rect 117320 55836 117372 55888
rect 250628 55836 250680 55888
rect 253940 55836 253992 55888
rect 488540 55836 488592 55888
rect 78680 54680 78732 54732
rect 290556 54680 290608 54732
rect 70400 54612 70452 54664
rect 304356 54612 304408 54664
rect 253020 54544 253072 54596
rect 489920 54544 489972 54596
rect 11060 54476 11112 54528
rect 253388 54476 253440 54528
rect 60740 53184 60792 53236
rect 264336 53184 264388 53236
rect 4160 53116 4212 53168
rect 247684 53116 247736 53168
rect 247776 53116 247828 53168
rect 491300 53116 491352 53168
rect 37280 53048 37332 53100
rect 296260 53048 296312 53100
rect 243544 52368 243596 52420
rect 467104 52368 467156 52420
rect 35808 52300 35860 52352
rect 252652 52300 252704 52352
rect 253020 52300 253072 52352
rect 202236 52232 202288 52284
rect 247040 52232 247092 52284
rect 247776 52232 247828 52284
rect 69112 51688 69164 51740
rect 300216 51688 300268 51740
rect 242900 51076 242952 51128
rect 243544 51076 243596 51128
rect 240784 51008 240836 51060
rect 492680 51008 492732 51060
rect 240140 50532 240192 50584
rect 240784 50532 240836 50584
rect 71780 50464 71832 50516
rect 249064 50464 249116 50516
rect 85580 50396 85632 50448
rect 300124 50396 300176 50448
rect 41420 50328 41472 50380
rect 269856 50328 269908 50380
rect 311164 49648 311216 49700
rect 312544 49648 312596 49700
rect 124220 49104 124272 49156
rect 260104 49104 260156 49156
rect 267188 49104 267240 49156
rect 353944 49104 353996 49156
rect 64604 49036 64656 49088
rect 311164 49036 311216 49088
rect 9680 48968 9732 49020
rect 292028 48968 292080 49020
rect 349160 48968 349212 49020
rect 495624 48968 495676 49020
rect 367836 48220 367888 48272
rect 495532 48220 495584 48272
rect 122840 47676 122892 47728
rect 268476 47676 268528 47728
rect 273904 47676 273956 47728
rect 276020 47676 276072 47728
rect 345664 47676 345716 47728
rect 34520 47608 34572 47660
rect 278136 47608 278188 47660
rect 64696 47540 64748 47592
rect 327724 47540 327776 47592
rect 345020 47540 345072 47592
rect 367100 47540 367152 47592
rect 367836 47540 367888 47592
rect 206376 46860 206428 46912
rect 349160 46860 349212 46912
rect 555424 46860 555476 46912
rect 580172 46860 580224 46912
rect 45468 46248 45520 46300
rect 291200 46248 291252 46300
rect 356796 46248 356848 46300
rect 2872 46180 2924 46232
rect 289268 46180 289320 46232
rect 340880 46180 340932 46232
rect 494152 46180 494204 46232
rect 3424 45500 3476 45552
rect 22744 45500 22796 45552
rect 67180 45500 67232 45552
rect 320180 45500 320232 45552
rect 362960 45500 363012 45552
rect 498200 45500 498252 45552
rect 338856 45432 338908 45484
rect 422300 45432 422352 45484
rect 320180 45228 320232 45280
rect 320824 45228 320876 45280
rect 115940 44888 115992 44940
rect 280804 44888 280856 44940
rect 62028 44820 62080 44872
rect 282184 44820 282236 44872
rect 343640 44820 343692 44872
rect 362960 44820 363012 44872
rect 338120 44140 338172 44192
rect 338856 44140 338908 44192
rect 106280 43460 106332 43512
rect 250536 43460 250588 43512
rect 85672 43392 85724 43444
rect 287888 43392 287940 43444
rect 317328 43392 317380 43444
rect 427820 43392 427872 43444
rect 195244 42712 195296 42764
rect 266360 42712 266412 42764
rect 266360 42100 266412 42152
rect 267188 42100 267240 42152
rect 305000 42100 305052 42152
rect 369860 42100 369912 42152
rect 313924 42032 313976 42084
rect 429200 42032 429252 42084
rect 284300 41352 284352 41404
rect 285128 41352 285180 41404
rect 331864 41352 331916 41404
rect 113180 40740 113232 40792
rect 286508 40740 286560 40792
rect 96620 40672 96672 40724
rect 285036 40672 285088 40724
rect 309876 40672 309928 40724
rect 430580 40672 430632 40724
rect 34428 39448 34480 39500
rect 133144 39448 133196 39500
rect 185584 39448 185636 39500
rect 299572 39448 299624 39500
rect 300676 39448 300728 39500
rect 110512 39380 110564 39432
rect 268384 39380 268436 39432
rect 302240 39380 302292 39432
rect 433340 39380 433392 39432
rect 89720 39312 89772 39364
rect 305736 39312 305788 39364
rect 182824 38564 182876 38616
rect 296720 38564 296772 38616
rect 297548 38564 297600 38616
rect 239404 38496 239456 38548
rect 302240 38496 302292 38548
rect 313280 38496 313332 38548
rect 434720 38564 434772 38616
rect 299480 37952 299532 38004
rect 313280 37952 313332 38004
rect 93952 37884 94004 37936
rect 303068 37884 303120 37936
rect 213276 36660 213328 36712
rect 295340 36660 295392 36712
rect 29000 36592 29052 36644
rect 260196 36592 260248 36644
rect 436192 36592 436244 36644
rect 44180 36524 44232 36576
rect 296168 36524 296220 36576
rect 22100 35164 22152 35216
rect 261484 35164 261536 35216
rect 295432 35164 295484 35216
rect 436284 35164 436336 35216
rect 289176 34416 289228 34468
rect 437480 34416 437532 34468
rect 53840 33804 53892 33856
rect 267096 33804 267148 33856
rect 60832 33736 60884 33788
rect 301596 33736 301648 33788
rect 288440 33124 288492 33176
rect 289176 33124 289228 33176
rect 3516 33056 3568 33108
rect 47584 33056 47636 33108
rect 184204 33056 184256 33108
rect 313924 33056 313976 33108
rect 327724 33056 327776 33108
rect 425060 33056 425112 33108
rect 99380 32444 99432 32496
rect 265624 32444 265676 32496
rect 291844 32444 291896 32496
rect 293960 32444 294012 32496
rect 360844 32444 360896 32496
rect 103520 32376 103572 32428
rect 294696 32376 294748 32428
rect 313280 32036 313332 32088
rect 313924 32036 313976 32088
rect 327080 31764 327132 31816
rect 327724 31764 327776 31816
rect 238024 31152 238076 31204
rect 284392 31152 284444 31204
rect 100760 31084 100812 31136
rect 302976 31084 303028 31136
rect 19340 31016 19392 31068
rect 271236 31016 271288 31068
rect 284392 31016 284444 31068
rect 438860 31016 438912 31068
rect 175924 30268 175976 30320
rect 241520 30268 241572 30320
rect 242164 30268 242216 30320
rect 277400 30268 277452 30320
rect 278044 30268 278096 30320
rect 441620 30268 441672 30320
rect 82820 29656 82872 29708
rect 282368 29656 282420 29708
rect 95240 29588 95292 29640
rect 295984 29588 296036 29640
rect 246304 28364 246356 28416
rect 274640 28364 274692 28416
rect 44272 28296 44324 28348
rect 272524 28296 272576 28348
rect 443000 28296 443052 28348
rect 59268 28228 59320 28280
rect 298836 28228 298888 28280
rect 188344 27548 188396 27600
rect 329840 27548 329892 27600
rect 330484 27548 330536 27600
rect 39856 27004 39908 27056
rect 128360 27004 128412 27056
rect 118792 26936 118844 26988
rect 276756 26936 276808 26988
rect 276940 26936 276992 26988
rect 444380 26936 444432 26988
rect 92480 26868 92532 26920
rect 283564 26868 283616 26920
rect 271144 26188 271196 26240
rect 276940 26188 276992 26240
rect 204904 25576 204956 25628
rect 267740 25576 267792 25628
rect 445852 25576 445904 25628
rect 77392 25508 77444 25560
rect 276664 25508 276716 25560
rect 81440 24216 81492 24268
rect 282276 24216 282328 24268
rect 57980 24148 58032 24200
rect 264244 24148 264296 24200
rect 264336 24148 264388 24200
rect 445944 24148 445996 24200
rect 52552 24080 52604 24132
rect 304264 24080 304316 24132
rect 244924 22924 244976 22976
rect 262312 22924 262364 22976
rect 447140 22924 447192 22976
rect 111800 22856 111852 22908
rect 302884 22856 302936 22908
rect 46940 22788 46992 22840
rect 262864 22788 262916 22840
rect 63500 22720 63552 22772
rect 289084 22720 289136 22772
rect 253204 22040 253256 22092
rect 449900 22040 449952 22092
rect 252560 21564 252612 21616
rect 253204 21564 253256 21616
rect 13820 21428 13872 21480
rect 254584 21428 254636 21480
rect 12440 21360 12492 21412
rect 267004 21360 267056 21412
rect 3424 20612 3476 20664
rect 11704 20612 11756 20664
rect 507768 20612 507820 20664
rect 579988 20612 580040 20664
rect 250536 20000 250588 20052
rect 451280 20000 451332 20052
rect 49700 19932 49752 19984
rect 294604 19932 294656 19984
rect 298836 19252 298888 19304
rect 359556 19252 359608 19304
rect 75920 18708 75972 18760
rect 269764 18708 269816 18760
rect 246304 18640 246356 18692
rect 452660 18640 452712 18692
rect 24860 18572 24912 18624
rect 251824 18572 251876 18624
rect 298100 18028 298152 18080
rect 298836 18028 298888 18080
rect 215944 17280 215996 17332
rect 242992 17280 243044 17332
rect 454132 17280 454184 17332
rect 26240 17212 26292 17264
rect 258724 17212 258776 17264
rect 89168 15988 89220 16040
rect 284944 15988 284996 16040
rect 36728 15920 36780 15972
rect 298744 15920 298796 15972
rect 11888 15852 11940 15904
rect 275284 15852 275336 15904
rect 282276 15852 282328 15904
rect 454040 15852 454092 15904
rect 164424 14492 164476 14544
rect 417424 14492 417476 14544
rect 17040 14424 17092 14476
rect 305644 14424 305696 14476
rect 314660 13744 314712 13796
rect 315304 13744 315356 13796
rect 467840 13744 467892 13796
rect 213184 13132 213236 13184
rect 245200 13132 245252 13184
rect 340144 13132 340196 13184
rect 48504 13064 48556 13116
rect 301504 13064 301556 13116
rect 64788 12384 64840 12436
rect 264152 12384 264204 12436
rect 249064 12316 249116 12368
rect 358084 12316 358136 12368
rect 248420 11908 248472 11960
rect 249064 11908 249116 11960
rect 242900 11772 242952 11824
rect 244096 11772 244148 11824
rect 181444 11704 181496 11756
rect 283104 11704 283156 11756
rect 478880 11704 478932 11756
rect 238024 10412 238076 10464
rect 251272 10412 251324 10464
rect 198004 10344 198056 10396
rect 258264 10344 258316 10396
rect 486424 10344 486476 10396
rect 56048 10276 56100 10328
rect 287796 10276 287848 10328
rect 308404 9596 308456 9648
rect 309048 9596 309100 9648
rect 331588 9596 331640 9648
rect 423680 9596 423732 9648
rect 356704 9528 356756 9580
rect 91560 8984 91612 9036
rect 307024 8984 307076 9036
rect 3332 8916 3384 8968
rect 29644 8916 29696 8968
rect 65524 8916 65576 8968
rect 283656 8916 283708 8968
rect 332600 8848 332652 8900
rect 333888 8848 333940 8900
rect 232504 7692 232556 7744
rect 39948 7624 40000 7676
rect 301504 7624 301556 7676
rect 8760 7556 8812 7608
rect 286416 7556 286468 7608
rect 306748 7556 306800 7608
rect 431960 7556 432012 7608
rect 281908 6808 281960 6860
rect 439504 6808 439556 6860
rect 543004 6808 543056 6860
rect 580172 6808 580224 6860
rect 301504 6740 301556 6792
rect 363604 6740 363656 6792
rect 308496 6672 308548 6724
rect 309784 6672 309836 6724
rect 34336 6264 34388 6316
rect 132960 6264 133012 6316
rect 108120 6196 108172 6248
rect 250444 6196 250496 6248
rect 28908 6128 28960 6180
rect 287704 6128 287756 6180
rect 257068 5448 257120 5500
rect 257344 5448 257396 5500
rect 448520 5448 448572 5500
rect 180064 4768 180116 4820
rect 239220 4768 239272 4820
rect 177396 4088 177448 4140
rect 249984 4088 250036 4140
rect 250536 4088 250588 4140
rect 332692 4088 332744 4140
rect 333244 4088 333296 4140
rect 346952 4088 347004 4140
rect 352564 4088 352616 4140
rect 191104 4020 191156 4072
rect 246396 4020 246448 4072
rect 239220 3952 239272 4004
rect 282276 3952 282328 4004
rect 109316 3612 109368 3664
rect 173164 3612 173216 3664
rect 66720 3544 66772 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 60740 3476 60792 3528
rect 61660 3476 61712 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 77300 3544 77352 3596
rect 78220 3544 78272 3596
rect 93860 3544 93912 3596
rect 94780 3544 94832 3596
rect 103336 3544 103388 3596
rect 187056 3544 187108 3596
rect 251272 3544 251324 3596
rect 252652 3544 252704 3596
rect 170404 3476 170456 3528
rect 251180 3476 251232 3528
rect 252376 3476 252428 3528
rect 276020 3476 276072 3528
rect 276848 3476 276900 3528
rect 316684 3476 316736 3528
rect 317328 3476 317380 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 329196 3476 329248 3528
rect 331312 3476 331364 3528
rect 349804 3476 349856 3528
rect 350448 3476 350500 3528
rect 6460 3408 6512 3460
rect 17224 3408 17276 3460
rect 24216 3408 24268 3460
rect 178684 3408 178736 3460
rect 324412 3408 324464 3460
rect 345756 3408 345808 3460
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 133144 3340 133196 3392
rect 136456 3340 136508 3392
rect 260656 3272 260708 3324
rect 262312 3272 262364 3324
rect 235816 3068 235868 3120
rect 238024 3068 238076 3120
rect 292580 3068 292632 3120
rect 295432 3068 295484 3120
rect 171968 3000 172020 3052
rect 177304 3000 177356 3052
rect 35992 2048 36044 2100
rect 297364 2048 297416 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3436 588606 3464 619103
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 588600 3476 588606
rect 3424 588542 3476 588548
rect 3424 582480 3476 582486
rect 3424 582422 3476 582428
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 553897 3464 582422
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 4816 539578 4844 632062
rect 6932 598262 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 697678 24348 703520
rect 24308 697672 24360 697678
rect 24308 697614 24360 697620
rect 15844 683188 15896 683194
rect 15844 683130 15896 683136
rect 6920 598256 6972 598262
rect 6920 598198 6972 598204
rect 15856 596834 15884 683130
rect 35164 605872 35216 605878
rect 35164 605814 35216 605820
rect 15844 596828 15896 596834
rect 15844 596770 15896 596776
rect 15844 579692 15896 579698
rect 15844 579634 15896 579640
rect 4804 539572 4856 539578
rect 4804 539514 4856 539520
rect 15856 538218 15884 579634
rect 34428 575544 34480 575550
rect 34428 575486 34480 575492
rect 25504 565888 25556 565894
rect 25504 565830 25556 565836
rect 25516 544406 25544 565830
rect 25504 544400 25556 544406
rect 25504 544342 25556 544348
rect 15844 538212 15896 538218
rect 15844 538154 15896 538160
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 34244 525836 34296 525842
rect 34244 525778 34296 525784
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 4804 514820 4856 514826
rect 2780 514762 2832 514768
rect 4804 514762 4856 514768
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3528 494766 3556 501735
rect 4816 496126 4844 514762
rect 4804 496120 4856 496126
rect 4804 496062 4856 496068
rect 3516 494760 3568 494766
rect 3516 494702 3568 494708
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 11704 474768 11756 474774
rect 11704 474710 11756 474716
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 4804 462596 4856 462602
rect 2780 462538 2832 462544
rect 4804 462538 4856 462544
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3436 435985 3464 449511
rect 4816 438190 4844 462538
rect 11716 438938 11744 474710
rect 33048 449948 33100 449954
rect 33048 449890 33100 449896
rect 11704 438932 11756 438938
rect 11704 438874 11756 438880
rect 4804 438184 4856 438190
rect 4804 438126 4856 438132
rect 3422 435976 3478 435985
rect 3422 435911 3478 435920
rect 3424 429888 3476 429894
rect 3424 429830 3476 429836
rect 3436 410553 3464 429830
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 4804 388068 4856 388074
rect 4804 388010 4856 388016
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 357882 3464 358391
rect 3424 357876 3476 357882
rect 3424 357818 3476 357824
rect 4816 346322 4844 388010
rect 7564 357876 7616 357882
rect 7564 357818 7616 357824
rect 7576 346390 7604 357818
rect 33060 352578 33088 449890
rect 34256 442270 34284 525778
rect 34336 476128 34388 476134
rect 34336 476070 34388 476076
rect 34244 442264 34296 442270
rect 34244 442206 34296 442212
rect 34256 431954 34284 442206
rect 34164 431926 34284 431954
rect 33048 352572 33100 352578
rect 33048 352514 33100 352520
rect 15844 351960 15896 351966
rect 15844 351902 15896 351908
rect 7564 346384 7616 346390
rect 7564 346326 7616 346332
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 4804 331288 4856 331294
rect 4804 331230 4856 331236
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 319122 3464 319223
rect 3424 319116 3476 319122
rect 3424 319058 3476 319064
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 4816 293214 4844 331230
rect 7564 319116 7616 319122
rect 7564 319058 7616 319064
rect 7576 314634 7604 319058
rect 7564 314628 7616 314634
rect 7564 314570 7616 314576
rect 15856 306338 15884 351902
rect 34164 342242 34192 431926
rect 34244 386504 34296 386510
rect 34244 386446 34296 386452
rect 34152 342236 34204 342242
rect 34152 342178 34204 342184
rect 15844 306332 15896 306338
rect 15844 306274 15896 306280
rect 11704 299532 11756 299538
rect 11704 299474 11756 299480
rect 2780 293208 2832 293214
rect 2778 293176 2780 293185
rect 4804 293208 4856 293214
rect 2832 293176 2834 293185
rect 4804 293150 4856 293156
rect 2778 293111 2834 293120
rect 5448 292664 5500 292670
rect 5448 292606 5500 292612
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 248414 3464 254079
rect 3436 248386 3556 248414
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3528 240106 3556 248386
rect 3516 240100 3568 240106
rect 3516 240042 3568 240048
rect 1306 217288 1362 217297
rect 1306 217223 1362 217232
rect 1320 75886 1348 217223
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111036 3476 111042
rect 3424 110978 3476 110984
rect 3436 110673 3464 110978
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 2780 76560 2832 76566
rect 2780 76502 2832 76508
rect 20 75880 72 75886
rect 20 75822 72 75828
rect 1308 75880 1360 75886
rect 1308 75822 1360 75828
rect 32 16574 60 75822
rect 2688 67584 2740 67590
rect 2688 67526 2740 67532
rect 32 16546 152 16574
rect 124 354 152 16546
rect 2700 3534 2728 67526
rect 2792 6914 2820 76502
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 5460 67590 5488 292606
rect 7564 210452 7616 210458
rect 7564 210394 7616 210400
rect 7576 111042 7604 210394
rect 7564 111036 7616 111042
rect 7564 110978 7616 110984
rect 5448 67584 5500 67590
rect 5448 67526 5500 67532
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 6920 57248 6972 57254
rect 6920 57190 6972 57196
rect 4160 53168 4212 53174
rect 4160 53110 4212 53116
rect 2872 46232 2924 46238
rect 2872 46174 2924 46180
rect 2884 16574 2912 46174
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 53110
rect 6932 16574 6960 57190
rect 11060 54528 11112 54534
rect 11060 54470 11112 54476
rect 9680 49020 9732 49026
rect 9680 48962 9732 48968
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 2792 6886 2912 6914
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1688 480 1716 3470
rect 2884 480 2912 6886
rect 3344 6497 3372 8910
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8760 7608 8812 7614
rect 8760 7550 8812 7556
rect 8772 480 8800 7550
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 48962
rect 11072 16574 11100 54470
rect 11716 20670 11744 299474
rect 25504 297424 25556 297430
rect 25504 297366 25556 297372
rect 15844 290488 15896 290494
rect 15844 290430 15896 290436
rect 14464 257372 14516 257378
rect 14464 257314 14516 257320
rect 14476 137970 14504 257314
rect 15856 150414 15884 290430
rect 21364 264240 21416 264246
rect 21364 264182 21416 264188
rect 17224 229764 17276 229770
rect 17224 229706 17276 229712
rect 15844 150408 15896 150414
rect 15844 150350 15896 150356
rect 14464 137964 14516 137970
rect 14464 137906 14516 137912
rect 17236 97986 17264 229706
rect 21376 215286 21404 264182
rect 21364 215280 21416 215286
rect 21364 215222 21416 215228
rect 22744 182844 22796 182850
rect 22744 182786 22796 182792
rect 17224 97980 17276 97986
rect 17224 97922 17276 97928
rect 20720 68332 20772 68338
rect 20720 68274 20772 68280
rect 17960 61396 18012 61402
rect 17960 61338 18012 61344
rect 15200 60036 15252 60042
rect 15200 59978 15252 59984
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 11704 20664 11756 20670
rect 11704 20606 11756 20612
rect 12452 16574 12480 21354
rect 13832 16574 13860 21422
rect 15212 16574 15240 59978
rect 17222 18592 17278 18601
rect 17222 18527 17278 18536
rect 11072 16546 11192 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 11164 480 11192 16546
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 15846
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17052 480 17080 14418
rect 17236 3466 17264 18527
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 61338
rect 19340 31068 19392 31074
rect 19340 31010 19392 31016
rect 19352 16574 19380 31010
rect 20732 16574 20760 68274
rect 22756 45558 22784 182786
rect 25516 59362 25544 297366
rect 33784 294024 33836 294030
rect 33784 293966 33836 293972
rect 29644 279472 29696 279478
rect 29644 279414 29696 279420
rect 25504 59356 25556 59362
rect 25504 59298 25556 59304
rect 22744 45552 22796 45558
rect 22744 45494 22796 45500
rect 29000 36644 29052 36650
rect 29000 36586 29052 36592
rect 22100 35216 22152 35222
rect 22100 35158 22152 35164
rect 22112 16574 22140 35158
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24872 16574 24900 18566
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 19444 480 19472 16546
rect 20166 10296 20222 10305
rect 20166 10231 20222 10240
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 10231
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 17206
rect 29012 6914 29040 36586
rect 29656 8974 29684 279414
rect 32404 253224 32456 253230
rect 32404 253166 32456 253172
rect 32416 85542 32444 253166
rect 33796 164218 33824 293966
rect 34256 258058 34284 386446
rect 34244 258052 34296 258058
rect 34244 257994 34296 258000
rect 34256 257378 34284 257994
rect 34244 257372 34296 257378
rect 34244 257314 34296 257320
rect 33784 164212 33836 164218
rect 33784 164154 33836 164160
rect 32404 85536 32456 85542
rect 32404 85478 32456 85484
rect 31760 65544 31812 65550
rect 31760 65486 31812 65492
rect 31772 16574 31800 65486
rect 33138 42120 33194 42129
rect 33138 42055 33194 42064
rect 33152 16574 33180 42055
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 30838 11656 30894 11665
rect 30838 11591 30894 11600
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29012 6886 30144 6914
rect 28908 6180 28960 6186
rect 28908 6122 28960 6128
rect 27710 4856 27766 4865
rect 27710 4791 27766 4800
rect 27724 480 27752 4791
rect 28920 480 28948 6122
rect 30116 480 30144 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 11591
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 34348 6322 34376 476070
rect 34440 39506 34468 575486
rect 35176 536790 35204 605814
rect 40052 592074 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 77944 703316 77996 703322
rect 77944 703258 77996 703264
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 76564 703044 76616 703050
rect 76564 702986 76616 702992
rect 68928 702500 68980 702506
rect 68928 702442 68980 702448
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 57888 697604 57940 697610
rect 57888 697546 57940 697552
rect 54484 670744 54536 670750
rect 54484 670686 54536 670692
rect 53104 598256 53156 598262
rect 53104 598198 53156 598204
rect 53116 597582 53144 598198
rect 53104 597576 53156 597582
rect 53104 597518 53156 597524
rect 50988 596828 51040 596834
rect 50988 596770 51040 596776
rect 51000 596222 51028 596770
rect 50988 596216 51040 596222
rect 50988 596158 51040 596164
rect 40040 592068 40092 592074
rect 40040 592010 40092 592016
rect 48228 592068 48280 592074
rect 48228 592010 48280 592016
rect 48044 586628 48096 586634
rect 48044 586570 48096 586576
rect 42616 586560 42668 586566
rect 42616 586502 42668 586508
rect 41236 585200 41288 585206
rect 41236 585142 41288 585148
rect 39764 581256 39816 581262
rect 39764 581198 39816 581204
rect 37004 581052 37056 581058
rect 37004 580994 37056 581000
rect 35716 549296 35768 549302
rect 35716 549238 35768 549244
rect 35164 536784 35216 536790
rect 35164 536726 35216 536732
rect 35624 475380 35676 475386
rect 35624 475322 35676 475328
rect 35636 379506 35664 475322
rect 35728 451246 35756 549238
rect 35808 545148 35860 545154
rect 35808 545090 35860 545096
rect 35716 451240 35768 451246
rect 35716 451182 35768 451188
rect 35728 449954 35756 451182
rect 35716 449948 35768 449954
rect 35716 449890 35768 449896
rect 35820 445738 35848 545090
rect 37016 483682 37044 580994
rect 37096 556232 37148 556238
rect 37096 556174 37148 556180
rect 37004 483676 37056 483682
rect 37004 483618 37056 483624
rect 36912 482316 36964 482322
rect 36912 482258 36964 482264
rect 35808 445732 35860 445738
rect 35808 445674 35860 445680
rect 36924 392630 36952 482258
rect 37108 460934 37136 556174
rect 37188 554804 37240 554810
rect 37188 554746 37240 554752
rect 37016 460906 37136 460934
rect 37016 457502 37044 460906
rect 37004 457496 37056 457502
rect 37004 457438 37056 457444
rect 36912 392624 36964 392630
rect 36912 392566 36964 392572
rect 35716 385144 35768 385150
rect 35716 385086 35768 385092
rect 35624 379500 35676 379506
rect 35624 379442 35676 379448
rect 35728 249082 35756 385086
rect 37016 361554 37044 457438
rect 37200 455394 37228 554746
rect 38568 550656 38620 550662
rect 38568 550598 38620 550604
rect 38476 497480 38528 497486
rect 38476 497422 38528 497428
rect 37188 455388 37240 455394
rect 37188 455330 37240 455336
rect 38488 440910 38516 497422
rect 38580 451178 38608 550598
rect 39672 526448 39724 526454
rect 39672 526390 39724 526396
rect 38568 451172 38620 451178
rect 38568 451114 38620 451120
rect 38476 440904 38528 440910
rect 38476 440846 38528 440852
rect 38488 440298 38516 440846
rect 37096 440292 37148 440298
rect 37096 440234 37148 440240
rect 38476 440292 38528 440298
rect 38476 440234 38528 440240
rect 37004 361548 37056 361554
rect 37004 361490 37056 361496
rect 35808 349172 35860 349178
rect 35808 349114 35860 349120
rect 35716 249076 35768 249082
rect 35716 249018 35768 249024
rect 35820 52358 35848 349114
rect 37108 339658 37136 440234
rect 38476 389836 38528 389842
rect 38476 389778 38528 389784
rect 37188 378820 37240 378826
rect 37188 378762 37240 378768
rect 37096 339652 37148 339658
rect 37096 339594 37148 339600
rect 37096 331900 37148 331906
rect 37096 331842 37148 331848
rect 37108 331294 37136 331842
rect 37096 331288 37148 331294
rect 37096 331230 37148 331236
rect 37108 244254 37136 331230
rect 37096 244248 37148 244254
rect 37096 244190 37148 244196
rect 37200 240106 37228 378762
rect 38488 306374 38516 389778
rect 38580 386374 38608 451114
rect 39684 436762 39712 526390
rect 39776 483002 39804 581198
rect 41144 564528 41196 564534
rect 41144 564470 41196 564476
rect 39856 547936 39908 547942
rect 39856 547878 39908 547884
rect 39764 482996 39816 483002
rect 39764 482938 39816 482944
rect 39764 458176 39816 458182
rect 39764 458118 39816 458124
rect 39672 436756 39724 436762
rect 39672 436698 39724 436704
rect 38568 386368 38620 386374
rect 38568 386310 38620 386316
rect 39776 359514 39804 458118
rect 39868 448526 39896 547878
rect 40960 529236 41012 529242
rect 40960 529178 41012 529184
rect 39948 492108 40000 492114
rect 39948 492050 40000 492056
rect 39856 448520 39908 448526
rect 39856 448462 39908 448468
rect 39960 389910 39988 492050
rect 40972 434722 41000 529178
rect 41156 470594 41184 564470
rect 41248 491366 41276 585142
rect 41328 569968 41380 569974
rect 41328 569910 41380 569916
rect 41236 491360 41288 491366
rect 41236 491302 41288 491308
rect 41064 470566 41184 470594
rect 41064 465730 41092 470566
rect 41052 465724 41104 465730
rect 41052 465666 41104 465672
rect 40960 434716 41012 434722
rect 40960 434658 41012 434664
rect 39948 389904 40000 389910
rect 39948 389846 40000 389852
rect 39948 387932 40000 387938
rect 39948 387874 40000 387880
rect 39856 382288 39908 382294
rect 39856 382230 39908 382236
rect 39764 359508 39816 359514
rect 39764 359450 39816 359456
rect 38488 306346 38608 306374
rect 38580 291174 38608 306346
rect 38568 291168 38620 291174
rect 38568 291110 38620 291116
rect 38580 290494 38608 291110
rect 38568 290488 38620 290494
rect 38568 290430 38620 290436
rect 38568 284368 38620 284374
rect 38568 284310 38620 284316
rect 37188 240100 37240 240106
rect 37188 240042 37240 240048
rect 37200 238882 37228 240042
rect 37188 238876 37240 238882
rect 37188 238818 37240 238824
rect 38580 230450 38608 284310
rect 39776 235754 39804 359450
rect 39764 235748 39816 235754
rect 39764 235690 39816 235696
rect 38568 230444 38620 230450
rect 38568 230386 38620 230392
rect 37280 53100 37332 53106
rect 37280 53042 37332 53048
rect 35808 52352 35860 52358
rect 35808 52294 35860 52300
rect 34520 47660 34572 47666
rect 34520 47602 34572 47608
rect 34428 39500 34480 39506
rect 34428 39442 34480 39448
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 47602
rect 37292 16574 37320 53042
rect 39868 27062 39896 382230
rect 39856 27056 39908 27062
rect 39856 26998 39908 27004
rect 37292 16546 38424 16574
rect 36728 15972 36780 15978
rect 36728 15914 36780 15920
rect 35992 2100 36044 2106
rect 35992 2042 36044 2048
rect 36004 480 36032 2042
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 15914
rect 38396 480 38424 16546
rect 39118 14512 39174 14521
rect 39118 14447 39174 14456
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 14447
rect 39960 7682 39988 387874
rect 40972 339425 41000 434658
rect 41064 371210 41092 465666
rect 41144 396092 41196 396098
rect 41144 396034 41196 396040
rect 41052 371204 41104 371210
rect 41052 371146 41104 371152
rect 40958 339416 41014 339425
rect 40958 339351 41014 339360
rect 41156 282878 41184 396034
rect 41248 393310 41276 491302
rect 41340 470558 41368 569910
rect 42628 490006 42656 586502
rect 46756 585268 46808 585274
rect 46756 585210 46808 585216
rect 45468 584044 45520 584050
rect 45468 583986 45520 583992
rect 43812 581120 43864 581126
rect 43812 581062 43864 581068
rect 42708 558952 42760 558958
rect 42708 558894 42760 558900
rect 42616 490000 42668 490006
rect 42616 489942 42668 489948
rect 42628 489914 42656 489942
rect 42536 489886 42656 489914
rect 41328 470552 41380 470558
rect 41328 470494 41380 470500
rect 42536 403617 42564 489886
rect 42616 473408 42668 473414
rect 42616 473350 42668 473356
rect 42522 403608 42578 403617
rect 42522 403543 42578 403552
rect 41236 393304 41288 393310
rect 41236 393246 41288 393252
rect 42628 379438 42656 473350
rect 42720 460222 42748 558894
rect 43720 556300 43772 556306
rect 43720 556242 43772 556248
rect 42708 460216 42760 460222
rect 42708 460158 42760 460164
rect 43732 458182 43760 556242
rect 43824 489870 43852 581062
rect 45376 537668 45428 537674
rect 45376 537610 45428 537616
rect 44088 537600 44140 537606
rect 44088 537542 44140 537548
rect 43904 494828 43956 494834
rect 43904 494770 43956 494776
rect 43812 489864 43864 489870
rect 43812 489806 43864 489812
rect 43720 458176 43772 458182
rect 43720 458118 43772 458124
rect 43720 439068 43772 439074
rect 43720 439010 43772 439016
rect 42708 432608 42760 432614
rect 42708 432550 42760 432556
rect 42616 379432 42668 379438
rect 42616 379374 42668 379380
rect 41236 364404 41288 364410
rect 41236 364346 41288 364352
rect 41144 282872 41196 282878
rect 41144 282814 41196 282820
rect 41248 241466 41276 364346
rect 42616 356108 42668 356114
rect 42616 356050 42668 356056
rect 41328 343664 41380 343670
rect 41328 343606 41380 343612
rect 40868 241460 40920 241466
rect 40868 241402 40920 241408
rect 41236 241460 41288 241466
rect 41236 241402 41288 241408
rect 40880 240786 40908 241402
rect 40868 240780 40920 240786
rect 40868 240722 40920 240728
rect 41340 71670 41368 343606
rect 42628 280158 42656 356050
rect 42720 335170 42748 432550
rect 43732 337958 43760 439010
rect 43916 399498 43944 494770
rect 43996 458924 44048 458930
rect 43996 458866 44048 458872
rect 43904 399492 43956 399498
rect 43904 399434 43956 399440
rect 43812 396840 43864 396846
rect 43812 396782 43864 396788
rect 43824 340270 43852 396782
rect 44008 363662 44036 458866
rect 44100 437238 44128 537542
rect 45284 489932 45336 489938
rect 45284 489874 45336 489880
rect 44088 437232 44140 437238
rect 44088 437174 44140 437180
rect 45296 402286 45324 489874
rect 45388 439074 45416 537610
rect 45480 492114 45508 583986
rect 46572 534744 46624 534750
rect 46572 534686 46624 534692
rect 45468 492108 45520 492114
rect 45468 492050 45520 492056
rect 45468 458856 45520 458862
rect 45468 458798 45520 458804
rect 45376 439068 45428 439074
rect 45376 439010 45428 439016
rect 45284 402280 45336 402286
rect 45284 402222 45336 402228
rect 45284 395412 45336 395418
rect 45284 395354 45336 395360
rect 43996 363656 44048 363662
rect 43996 363598 44048 363604
rect 43904 345092 43956 345098
rect 43904 345034 43956 345040
rect 43812 340264 43864 340270
rect 43812 340206 43864 340212
rect 43720 337952 43772 337958
rect 43720 337894 43772 337900
rect 42708 335164 42760 335170
rect 42708 335106 42760 335112
rect 42708 289876 42760 289882
rect 42708 289818 42760 289824
rect 41420 280152 41472 280158
rect 41420 280094 41472 280100
rect 42616 280152 42668 280158
rect 42616 280094 42668 280100
rect 41432 279478 41460 280094
rect 41420 279472 41472 279478
rect 41420 279414 41472 279420
rect 42720 225690 42748 289818
rect 43812 273284 43864 273290
rect 43812 273226 43864 273232
rect 42708 225684 42760 225690
rect 42708 225626 42760 225632
rect 43824 210526 43852 273226
rect 43916 268462 43944 345034
rect 43904 268456 43956 268462
rect 43904 268398 43956 268404
rect 44008 264246 44036 363598
rect 45296 333946 45324 395354
rect 45376 385892 45428 385898
rect 45376 385834 45428 385840
rect 45284 333940 45336 333946
rect 45284 333882 45336 333888
rect 44088 293276 44140 293282
rect 44088 293218 44140 293224
rect 43996 264240 44048 264246
rect 43996 264182 44048 264188
rect 43812 210520 43864 210526
rect 43812 210462 43864 210468
rect 44100 72554 44128 293218
rect 45388 267714 45416 385834
rect 45480 361486 45508 458798
rect 46584 437374 46612 534686
rect 46768 533390 46796 585210
rect 47952 583840 48004 583846
rect 47952 583782 48004 583788
rect 46848 542428 46900 542434
rect 46848 542370 46900 542376
rect 46756 533384 46808 533390
rect 46756 533326 46808 533332
rect 46664 529304 46716 529310
rect 46664 529246 46716 529252
rect 46676 442377 46704 529246
rect 46860 443698 46888 542370
rect 47860 494556 47912 494562
rect 47860 494498 47912 494504
rect 47872 494086 47900 494498
rect 47860 494080 47912 494086
rect 47860 494022 47912 494028
rect 46848 443692 46900 443698
rect 46848 443634 46900 443640
rect 46662 442368 46718 442377
rect 46662 442303 46718 442312
rect 46572 437368 46624 437374
rect 46572 437310 46624 437316
rect 46756 436756 46808 436762
rect 46756 436698 46808 436704
rect 46664 387116 46716 387122
rect 46664 387058 46716 387064
rect 45468 361480 45520 361486
rect 45468 361422 45520 361428
rect 46572 349240 46624 349246
rect 46572 349182 46624 349188
rect 45468 337544 45520 337550
rect 45468 337486 45520 337492
rect 45376 267708 45428 267714
rect 45376 267650 45428 267656
rect 44088 72548 44140 72554
rect 44088 72490 44140 72496
rect 41328 71664 41380 71670
rect 41328 71606 41380 71612
rect 40040 69692 40092 69698
rect 40040 69634 40092 69640
rect 40052 16574 40080 69634
rect 41420 50380 41472 50386
rect 41420 50322 41472 50328
rect 41432 16574 41460 50322
rect 45480 46306 45508 337486
rect 46584 234598 46612 349182
rect 46676 335238 46704 387058
rect 46768 336462 46796 436698
rect 46860 344350 46888 443634
rect 47872 404977 47900 494022
rect 47964 492726 47992 583782
rect 48056 494562 48084 586570
rect 48136 534880 48188 534886
rect 48136 534822 48188 534828
rect 48044 494556 48096 494562
rect 48044 494498 48096 494504
rect 47952 492720 48004 492726
rect 47952 492662 48004 492668
rect 47964 489914 47992 492662
rect 47964 489886 48084 489914
rect 47858 404968 47914 404977
rect 47858 404903 47914 404912
rect 48056 395350 48084 489886
rect 48148 438734 48176 534822
rect 48240 487830 48268 592010
rect 49608 586696 49660 586702
rect 49608 586638 49660 586644
rect 49424 563100 49476 563106
rect 49424 563042 49476 563048
rect 48228 487824 48280 487830
rect 48228 487766 48280 487772
rect 48136 438728 48188 438734
rect 48136 438670 48188 438676
rect 48044 395344 48096 395350
rect 48044 395286 48096 395292
rect 47860 392148 47912 392154
rect 47860 392090 47912 392096
rect 46848 344344 46900 344350
rect 46848 344286 46900 344292
rect 46756 336456 46808 336462
rect 46756 336398 46808 336404
rect 46664 335232 46716 335238
rect 46664 335174 46716 335180
rect 46756 294092 46808 294098
rect 46756 294034 46808 294040
rect 46572 234592 46624 234598
rect 46572 234534 46624 234540
rect 46768 207738 46796 294034
rect 47872 269074 47900 392090
rect 47952 391332 48004 391338
rect 47952 391274 48004 391280
rect 47964 332586 47992 391274
rect 48044 379568 48096 379574
rect 48044 379510 48096 379516
rect 47952 332580 48004 332586
rect 47952 332522 48004 332528
rect 48056 314634 48084 379510
rect 48148 336530 48176 438670
rect 48240 388482 48268 487766
rect 49436 464370 49464 563042
rect 49516 532160 49568 532166
rect 49516 532102 49568 532108
rect 49424 464364 49476 464370
rect 49424 464306 49476 464312
rect 49436 463690 49464 464306
rect 49424 463684 49476 463690
rect 49424 463626 49476 463632
rect 49528 433294 49556 532102
rect 49620 494834 49648 586638
rect 50804 582548 50856 582554
rect 50804 582490 50856 582496
rect 49608 494828 49660 494834
rect 49608 494770 49660 494776
rect 49608 492040 49660 492046
rect 49608 491982 49660 491988
rect 49516 433288 49568 433294
rect 49516 433230 49568 433236
rect 49528 432614 49556 433230
rect 49516 432608 49568 432614
rect 49516 432550 49568 432556
rect 49516 393984 49568 393990
rect 49516 393926 49568 393932
rect 48964 389292 49016 389298
rect 48964 389234 49016 389240
rect 48228 388476 48280 388482
rect 48228 388418 48280 388424
rect 48976 372570 49004 389234
rect 49332 385756 49384 385762
rect 49332 385698 49384 385704
rect 48964 372564 49016 372570
rect 48964 372506 49016 372512
rect 48136 336524 48188 336530
rect 48136 336466 48188 336472
rect 49344 333810 49372 385698
rect 49424 351960 49476 351966
rect 49424 351902 49476 351908
rect 49332 333804 49384 333810
rect 49332 333746 49384 333752
rect 48136 332648 48188 332654
rect 48136 332590 48188 332596
rect 48044 314628 48096 314634
rect 48044 314570 48096 314576
rect 48056 313954 48084 314570
rect 48044 313948 48096 313954
rect 48044 313890 48096 313896
rect 48044 302320 48096 302326
rect 48044 302262 48096 302268
rect 47860 269068 47912 269074
rect 47860 269010 47912 269016
rect 48056 253910 48084 302262
rect 47676 253904 47728 253910
rect 47676 253846 47728 253852
rect 48044 253904 48096 253910
rect 48044 253846 48096 253852
rect 47688 253230 47716 253846
rect 47676 253224 47728 253230
rect 47676 253166 47728 253172
rect 48148 238678 48176 332590
rect 49436 323746 49464 351902
rect 49528 338094 49556 393926
rect 49620 385898 49648 491982
rect 50816 491298 50844 582490
rect 50896 553444 50948 553450
rect 50896 553386 50948 553392
rect 50804 491292 50856 491298
rect 50804 491234 50856 491240
rect 50804 490612 50856 490618
rect 50804 490554 50856 490560
rect 50344 463684 50396 463690
rect 50344 463626 50396 463632
rect 49608 385892 49660 385898
rect 49608 385834 49660 385840
rect 49620 385082 49648 385834
rect 49608 385076 49660 385082
rect 49608 385018 49660 385024
rect 50356 368558 50384 463626
rect 50816 436082 50844 490554
rect 50908 452606 50936 553386
rect 51000 484362 51028 596158
rect 52368 586764 52420 586770
rect 52368 586706 52420 586712
rect 52184 579692 52236 579698
rect 52184 579634 52236 579640
rect 52092 537532 52144 537538
rect 52092 537474 52144 537480
rect 50988 484356 51040 484362
rect 50988 484298 51040 484304
rect 50896 452600 50948 452606
rect 50896 452542 50948 452548
rect 51724 452600 51776 452606
rect 51724 452542 51776 452548
rect 50988 438864 51040 438870
rect 50988 438806 51040 438812
rect 51000 438190 51028 438806
rect 50988 438184 51040 438190
rect 50988 438126 51040 438132
rect 50804 436076 50856 436082
rect 50804 436018 50856 436024
rect 51000 431954 51028 438126
rect 50908 431926 51028 431954
rect 50804 388612 50856 388618
rect 50804 388554 50856 388560
rect 50344 368552 50396 368558
rect 50344 368494 50396 368500
rect 49608 352640 49660 352646
rect 49608 352582 49660 352588
rect 49620 351966 49648 352582
rect 49608 351960 49660 351966
rect 49608 351902 49660 351908
rect 49516 338088 49568 338094
rect 49516 338030 49568 338036
rect 49608 336728 49660 336734
rect 49608 336670 49660 336676
rect 49424 323740 49476 323746
rect 49424 323682 49476 323688
rect 49516 320884 49568 320890
rect 49516 320826 49568 320832
rect 49424 287088 49476 287094
rect 49424 287030 49476 287036
rect 48228 269068 48280 269074
rect 48228 269010 48280 269016
rect 48240 268394 48268 269010
rect 48228 268388 48280 268394
rect 48228 268330 48280 268336
rect 48136 238672 48188 238678
rect 48136 238614 48188 238620
rect 48240 234530 48268 268330
rect 48228 234524 48280 234530
rect 48228 234466 48280 234472
rect 48240 234122 48268 234466
rect 47584 234116 47636 234122
rect 47584 234058 47636 234064
rect 48228 234116 48280 234122
rect 48228 234058 48280 234064
rect 46756 207732 46808 207738
rect 46756 207674 46808 207680
rect 45560 77988 45612 77994
rect 45560 77930 45612 77936
rect 45468 46300 45520 46306
rect 45468 46242 45520 46248
rect 44180 36576 44232 36582
rect 44180 36518 44232 36524
rect 42798 17232 42854 17241
rect 42798 17167 42854 17176
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39948 7676 40000 7682
rect 39948 7618 40000 7624
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 17167
rect 44192 6914 44220 36518
rect 44272 28348 44324 28354
rect 44272 28290 44324 28296
rect 44284 16574 44312 28290
rect 45572 16574 45600 77930
rect 47596 33114 47624 234058
rect 49436 221542 49464 287030
rect 49528 244186 49556 320826
rect 49516 244180 49568 244186
rect 49516 244122 49568 244128
rect 49620 237250 49648 336670
rect 50712 334008 50764 334014
rect 50712 333950 50764 333956
rect 50344 266416 50396 266422
rect 50344 266358 50396 266364
rect 49608 237244 49660 237250
rect 49608 237186 49660 237192
rect 50356 234462 50384 266358
rect 50724 255270 50752 333950
rect 50816 297566 50844 388554
rect 50908 337890 50936 431926
rect 50988 397520 51040 397526
rect 50988 397462 51040 397468
rect 50896 337884 50948 337890
rect 50896 337826 50948 337832
rect 50804 297560 50856 297566
rect 50804 297502 50856 297508
rect 50896 280220 50948 280226
rect 50896 280162 50948 280168
rect 50712 255264 50764 255270
rect 50712 255206 50764 255212
rect 50344 234456 50396 234462
rect 50344 234398 50396 234404
rect 49424 221536 49476 221542
rect 49424 221478 49476 221484
rect 50908 186998 50936 280162
rect 51000 238746 51028 397462
rect 51736 396001 51764 452542
rect 52104 437306 52132 537474
rect 52196 481642 52224 579634
rect 52276 548004 52328 548010
rect 52276 547946 52328 547952
rect 52184 481636 52236 481642
rect 52184 481578 52236 481584
rect 52184 472660 52236 472666
rect 52184 472602 52236 472608
rect 52092 437300 52144 437306
rect 52092 437242 52144 437248
rect 51722 395992 51778 396001
rect 51722 395927 51778 395936
rect 52092 385688 52144 385694
rect 52092 385630 52144 385636
rect 52104 335306 52132 385630
rect 52196 376718 52224 472602
rect 52288 447817 52316 547946
rect 52380 532098 52408 586706
rect 52368 532092 52420 532098
rect 52368 532034 52420 532040
rect 53116 492046 53144 597518
rect 53656 585336 53708 585342
rect 53656 585278 53708 585284
rect 53564 534812 53616 534818
rect 53564 534754 53616 534760
rect 53104 492040 53156 492046
rect 53104 491982 53156 491988
rect 53104 484356 53156 484362
rect 53104 484298 53156 484304
rect 52460 460216 52512 460222
rect 52460 460158 52512 460164
rect 52472 459610 52500 460158
rect 52460 459604 52512 459610
rect 52460 459546 52512 459552
rect 52274 447808 52330 447817
rect 52274 447743 52330 447752
rect 53116 394126 53144 484298
rect 53576 438870 53604 534754
rect 53668 488510 53696 585278
rect 53748 552084 53800 552090
rect 53748 552026 53800 552032
rect 53656 488504 53708 488510
rect 53656 488446 53708 488452
rect 53668 487257 53696 488446
rect 53654 487248 53710 487257
rect 53654 487183 53710 487192
rect 53656 459604 53708 459610
rect 53656 459546 53708 459552
rect 53564 438864 53616 438870
rect 53564 438806 53616 438812
rect 53668 398138 53696 459546
rect 53760 452742 53788 552026
rect 54496 538898 54524 670686
rect 57704 588600 57756 588606
rect 57704 588542 57756 588548
rect 57716 587926 57744 588542
rect 57704 587920 57756 587926
rect 57704 587862 57756 587868
rect 55128 584112 55180 584118
rect 55128 584054 55180 584060
rect 55036 556164 55088 556170
rect 55036 556106 55088 556112
rect 54484 538892 54536 538898
rect 54484 538834 54536 538840
rect 54944 532024 54996 532030
rect 54944 531966 54996 531972
rect 54760 493332 54812 493338
rect 54760 493274 54812 493280
rect 53840 473408 53892 473414
rect 53840 473350 53892 473356
rect 53852 473249 53880 473350
rect 53838 473240 53894 473249
rect 53838 473175 53894 473184
rect 53748 452736 53800 452742
rect 53748 452678 53800 452684
rect 53748 439544 53800 439550
rect 53748 439486 53800 439492
rect 53656 398132 53708 398138
rect 53656 398074 53708 398080
rect 53472 396772 53524 396778
rect 53472 396714 53524 396720
rect 53104 394120 53156 394126
rect 53104 394062 53156 394068
rect 52368 394052 52420 394058
rect 52368 393994 52420 394000
rect 52274 390688 52330 390697
rect 52274 390623 52330 390632
rect 52288 390590 52316 390623
rect 52276 390584 52328 390590
rect 52276 390526 52328 390532
rect 52184 376712 52236 376718
rect 52184 376654 52236 376660
rect 52184 355360 52236 355366
rect 52184 355302 52236 355308
rect 52092 335300 52144 335306
rect 52092 335242 52144 335248
rect 52092 330608 52144 330614
rect 52092 330550 52144 330556
rect 52104 287026 52132 330550
rect 52196 300121 52224 355302
rect 52182 300112 52238 300121
rect 52182 300047 52238 300056
rect 52092 287020 52144 287026
rect 52092 286962 52144 286968
rect 52184 285728 52236 285734
rect 52184 285670 52236 285676
rect 52092 271924 52144 271930
rect 52092 271866 52144 271872
rect 50988 238740 51040 238746
rect 50988 238682 51040 238688
rect 52104 227050 52132 271866
rect 52092 227044 52144 227050
rect 52092 226986 52144 226992
rect 52196 206281 52224 285670
rect 52288 255202 52316 390526
rect 52380 335102 52408 393994
rect 53380 338088 53432 338094
rect 53380 338030 53432 338036
rect 53392 337482 53420 338030
rect 53380 337476 53432 337482
rect 53380 337418 53432 337424
rect 52368 335096 52420 335102
rect 52368 335038 52420 335044
rect 52380 334014 52408 335038
rect 52368 334008 52420 334014
rect 52368 333950 52420 333956
rect 52368 299668 52420 299674
rect 52368 299610 52420 299616
rect 52276 255196 52328 255202
rect 52276 255138 52328 255144
rect 52182 206272 52238 206281
rect 52182 206207 52238 206216
rect 50896 186992 50948 186998
rect 50896 186934 50948 186940
rect 52380 71738 52408 299610
rect 53104 292868 53156 292874
rect 53104 292810 53156 292816
rect 53116 189038 53144 292810
rect 53392 245546 53420 337418
rect 53484 333878 53512 396714
rect 53564 391944 53616 391950
rect 53564 391886 53616 391892
rect 53576 358086 53604 391886
rect 53656 388000 53708 388006
rect 53656 387942 53708 387948
rect 53564 358080 53616 358086
rect 53564 358022 53616 358028
rect 53472 333872 53524 333878
rect 53472 333814 53524 333820
rect 53484 332654 53512 333814
rect 53472 332648 53524 332654
rect 53472 332590 53524 332596
rect 53576 271862 53604 358022
rect 53668 298110 53696 387942
rect 53760 337414 53788 439486
rect 54772 389366 54800 493274
rect 54852 480276 54904 480282
rect 54852 480218 54904 480224
rect 54760 389360 54812 389366
rect 54760 389302 54812 389308
rect 54864 388618 54892 480218
rect 54956 437442 54984 531966
rect 55048 455326 55076 556106
rect 55140 487150 55168 584054
rect 56416 583024 56468 583030
rect 56416 582966 56468 582972
rect 56324 557592 56376 557598
rect 56324 557534 56376 557540
rect 56232 491972 56284 491978
rect 56232 491914 56284 491920
rect 55128 487144 55180 487150
rect 55128 487086 55180 487092
rect 55036 455320 55088 455326
rect 55036 455262 55088 455268
rect 56244 437510 56272 491914
rect 56336 468382 56364 557534
rect 56428 538121 56456 582966
rect 57244 578264 57296 578270
rect 57244 578206 57296 578212
rect 56508 561672 56560 561678
rect 56508 561614 56560 561620
rect 56414 538112 56470 538121
rect 56414 538047 56470 538056
rect 56428 537674 56456 538047
rect 56416 537668 56468 537674
rect 56416 537610 56468 537616
rect 56416 529372 56468 529378
rect 56416 529314 56468 529320
rect 56324 468376 56376 468382
rect 56324 468318 56376 468324
rect 56428 441614 56456 529314
rect 56520 463010 56548 561614
rect 57256 480282 57284 578206
rect 57716 538966 57744 587862
rect 57796 560312 57848 560318
rect 57796 560254 57848 560260
rect 57704 538960 57756 538966
rect 57704 538902 57756 538908
rect 57704 537668 57756 537674
rect 57704 537610 57756 537616
rect 57244 480276 57296 480282
rect 57244 480218 57296 480224
rect 56508 463004 56560 463010
rect 56508 462946 56560 462952
rect 56336 441586 56456 441614
rect 56232 437504 56284 437510
rect 56232 437446 56284 437452
rect 54944 437436 54996 437442
rect 54944 437378 54996 437384
rect 55864 437232 55916 437238
rect 55864 437174 55916 437180
rect 54944 399560 54996 399566
rect 54944 399502 54996 399508
rect 54852 388612 54904 388618
rect 54852 388554 54904 388560
rect 54852 387184 54904 387190
rect 54852 387126 54904 387132
rect 54206 355464 54262 355473
rect 54206 355399 54262 355408
rect 54220 355366 54248 355399
rect 54208 355360 54260 355366
rect 54208 355302 54260 355308
rect 54864 339318 54892 387126
rect 54852 339312 54904 339318
rect 54852 339254 54904 339260
rect 54852 338768 54904 338774
rect 54852 338710 54904 338716
rect 53748 337408 53800 337414
rect 53748 337350 53800 337356
rect 53656 298104 53708 298110
rect 53656 298046 53708 298052
rect 53656 274712 53708 274718
rect 53656 274654 53708 274660
rect 53564 271856 53616 271862
rect 53564 271798 53616 271804
rect 53564 256760 53616 256766
rect 53564 256702 53616 256708
rect 53380 245540 53432 245546
rect 53380 245482 53432 245488
rect 53576 216646 53604 256702
rect 53564 216640 53616 216646
rect 53564 216582 53616 216588
rect 53668 214742 53696 274654
rect 54864 266354 54892 338710
rect 54956 336666 54984 399502
rect 55128 391264 55180 391270
rect 55128 391206 55180 391212
rect 55036 368552 55088 368558
rect 55036 368494 55088 368500
rect 54944 336660 54996 336666
rect 54944 336602 54996 336608
rect 54944 326528 54996 326534
rect 54944 326470 54996 326476
rect 54852 266348 54904 266354
rect 54852 266290 54904 266296
rect 53840 264240 53892 264246
rect 53840 264182 53892 264188
rect 53852 263634 53880 264182
rect 53840 263628 53892 263634
rect 53840 263570 53892 263576
rect 54852 263628 54904 263634
rect 54852 263570 54904 263576
rect 54864 231810 54892 263570
rect 54956 245614 54984 326470
rect 55048 304298 55076 368494
rect 55140 338842 55168 391206
rect 55876 339386 55904 437174
rect 56336 434654 56364 441586
rect 56416 438252 56468 438258
rect 56416 438194 56468 438200
rect 56428 437238 56456 438194
rect 56416 437232 56468 437238
rect 56416 437174 56468 437180
rect 56324 434648 56376 434654
rect 56324 434590 56376 434596
rect 56416 399628 56468 399634
rect 56416 399570 56468 399576
rect 56324 389224 56376 389230
rect 56324 389166 56376 389172
rect 56336 367062 56364 389166
rect 56324 367056 56376 367062
rect 56324 366998 56376 367004
rect 56324 363724 56376 363730
rect 56324 363666 56376 363672
rect 55864 339380 55916 339386
rect 55864 339322 55916 339328
rect 55128 338836 55180 338842
rect 55128 338778 55180 338784
rect 55128 337408 55180 337414
rect 55128 337350 55180 337356
rect 55036 304292 55088 304298
rect 55036 304234 55088 304240
rect 55036 294160 55088 294166
rect 55036 294102 55088 294108
rect 54944 245608 54996 245614
rect 54944 245550 54996 245556
rect 54852 231804 54904 231810
rect 54852 231746 54904 231752
rect 53656 214736 53708 214742
rect 53656 214678 53708 214684
rect 55048 202230 55076 294102
rect 55140 237318 55168 337350
rect 56232 297560 56284 297566
rect 56232 297502 56284 297508
rect 56244 280090 56272 297502
rect 56336 297430 56364 363666
rect 56428 336598 56456 399570
rect 56520 390522 56548 462946
rect 57336 455320 57388 455326
rect 57336 455262 57388 455268
rect 57348 454102 57376 455262
rect 57336 454096 57388 454102
rect 57336 454038 57388 454044
rect 57244 438184 57296 438190
rect 57244 438126 57296 438132
rect 57256 437510 57284 438126
rect 57244 437504 57296 437510
rect 57244 437446 57296 437452
rect 56508 390516 56560 390522
rect 56508 390458 56560 390464
rect 56520 389230 56548 390458
rect 56508 389224 56560 389230
rect 56508 389166 56560 389172
rect 56506 387696 56562 387705
rect 56506 387631 56562 387640
rect 56520 386578 56548 387631
rect 56508 386572 56560 386578
rect 56508 386514 56560 386520
rect 56416 336592 56468 336598
rect 56416 336534 56468 336540
rect 56416 331968 56468 331974
rect 56416 331910 56468 331916
rect 56324 297424 56376 297430
rect 56324 297366 56376 297372
rect 56232 280084 56284 280090
rect 56232 280026 56284 280032
rect 56140 276072 56192 276078
rect 56140 276014 56192 276020
rect 55220 268456 55272 268462
rect 55220 268398 55272 268404
rect 55232 267034 55260 268398
rect 55220 267028 55272 267034
rect 55220 266970 55272 266976
rect 55128 237312 55180 237318
rect 55128 237254 55180 237260
rect 56152 209098 56180 276014
rect 56324 267028 56376 267034
rect 56324 266970 56376 266976
rect 56232 249076 56284 249082
rect 56232 249018 56284 249024
rect 56244 248470 56272 249018
rect 56232 248464 56284 248470
rect 56232 248406 56284 248412
rect 56244 226234 56272 248406
rect 56336 229090 56364 266970
rect 56428 260846 56456 331910
rect 56520 297401 56548 386514
rect 57256 336734 57284 437446
rect 57348 391950 57376 454038
rect 57716 439550 57744 537610
rect 57808 460222 57836 560254
rect 57900 556170 57928 697546
rect 59176 583976 59228 583982
rect 59176 583918 59228 583924
rect 59084 581188 59136 581194
rect 59084 581130 59136 581136
rect 57888 556164 57940 556170
rect 57888 556106 57940 556112
rect 59096 539034 59124 581130
rect 59084 539028 59136 539034
rect 59084 538970 59136 538976
rect 57888 538892 57940 538898
rect 57888 538834 57940 538840
rect 57796 460216 57848 460222
rect 57796 460158 57848 460164
rect 57808 458930 57836 460158
rect 57796 458924 57848 458930
rect 57796 458866 57848 458872
rect 57796 452736 57848 452742
rect 57796 452678 57848 452684
rect 57704 439544 57756 439550
rect 57704 439486 57756 439492
rect 57704 392692 57756 392698
rect 57704 392634 57756 392640
rect 57336 391944 57388 391950
rect 57336 391886 57388 391892
rect 57716 338026 57744 392634
rect 57808 355434 57836 452678
rect 57900 439006 57928 538834
rect 58992 494896 59044 494902
rect 58992 494838 59044 494844
rect 58624 491428 58676 491434
rect 58624 491370 58676 491376
rect 58636 491298 58664 491370
rect 58624 491292 58676 491298
rect 58624 491234 58676 491240
rect 57888 439000 57940 439006
rect 57888 438942 57940 438948
rect 57888 389360 57940 389366
rect 57888 389302 57940 389308
rect 57900 389201 57928 389302
rect 57886 389192 57942 389201
rect 57886 389127 57942 389136
rect 58636 388550 58664 491234
rect 59004 437238 59032 494838
rect 59188 493338 59216 583918
rect 59268 574116 59320 574122
rect 59268 574058 59320 574064
rect 59176 493332 59228 493338
rect 59176 493274 59228 493280
rect 59280 480254 59308 574058
rect 61844 572756 61896 572762
rect 61844 572698 61896 572704
rect 61752 568608 61804 568614
rect 61752 568550 61804 568556
rect 61108 562352 61160 562358
rect 61108 562294 61160 562300
rect 60372 561740 60424 561746
rect 60372 561682 60424 561688
rect 59096 480226 59308 480254
rect 59096 475454 59124 480226
rect 59084 475448 59136 475454
rect 59084 475390 59136 475396
rect 58992 437232 59044 437238
rect 58992 437174 59044 437180
rect 59096 434042 59124 475390
rect 59268 467900 59320 467906
rect 59268 467842 59320 467848
rect 59084 434036 59136 434042
rect 59084 433978 59136 433984
rect 58624 388544 58676 388550
rect 58624 388486 58676 388492
rect 58622 386472 58678 386481
rect 58622 386407 58678 386416
rect 58636 386374 58664 386407
rect 58624 386368 58676 386374
rect 58624 386310 58676 386316
rect 57888 378140 57940 378146
rect 57888 378082 57940 378088
rect 57796 355428 57848 355434
rect 57796 355370 57848 355376
rect 57704 338020 57756 338026
rect 57704 337962 57756 337968
rect 57244 336728 57296 336734
rect 57244 336670 57296 336676
rect 57808 330546 57836 355370
rect 57796 330540 57848 330546
rect 57796 330482 57848 330488
rect 57704 326460 57756 326466
rect 57704 326402 57756 326408
rect 56506 297392 56562 297401
rect 56506 297327 56562 297336
rect 56508 294704 56560 294710
rect 56508 294646 56560 294652
rect 56520 276010 56548 294646
rect 56508 276004 56560 276010
rect 56508 275946 56560 275952
rect 57716 263566 57744 326402
rect 57796 277432 57848 277438
rect 57796 277374 57848 277380
rect 57704 263560 57756 263566
rect 57704 263502 57756 263508
rect 56508 260908 56560 260914
rect 56508 260850 56560 260856
rect 56416 260840 56468 260846
rect 56416 260782 56468 260788
rect 56520 233170 56548 260850
rect 57704 258120 57756 258126
rect 57704 258062 57756 258068
rect 56508 233164 56560 233170
rect 56508 233106 56560 233112
rect 56324 229084 56376 229090
rect 56324 229026 56376 229032
rect 56232 226228 56284 226234
rect 56232 226170 56284 226176
rect 57716 220182 57744 258062
rect 57704 220176 57756 220182
rect 57704 220118 57756 220124
rect 56140 209092 56192 209098
rect 56140 209034 56192 209040
rect 55036 202224 55088 202230
rect 55036 202166 55088 202172
rect 53104 189032 53156 189038
rect 53104 188974 53156 188980
rect 57808 188358 57836 277374
rect 57796 188352 57848 188358
rect 57796 188294 57848 188300
rect 57796 125656 57848 125662
rect 57796 125598 57848 125604
rect 56508 122868 56560 122874
rect 56508 122810 56560 122816
rect 56520 93838 56548 122810
rect 56508 93832 56560 93838
rect 56508 93774 56560 93780
rect 57808 93770 57836 125598
rect 57796 93764 57848 93770
rect 57796 93706 57848 93712
rect 52368 71732 52420 71738
rect 52368 71674 52420 71680
rect 56600 58744 56652 58750
rect 56600 58686 56652 58692
rect 52460 57316 52512 57322
rect 52460 57258 52512 57264
rect 51080 56024 51132 56030
rect 51080 55966 51132 55972
rect 47584 33108 47636 33114
rect 47584 33050 47636 33056
rect 46940 22840 46992 22846
rect 46940 22782 46992 22788
rect 46952 16574 46980 22782
rect 49700 19984 49752 19990
rect 49700 19926 49752 19932
rect 49712 16574 49740 19926
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48504 13116 48556 13122
rect 48504 13058 48556 13064
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 13058
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 55966
rect 52472 3534 52500 57258
rect 53840 33856 53892 33862
rect 53840 33798 53892 33804
rect 52552 24132 52604 24138
rect 52552 24074 52604 24080
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 24074
rect 53852 16574 53880 33798
rect 56612 16574 56640 58686
rect 57900 58682 57928 378082
rect 58636 353297 58664 386310
rect 59082 383208 59138 383217
rect 59082 383143 59138 383152
rect 58622 353288 58678 353297
rect 58622 353223 58678 353232
rect 58992 344344 59044 344350
rect 58992 344286 59044 344292
rect 59004 343738 59032 344286
rect 58992 343732 59044 343738
rect 58992 343674 59044 343680
rect 59004 336025 59032 343674
rect 59096 339590 59124 383143
rect 59280 373318 59308 467842
rect 60384 463593 60412 561682
rect 61120 561678 61148 562294
rect 61108 561672 61160 561678
rect 61108 561614 61160 561620
rect 60464 560380 60516 560386
rect 60464 560322 60516 560328
rect 60370 463584 60426 463593
rect 60370 463519 60426 463528
rect 60476 461650 60504 560322
rect 60648 546508 60700 546514
rect 60648 546450 60700 546456
rect 60556 478848 60608 478854
rect 60556 478790 60608 478796
rect 60464 461644 60516 461650
rect 60464 461586 60516 461592
rect 60476 451274 60504 461586
rect 60384 451246 60504 451274
rect 59268 373312 59320 373318
rect 59268 373254 59320 373260
rect 59174 368384 59230 368393
rect 59174 368319 59230 368328
rect 59188 367713 59216 368319
rect 59174 367704 59230 367713
rect 59174 367639 59230 367648
rect 59084 339584 59136 339590
rect 59084 339526 59136 339532
rect 58990 336016 59046 336025
rect 58990 335951 59046 335960
rect 58992 301708 59044 301714
rect 58992 301650 59044 301656
rect 59004 285666 59032 301650
rect 59084 295996 59136 296002
rect 59084 295938 59136 295944
rect 58992 285660 59044 285666
rect 58992 285602 59044 285608
rect 59096 278730 59124 295938
rect 59084 278724 59136 278730
rect 59084 278666 59136 278672
rect 59084 269136 59136 269142
rect 59084 269078 59136 269084
rect 58716 240780 58768 240786
rect 58716 240722 58768 240728
rect 58728 237386 58756 240722
rect 58716 237380 58768 237386
rect 58716 237322 58768 237328
rect 59096 228410 59124 269078
rect 59084 228404 59136 228410
rect 59084 228346 59136 228352
rect 59188 61470 59216 367639
rect 59176 61464 59228 61470
rect 59176 61406 59228 61412
rect 57888 58676 57940 58682
rect 57888 58618 57940 58624
rect 59280 28286 59308 373254
rect 60384 365702 60412 451246
rect 60464 448588 60516 448594
rect 60464 448530 60516 448536
rect 60372 365696 60424 365702
rect 60372 365638 60424 365644
rect 60476 350606 60504 448530
rect 60568 384334 60596 478790
rect 60660 445754 60688 546450
rect 61384 470620 61436 470626
rect 61384 470562 61436 470568
rect 60740 445868 60792 445874
rect 60740 445810 60792 445816
rect 60752 445754 60780 445810
rect 60660 445726 60780 445754
rect 60556 384328 60608 384334
rect 60556 384270 60608 384276
rect 60464 350600 60516 350606
rect 60464 350542 60516 350548
rect 60464 312724 60516 312730
rect 60464 312666 60516 312672
rect 60476 274650 60504 312666
rect 60464 274644 60516 274650
rect 60464 274586 60516 274592
rect 60464 263696 60516 263702
rect 60464 263638 60516 263644
rect 60372 262268 60424 262274
rect 60372 262210 60424 262216
rect 60384 239562 60412 262210
rect 60372 239556 60424 239562
rect 60372 239498 60424 239504
rect 60476 233238 60504 263638
rect 60464 233232 60516 233238
rect 60464 233174 60516 233180
rect 59360 72480 59412 72486
rect 59360 72422 59412 72428
rect 59268 28280 59320 28286
rect 59268 28222 59320 28228
rect 57980 24200 58032 24206
rect 57980 24142 58032 24148
rect 57992 16574 58020 24142
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 16546
rect 56048 10328 56100 10334
rect 56048 10270 56100 10276
rect 56060 480 56088 10270
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 72422
rect 60568 69018 60596 384270
rect 60648 379636 60700 379642
rect 60648 379578 60700 379584
rect 60556 69012 60608 69018
rect 60556 68954 60608 68960
rect 60660 64870 60688 379578
rect 61396 375426 61424 470562
rect 61764 469606 61792 568550
rect 61856 474366 61884 572698
rect 62040 562358 62068 700266
rect 68836 594108 68888 594114
rect 68836 594050 68888 594056
rect 68468 585812 68520 585818
rect 68468 585754 68520 585760
rect 65892 583772 65944 583778
rect 65892 583714 65944 583720
rect 65524 581732 65576 581738
rect 65524 581674 65576 581680
rect 65536 581126 65564 581674
rect 65524 581120 65576 581126
rect 65524 581062 65576 581068
rect 64696 572008 64748 572014
rect 64696 571950 64748 571956
rect 64604 568676 64656 568682
rect 64604 568618 64656 568624
rect 63224 567248 63276 567254
rect 63224 567190 63276 567196
rect 62028 562352 62080 562358
rect 62028 562294 62080 562300
rect 61936 546576 61988 546582
rect 61936 546518 61988 546524
rect 61844 474360 61896 474366
rect 61844 474302 61896 474308
rect 61752 469600 61804 469606
rect 61752 469542 61804 469548
rect 61764 466454 61792 469542
rect 61764 466426 61884 466454
rect 61750 448624 61806 448633
rect 61750 448559 61752 448568
rect 61804 448559 61806 448568
rect 61752 448530 61804 448536
rect 61752 441516 61804 441522
rect 61752 441458 61804 441464
rect 61474 381032 61530 381041
rect 61474 380967 61530 380976
rect 61488 378146 61516 380967
rect 61476 378140 61528 378146
rect 61476 378082 61528 378088
rect 61384 375420 61436 375426
rect 61384 375362 61436 375368
rect 61764 340950 61792 441458
rect 61856 375358 61884 466426
rect 61948 448458 61976 546518
rect 62028 539640 62080 539646
rect 62028 539582 62080 539588
rect 61936 448452 61988 448458
rect 61936 448394 61988 448400
rect 61936 445868 61988 445874
rect 61936 445810 61988 445816
rect 61948 445777 61976 445810
rect 61934 445768 61990 445777
rect 61934 445703 61990 445712
rect 62040 441590 62068 539582
rect 63130 477456 63186 477465
rect 63130 477391 63186 477400
rect 62488 451512 62540 451518
rect 62488 451454 62540 451460
rect 62500 451178 62528 451454
rect 62488 451172 62540 451178
rect 62488 451114 62540 451120
rect 62120 448452 62172 448458
rect 62120 448394 62172 448400
rect 62132 447234 62160 448394
rect 62120 447228 62172 447234
rect 62120 447170 62172 447176
rect 62028 441584 62080 441590
rect 62028 441526 62080 441532
rect 61844 375352 61896 375358
rect 61844 375294 61896 375300
rect 62028 374672 62080 374678
rect 62028 374614 62080 374620
rect 61936 371884 61988 371890
rect 61936 371826 61988 371832
rect 61844 350600 61896 350606
rect 61844 350542 61896 350548
rect 61752 340944 61804 340950
rect 61752 340886 61804 340892
rect 61856 66230 61884 350542
rect 61948 73846 61976 371826
rect 61936 73840 61988 73846
rect 61936 73782 61988 73788
rect 61844 66224 61896 66230
rect 61844 66166 61896 66172
rect 60648 64864 60700 64870
rect 60648 64806 60700 64812
rect 60740 53236 60792 53242
rect 60740 53178 60792 53184
rect 60752 3534 60780 53178
rect 62040 44878 62068 374614
rect 62132 349178 62160 447170
rect 62764 442468 62816 442474
rect 62764 442410 62816 442416
rect 62120 349172 62172 349178
rect 62120 349114 62172 349120
rect 62776 343670 62804 442410
rect 63144 382265 63172 477391
rect 63236 467906 63264 567190
rect 63408 542496 63460 542502
rect 63408 542438 63460 542444
rect 63316 541000 63368 541006
rect 63316 540942 63368 540948
rect 63224 467900 63276 467906
rect 63224 467842 63276 467848
rect 63328 441522 63356 540942
rect 63420 442474 63448 542438
rect 64420 478916 64472 478922
rect 64420 478858 64472 478864
rect 64144 468376 64196 468382
rect 64144 468318 64196 468324
rect 64156 458930 64184 468318
rect 64144 458924 64196 458930
rect 64144 458866 64196 458872
rect 64144 455388 64196 455394
rect 64144 455330 64196 455336
rect 63408 442468 63460 442474
rect 63408 442410 63460 442416
rect 63316 441516 63368 441522
rect 63316 441458 63368 441464
rect 63224 389224 63276 389230
rect 63224 389166 63276 389172
rect 63130 382256 63186 382265
rect 63130 382191 63186 382200
rect 62764 343664 62816 343670
rect 62764 343606 62816 343612
rect 63132 255332 63184 255338
rect 63132 255274 63184 255280
rect 63144 239630 63172 255274
rect 63236 253842 63264 389166
rect 63408 375352 63460 375358
rect 63408 375294 63460 375300
rect 63420 374066 63448 375294
rect 63408 374060 63460 374066
rect 63408 374002 63460 374008
rect 63316 340944 63368 340950
rect 63316 340886 63368 340892
rect 63224 253836 63276 253842
rect 63224 253778 63276 253784
rect 63132 239624 63184 239630
rect 63132 239566 63184 239572
rect 63328 69766 63356 340886
rect 63420 75206 63448 374002
rect 64156 358766 64184 455330
rect 64432 386345 64460 478858
rect 64616 470558 64644 568618
rect 64708 473346 64736 571950
rect 64788 565888 64840 565894
rect 64788 565830 64840 565836
rect 64696 473340 64748 473346
rect 64696 473282 64748 473288
rect 64708 472666 64736 473282
rect 64696 472660 64748 472666
rect 64696 472602 64748 472608
rect 64604 470552 64656 470558
rect 64604 470494 64656 470500
rect 64800 467838 64828 565830
rect 65904 557433 65932 583714
rect 67640 581256 67692 581262
rect 67638 581224 67640 581233
rect 67692 581224 67694 581233
rect 67638 581159 67694 581168
rect 66902 579184 66958 579193
rect 66902 579119 66958 579128
rect 65984 573368 66036 573374
rect 65984 573310 66036 573316
rect 65890 557424 65946 557433
rect 65890 557359 65946 557368
rect 65892 483676 65944 483682
rect 65892 483618 65944 483624
rect 65798 478952 65854 478961
rect 65798 478887 65800 478896
rect 65852 478887 65854 478896
rect 65800 478858 65852 478864
rect 64788 467832 64840 467838
rect 64788 467774 64840 467780
rect 64788 458924 64840 458930
rect 64788 458866 64840 458872
rect 64512 441584 64564 441590
rect 64512 441526 64564 441532
rect 64524 440978 64552 441526
rect 64512 440972 64564 440978
rect 64512 440914 64564 440920
rect 64418 386336 64474 386345
rect 64418 386271 64474 386280
rect 64144 358760 64196 358766
rect 64144 358702 64196 358708
rect 63500 352572 63552 352578
rect 63500 352514 63552 352520
rect 63512 351966 63540 352514
rect 63500 351960 63552 351966
rect 63500 351902 63552 351908
rect 64420 351960 64472 351966
rect 64420 351902 64472 351908
rect 64432 349897 64460 351902
rect 64418 349888 64474 349897
rect 64418 349823 64474 349832
rect 64524 339522 64552 440914
rect 64696 375420 64748 375426
rect 64696 375362 64748 375368
rect 64602 349752 64658 349761
rect 64602 349687 64658 349696
rect 64512 339516 64564 339522
rect 64512 339458 64564 339464
rect 64512 302252 64564 302258
rect 64512 302194 64564 302200
rect 64524 262206 64552 302194
rect 64512 262200 64564 262206
rect 64512 262142 64564 262148
rect 63408 75200 63460 75206
rect 63408 75142 63460 75148
rect 63316 69760 63368 69766
rect 63316 69702 63368 69708
rect 62120 66904 62172 66910
rect 62120 66846 62172 66852
rect 62028 44872 62080 44878
rect 62028 44814 62080 44820
rect 60832 33788 60884 33794
rect 60832 33730 60884 33736
rect 60740 3528 60792 3534
rect 60740 3470 60792 3476
rect 60844 480 60872 33730
rect 62132 16574 62160 66846
rect 64616 49094 64644 349687
rect 64604 49088 64656 49094
rect 64604 49030 64656 49036
rect 64708 47598 64736 375362
rect 64800 360874 64828 458866
rect 65524 445800 65576 445806
rect 65524 445742 65576 445748
rect 64788 360868 64840 360874
rect 64788 360810 64840 360816
rect 64696 47592 64748 47598
rect 64696 47534 64748 47540
rect 63500 22772 63552 22778
rect 63500 22714 63552 22720
rect 63512 16574 63540 22714
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 61660 3528 61712 3534
rect 61660 3470 61712 3476
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3470
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 64800 12442 64828 360810
rect 65536 347750 65564 445742
rect 65904 438326 65932 483618
rect 65996 475386 66024 573310
rect 66076 567316 66128 567322
rect 66076 567258 66128 567264
rect 65984 475380 66036 475386
rect 65984 475322 66036 475328
rect 65984 474360 66036 474366
rect 65982 474328 65984 474337
rect 66036 474328 66038 474337
rect 65982 474263 66038 474272
rect 65984 470552 66036 470558
rect 65984 470494 66036 470500
rect 65892 438320 65944 438326
rect 65892 438262 65944 438268
rect 65996 383654 66024 470494
rect 66088 467945 66116 567258
rect 66168 558340 66220 558346
rect 66168 558282 66220 558288
rect 66074 467936 66130 467945
rect 66074 467871 66130 467880
rect 66076 465384 66128 465390
rect 66076 465326 66128 465332
rect 65904 383626 66024 383654
rect 65616 379500 65668 379506
rect 65616 379442 65668 379448
rect 65524 347744 65576 347750
rect 65524 347686 65576 347692
rect 65628 318102 65656 379442
rect 65904 374678 65932 383626
rect 65984 379704 66036 379710
rect 65984 379646 66036 379652
rect 65996 379506 66024 379646
rect 65984 379500 66036 379506
rect 65984 379442 66036 379448
rect 65892 374672 65944 374678
rect 65892 374614 65944 374620
rect 66088 369510 66116 465326
rect 66180 459542 66208 558282
rect 66916 482322 66944 579119
rect 67638 578504 67694 578513
rect 67638 578439 67694 578448
rect 67652 578270 67680 578439
rect 67640 578264 67692 578270
rect 67640 578206 67692 578212
rect 67454 577144 67510 577153
rect 67454 577079 67510 577088
rect 67468 489914 67496 577079
rect 67638 575784 67694 575793
rect 67638 575719 67694 575728
rect 67652 575550 67680 575719
rect 67640 575544 67692 575550
rect 67640 575486 67692 575492
rect 67638 574424 67694 574433
rect 67638 574359 67694 574368
rect 67652 574122 67680 574359
rect 67640 574116 67692 574122
rect 67640 574058 67692 574064
rect 68098 573472 68154 573481
rect 68098 573407 68154 573416
rect 68112 573374 68140 573407
rect 68100 573368 68152 573374
rect 68100 573310 68152 573316
rect 67638 572792 67694 572801
rect 67638 572727 67640 572736
rect 67692 572727 67694 572736
rect 67640 572698 67692 572704
rect 67824 572008 67876 572014
rect 67824 571950 67876 571956
rect 67836 571713 67864 571950
rect 68480 571713 68508 585754
rect 68848 582374 68876 594050
rect 68756 582346 68876 582374
rect 68756 576586 68784 582346
rect 68756 576558 68876 576586
rect 68742 576464 68798 576473
rect 68742 576399 68798 576408
rect 67822 571704 67878 571713
rect 67822 571639 67878 571648
rect 68466 571704 68522 571713
rect 68466 571639 68522 571648
rect 67638 570072 67694 570081
rect 67638 570007 67694 570016
rect 67652 569974 67680 570007
rect 67640 569968 67692 569974
rect 67640 569910 67692 569916
rect 67730 568984 67786 568993
rect 67730 568919 67786 568928
rect 67638 568712 67694 568721
rect 67744 568682 67772 568919
rect 67638 568647 67694 568656
rect 67732 568676 67784 568682
rect 67652 568614 67680 568647
rect 67732 568618 67784 568624
rect 67640 568608 67692 568614
rect 67640 568550 67692 568556
rect 67638 567624 67694 567633
rect 67638 567559 67694 567568
rect 67652 567254 67680 567559
rect 67732 567316 67784 567322
rect 67732 567258 67784 567264
rect 67640 567248 67692 567254
rect 67744 567225 67772 567258
rect 67640 567190 67692 567196
rect 67730 567216 67786 567225
rect 67730 567151 67786 567160
rect 67640 565888 67692 565894
rect 67638 565856 67640 565865
rect 67692 565856 67694 565865
rect 67638 565791 67694 565800
rect 67638 564904 67694 564913
rect 67638 564839 67694 564848
rect 67652 564534 67680 564839
rect 67640 564528 67692 564534
rect 67546 564496 67602 564505
rect 67640 564470 67692 564476
rect 67546 564431 67602 564440
rect 67284 489886 67496 489914
rect 66994 485752 67050 485761
rect 66994 485687 67050 485696
rect 66904 482316 66956 482322
rect 66904 482258 66956 482264
rect 66168 459536 66220 459542
rect 66168 459478 66220 459484
rect 66180 458862 66208 459478
rect 66168 458856 66220 458862
rect 66168 458798 66220 458804
rect 67008 439618 67036 485687
rect 67284 478854 67312 489886
rect 67364 482452 67416 482458
rect 67364 482394 67416 482400
rect 67272 478848 67324 478854
rect 67272 478790 67324 478796
rect 67284 478553 67312 478790
rect 67270 478544 67326 478553
rect 67270 478479 67326 478488
rect 66996 439612 67048 439618
rect 66996 439554 67048 439560
rect 67376 439142 67404 482394
rect 67456 482316 67508 482322
rect 67456 482258 67508 482264
rect 67468 481681 67496 482258
rect 67454 481672 67510 481681
rect 67454 481607 67510 481616
rect 67456 467832 67508 467838
rect 67456 467774 67508 467780
rect 67468 466857 67496 467774
rect 67454 466848 67510 466857
rect 67454 466783 67510 466792
rect 67364 439136 67416 439142
rect 67364 439078 67416 439084
rect 66166 379672 66222 379681
rect 66166 379607 66168 379616
rect 66220 379607 66222 379616
rect 66168 379578 66220 379584
rect 66904 376712 66956 376718
rect 66904 376654 66956 376660
rect 66166 369744 66222 369753
rect 66166 369679 66222 369688
rect 66076 369504 66128 369510
rect 66076 369446 66128 369452
rect 66076 365696 66128 365702
rect 66074 365664 66076 365673
rect 66128 365664 66130 365673
rect 66074 365599 66130 365608
rect 66076 347744 66128 347750
rect 66076 347686 66128 347692
rect 66088 347002 66116 347686
rect 66076 346996 66128 347002
rect 66076 346938 66128 346944
rect 65616 318096 65668 318102
rect 65616 318038 65668 318044
rect 66088 303006 66116 346938
rect 66180 337929 66208 369679
rect 66166 337920 66222 337929
rect 66166 337855 66222 337864
rect 66168 310548 66220 310554
rect 66168 310490 66220 310496
rect 66076 303000 66128 303006
rect 66076 302942 66128 302948
rect 65524 298240 65576 298246
rect 65524 298182 65576 298188
rect 65536 284306 65564 298182
rect 66076 291848 66128 291854
rect 66076 291790 66128 291796
rect 66088 286346 66116 291790
rect 66076 286340 66128 286346
rect 66076 286282 66128 286288
rect 65524 284300 65576 284306
rect 65524 284242 65576 284248
rect 65984 270564 66036 270570
rect 65984 270506 66036 270512
rect 65996 239494 66024 270506
rect 66076 258188 66128 258194
rect 66076 258130 66128 258136
rect 65984 239488 66036 239494
rect 65984 239430 66036 239436
rect 66088 224330 66116 258130
rect 66180 251190 66208 310490
rect 66916 301374 66944 376654
rect 67468 372722 67496 466783
rect 67560 465390 67588 564431
rect 67638 563544 67694 563553
rect 67638 563479 67694 563488
rect 67652 563106 67680 563479
rect 67640 563100 67692 563106
rect 67640 563042 67692 563048
rect 67640 562352 67692 562358
rect 67638 562320 67640 562329
rect 67692 562320 67694 562329
rect 67638 562255 67694 562264
rect 67638 562184 67694 562193
rect 67638 562119 67694 562128
rect 67652 561746 67680 562119
rect 67640 561740 67692 561746
rect 67640 561682 67692 561688
rect 67730 560824 67786 560833
rect 67730 560759 67786 560768
rect 67638 560416 67694 560425
rect 67744 560386 67772 560759
rect 67638 560351 67694 560360
rect 67732 560380 67784 560386
rect 67652 560318 67680 560351
rect 67732 560322 67784 560328
rect 67640 560312 67692 560318
rect 67640 560254 67692 560260
rect 67638 559464 67694 559473
rect 67638 559399 67694 559408
rect 67652 558958 67680 559399
rect 67640 558952 67692 558958
rect 67640 558894 67692 558900
rect 67640 557592 67692 557598
rect 67638 557560 67640 557569
rect 67692 557560 67694 557569
rect 67638 557495 67694 557504
rect 67822 556744 67878 556753
rect 67822 556679 67878 556688
rect 67640 556300 67692 556306
rect 67640 556242 67692 556248
rect 67652 556209 67680 556242
rect 67836 556238 67864 556679
rect 67824 556232 67876 556238
rect 67638 556200 67694 556209
rect 67824 556174 67876 556180
rect 67638 556135 67694 556144
rect 67732 556164 67784 556170
rect 67732 556106 67784 556112
rect 67638 555384 67694 555393
rect 67638 555319 67694 555328
rect 67652 554810 67680 555319
rect 67744 554849 67772 556106
rect 67730 554840 67786 554849
rect 67640 554804 67692 554810
rect 67730 554775 67786 554784
rect 67640 554746 67692 554752
rect 67638 553480 67694 553489
rect 67638 553415 67640 553424
rect 67692 553415 67694 553424
rect 67640 553386 67692 553392
rect 67638 552120 67694 552129
rect 67638 552055 67640 552064
rect 67692 552055 67694 552064
rect 67640 552026 67692 552032
rect 67638 551304 67694 551313
rect 67638 551239 67694 551248
rect 67652 550662 67680 551239
rect 68650 550760 68706 550769
rect 68650 550695 68706 550704
rect 67640 550656 67692 550662
rect 67640 550598 67692 550604
rect 67638 549944 67694 549953
rect 67638 549879 67694 549888
rect 67652 549302 67680 549879
rect 67640 549296 67692 549302
rect 67640 549238 67692 549244
rect 67730 548584 67786 548593
rect 67730 548519 67786 548528
rect 67638 548040 67694 548049
rect 67638 547975 67640 547984
rect 67692 547975 67694 547984
rect 67640 547946 67692 547952
rect 67744 547942 67772 548519
rect 67732 547936 67784 547942
rect 67732 547878 67784 547884
rect 67730 547224 67786 547233
rect 67730 547159 67786 547168
rect 67744 546582 67772 547159
rect 67732 546576 67784 546582
rect 67638 546544 67694 546553
rect 67732 546518 67784 546524
rect 67638 546479 67640 546488
rect 67692 546479 67694 546488
rect 67640 546450 67692 546456
rect 68558 545320 68614 545329
rect 68558 545255 68614 545264
rect 68572 545154 68600 545255
rect 68560 545148 68612 545154
rect 68560 545090 68612 545096
rect 68190 544504 68246 544513
rect 68190 544439 68246 544448
rect 68008 544400 68060 544406
rect 68008 544342 68060 544348
rect 68020 543969 68048 544342
rect 68006 543960 68062 543969
rect 68006 543895 68062 543904
rect 67730 543144 67786 543153
rect 67730 543079 67786 543088
rect 67638 542600 67694 542609
rect 67638 542535 67694 542544
rect 67652 542502 67680 542535
rect 67640 542496 67692 542502
rect 67640 542438 67692 542444
rect 67744 542434 67772 543079
rect 67732 542428 67784 542434
rect 67732 542370 67784 542376
rect 67638 541240 67694 541249
rect 67638 541175 67694 541184
rect 67652 541006 67680 541175
rect 67640 541000 67692 541006
rect 67640 540942 67692 540948
rect 67638 540152 67694 540161
rect 67638 540087 67694 540096
rect 67652 539646 67680 540087
rect 67640 539640 67692 539646
rect 67640 539582 67692 539588
rect 67640 488504 67692 488510
rect 67640 488446 67692 488452
rect 67652 488073 67680 488446
rect 67638 488064 67694 488073
rect 67638 487999 67694 488008
rect 67638 487928 67694 487937
rect 67638 487863 67694 487872
rect 67652 487830 67680 487863
rect 67640 487824 67692 487830
rect 67640 487766 67692 487772
rect 68008 487144 68060 487150
rect 68008 487086 68060 487092
rect 68020 486713 68048 487086
rect 68006 486704 68062 486713
rect 68006 486639 68062 486648
rect 67638 485208 67694 485217
rect 67638 485143 67694 485152
rect 67652 484430 67680 485143
rect 67640 484424 67692 484430
rect 67640 484366 67692 484372
rect 67638 483712 67694 483721
rect 67638 483647 67640 483656
rect 67692 483647 67694 483656
rect 67640 483618 67692 483624
rect 68100 482996 68152 483002
rect 68100 482938 68152 482944
rect 68112 482497 68140 482938
rect 68098 482488 68154 482497
rect 68098 482423 68154 482432
rect 67640 480208 67692 480214
rect 67640 480150 67692 480156
rect 67652 479913 67680 480150
rect 67638 479904 67694 479913
rect 67638 479839 67694 479848
rect 67730 477456 67786 477465
rect 67730 477391 67786 477400
rect 67638 476368 67694 476377
rect 67638 476303 67694 476312
rect 67652 476134 67680 476303
rect 67744 476241 67772 477391
rect 67730 476232 67786 476241
rect 67730 476167 67786 476176
rect 67640 476128 67692 476134
rect 67640 476070 67692 476076
rect 67638 475688 67694 475697
rect 67638 475623 67694 475632
rect 67652 475454 67680 475623
rect 67640 475448 67692 475454
rect 67640 475390 67692 475396
rect 67732 475380 67784 475386
rect 67732 475322 67784 475328
rect 67744 475153 67772 475322
rect 67730 475144 67786 475153
rect 67730 475079 67786 475088
rect 67640 474360 67692 474366
rect 67638 474328 67640 474337
rect 67692 474328 67694 474337
rect 67638 474263 67694 474272
rect 67640 473340 67692 473346
rect 67640 473282 67692 473288
rect 67652 472705 67680 473282
rect 67638 472696 67694 472705
rect 67638 472631 67694 472640
rect 67638 470928 67694 470937
rect 67638 470863 67694 470872
rect 67652 470626 67680 470863
rect 67640 470620 67692 470626
rect 67640 470562 67692 470568
rect 67732 470552 67784 470558
rect 67732 470494 67784 470500
rect 67744 470393 67772 470494
rect 67730 470384 67786 470393
rect 67730 470319 67786 470328
rect 67640 469600 67692 469606
rect 67638 469568 67640 469577
rect 67692 469568 67694 469577
rect 67638 469503 67694 469512
rect 67638 468208 67694 468217
rect 67638 468143 67694 468152
rect 67652 467906 67680 468143
rect 67640 467900 67692 467906
rect 67640 467842 67692 467848
rect 67640 465724 67692 465730
rect 67640 465666 67692 465672
rect 67652 465633 67680 465666
rect 67638 465624 67694 465633
rect 67638 465559 67694 465568
rect 67914 465488 67970 465497
rect 67914 465423 67970 465432
rect 67928 465390 67956 465423
rect 67548 465384 67600 465390
rect 67548 465326 67600 465332
rect 67916 465384 67968 465390
rect 67916 465326 67968 465332
rect 67640 464364 67692 464370
rect 67640 464306 67692 464312
rect 67652 464273 67680 464306
rect 67638 464264 67694 464273
rect 67638 464199 67694 464208
rect 67638 463448 67694 463457
rect 67638 463383 67694 463392
rect 67652 463010 67680 463383
rect 67640 463004 67692 463010
rect 67640 462946 67692 462952
rect 67640 461644 67692 461650
rect 67640 461586 67692 461592
rect 67652 461553 67680 461586
rect 67638 461544 67694 461553
rect 67638 461479 67694 461488
rect 67640 460216 67692 460222
rect 67638 460184 67640 460193
rect 67692 460184 67694 460193
rect 67638 460119 67694 460128
rect 67638 460048 67694 460057
rect 67638 459983 67694 459992
rect 67652 459610 67680 459983
rect 67640 459604 67692 459610
rect 67640 459546 67692 459552
rect 67732 459536 67784 459542
rect 67730 459504 67732 459513
rect 67784 459504 67786 459513
rect 67730 459439 67786 459448
rect 67640 458924 67692 458930
rect 67640 458866 67692 458872
rect 67652 458833 67680 458866
rect 67638 458824 67694 458833
rect 67638 458759 67694 458768
rect 67732 458176 67784 458182
rect 67732 458118 67784 458124
rect 67638 458008 67694 458017
rect 67638 457943 67694 457952
rect 67652 457502 67680 457943
rect 67640 457496 67692 457502
rect 67744 457473 67772 458118
rect 67640 457438 67692 457444
rect 67730 457464 67786 457473
rect 67730 457399 67786 457408
rect 67638 455968 67694 455977
rect 67638 455903 67694 455912
rect 67652 455462 67680 455903
rect 67640 455456 67692 455462
rect 67640 455398 67692 455404
rect 67638 454608 67694 454617
rect 67638 454543 67694 454552
rect 67652 454102 67680 454543
rect 67640 454096 67692 454102
rect 67640 454038 67692 454044
rect 67730 453248 67786 453257
rect 67730 453183 67786 453192
rect 67640 452736 67692 452742
rect 67638 452704 67640 452713
rect 67692 452704 67694 452713
rect 67744 452674 67772 453183
rect 67638 452639 67694 452648
rect 67732 452668 67784 452674
rect 67732 452610 67784 452616
rect 67638 451888 67694 451897
rect 67638 451823 67694 451832
rect 67652 451518 67680 451823
rect 67640 451512 67692 451518
rect 67640 451454 67692 451460
rect 67640 451240 67692 451246
rect 67640 451182 67692 451188
rect 67652 450809 67680 451182
rect 67638 450800 67694 450809
rect 67638 450735 67694 450744
rect 67822 448624 67878 448633
rect 67822 448559 67878 448568
rect 67836 448526 67864 448559
rect 67824 448520 67876 448526
rect 67824 448462 67876 448468
rect 67638 447264 67694 447273
rect 67638 447199 67640 447208
rect 67692 447199 67694 447208
rect 67640 447170 67692 447176
rect 67730 446448 67786 446457
rect 67730 446383 67786 446392
rect 67638 445904 67694 445913
rect 67744 445874 67772 446383
rect 67638 445839 67694 445848
rect 67732 445868 67784 445874
rect 67652 445806 67680 445839
rect 67732 445810 67784 445816
rect 67640 445800 67692 445806
rect 67640 445742 67692 445748
rect 67638 443728 67694 443737
rect 67638 443663 67640 443672
rect 67692 443663 67694 443672
rect 67640 443634 67692 443640
rect 67638 442504 67694 442513
rect 67638 442439 67640 442448
rect 67692 442439 67694 442448
rect 67640 442410 67692 442416
rect 67638 442368 67694 442377
rect 67638 442303 67694 442312
rect 67652 442270 67680 442303
rect 67640 442264 67692 442270
rect 67640 442206 67692 442212
rect 67640 441516 67692 441522
rect 67640 441458 67692 441464
rect 67652 441153 67680 441458
rect 67638 441144 67694 441153
rect 67638 441079 67694 441088
rect 67638 441008 67694 441017
rect 67638 440943 67640 440952
rect 67692 440943 67694 440952
rect 67640 440914 67692 440920
rect 67836 431954 67864 448462
rect 68204 444417 68232 544439
rect 68664 460934 68692 550695
rect 68756 477057 68784 576399
rect 68848 558929 68876 576558
rect 68940 572529 68968 702442
rect 69020 700392 69072 700398
rect 69020 700334 69072 700340
rect 69032 580689 69060 700334
rect 70308 583908 70360 583914
rect 70308 583850 70360 583856
rect 70216 582616 70268 582622
rect 70216 582558 70268 582564
rect 69112 582412 69164 582418
rect 69112 582354 69164 582360
rect 69018 580680 69074 580689
rect 69018 580615 69074 580624
rect 69032 579698 69060 580615
rect 69020 579692 69072 579698
rect 69020 579634 69072 579640
rect 68926 572520 68982 572529
rect 68926 572455 68982 572464
rect 68940 571849 68968 572455
rect 68926 571840 68982 571849
rect 68926 571775 68982 571784
rect 68834 558920 68890 558929
rect 68834 558855 68890 558864
rect 68848 558346 68876 558855
rect 68836 558340 68888 558346
rect 68836 558282 68888 558288
rect 69124 545329 69152 582354
rect 69846 581360 69902 581369
rect 69902 581318 70058 581346
rect 69846 581295 69902 581304
rect 69110 545320 69166 545329
rect 69110 545255 69166 545264
rect 68926 543960 68982 543969
rect 68926 543895 68982 543904
rect 68742 477048 68798 477057
rect 68742 476983 68798 476992
rect 68664 460906 68784 460934
rect 68756 451353 68784 460906
rect 68742 451344 68798 451353
rect 68742 451279 68798 451288
rect 68190 444408 68246 444417
rect 68190 444343 68246 444352
rect 68282 443864 68338 443873
rect 68282 443799 68338 443808
rect 67744 431926 67864 431954
rect 67744 400353 67772 431926
rect 67730 400344 67786 400353
rect 67730 400279 67786 400288
rect 67548 390652 67600 390658
rect 67548 390594 67600 390600
rect 67560 390522 67588 390594
rect 67548 390516 67600 390522
rect 67548 390458 67600 390464
rect 67638 384704 67694 384713
rect 67638 384639 67694 384648
rect 67652 384334 67680 384639
rect 67640 384328 67692 384334
rect 67640 384270 67692 384276
rect 67638 382528 67694 382537
rect 67638 382463 67694 382472
rect 67652 382294 67680 382463
rect 67640 382288 67692 382294
rect 67640 382230 67692 382236
rect 67730 379808 67786 379817
rect 67730 379743 67786 379752
rect 67744 379710 67772 379743
rect 67732 379704 67784 379710
rect 67638 379672 67694 379681
rect 67732 379646 67784 379652
rect 67638 379607 67640 379616
rect 67692 379607 67694 379616
rect 67640 379578 67692 379584
rect 67640 378140 67692 378146
rect 67640 378082 67692 378088
rect 67546 377360 67602 377369
rect 67546 377295 67602 377304
rect 67560 376718 67588 377295
rect 67652 377233 67680 378082
rect 67638 377224 67694 377233
rect 67638 377159 67694 377168
rect 67548 376712 67600 376718
rect 67548 376654 67600 376660
rect 67638 375592 67694 375601
rect 67638 375527 67694 375536
rect 67652 375426 67680 375527
rect 67640 375420 67692 375426
rect 67640 375362 67692 375368
rect 67640 374672 67692 374678
rect 67638 374640 67640 374649
rect 67692 374640 67694 374649
rect 67638 374575 67694 374584
rect 67638 374232 67694 374241
rect 67638 374167 67694 374176
rect 67652 374066 67680 374167
rect 67640 374060 67692 374066
rect 67640 374002 67692 374008
rect 67640 373312 67692 373318
rect 67640 373254 67692 373260
rect 67652 373017 67680 373254
rect 67638 373008 67694 373017
rect 67638 372943 67694 372952
rect 67468 372694 67680 372722
rect 67652 371890 67680 372694
rect 67640 371884 67692 371890
rect 67640 371826 67692 371832
rect 67652 371793 67680 371826
rect 67638 371784 67694 371793
rect 67638 371719 67694 371728
rect 67640 368552 67692 368558
rect 67638 368520 67640 368529
rect 67692 368520 67694 368529
rect 67638 368455 67694 368464
rect 67640 367056 67692 367062
rect 67638 367024 67640 367033
rect 67692 367024 67694 367033
rect 67638 366959 67694 366968
rect 68296 364334 68324 443799
rect 68756 394670 68784 451279
rect 68834 444408 68890 444417
rect 68834 444343 68890 444352
rect 68744 394664 68796 394670
rect 68744 394606 68796 394612
rect 68376 369504 68428 369510
rect 68374 369472 68376 369481
rect 68428 369472 68430 369481
rect 68374 369407 68430 369416
rect 68742 369472 68798 369481
rect 68742 369407 68798 369416
rect 68296 364306 68508 364334
rect 67638 363760 67694 363769
rect 67638 363695 67694 363704
rect 67652 363662 67680 363695
rect 67640 363656 67692 363662
rect 67640 363598 67692 363604
rect 67546 361992 67602 362001
rect 67546 361927 67602 361936
rect 67560 361486 67588 361927
rect 68008 361548 68060 361554
rect 68008 361490 68060 361496
rect 66996 361480 67048 361486
rect 66996 361422 67048 361428
rect 67548 361480 67600 361486
rect 67548 361422 67600 361428
rect 67008 336054 67036 361422
rect 67638 360904 67694 360913
rect 67638 360839 67640 360848
rect 67692 360839 67694 360848
rect 67640 360810 67692 360816
rect 68020 360641 68048 361490
rect 68006 360632 68062 360641
rect 68006 360567 68062 360576
rect 67638 359544 67694 359553
rect 67638 359479 67640 359488
rect 67692 359479 67694 359488
rect 67640 359450 67692 359456
rect 67456 358760 67508 358766
rect 67640 358760 67692 358766
rect 67456 358702 67508 358708
rect 67638 358728 67640 358737
rect 67692 358728 67694 358737
rect 67180 339516 67232 339522
rect 67180 339458 67232 339464
rect 66996 336048 67048 336054
rect 66996 335990 67048 335996
rect 66904 301368 66956 301374
rect 66904 301310 66956 301316
rect 66168 251184 66220 251190
rect 66168 251126 66220 251132
rect 66168 247104 66220 247110
rect 66168 247046 66220 247052
rect 66076 224324 66128 224330
rect 66076 224266 66128 224272
rect 66180 189689 66208 247046
rect 66166 189680 66222 189689
rect 66166 189615 66222 189624
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65154 126304 65210 126313
rect 65154 126239 65210 126248
rect 65168 125662 65196 126239
rect 65156 125656 65208 125662
rect 65156 125598 65208 125604
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66074 102368 66130 102377
rect 66074 102303 66130 102312
rect 66088 84182 66116 102303
rect 66180 94897 66208 129231
rect 66166 94888 66222 94897
rect 66166 94823 66222 94832
rect 66076 84176 66128 84182
rect 66076 84118 66128 84124
rect 67192 45558 67220 339458
rect 67468 319666 67496 358702
rect 67638 358663 67694 358672
rect 67640 358080 67692 358086
rect 67638 358048 67640 358057
rect 67692 358048 67694 358057
rect 67638 357983 67694 357992
rect 67914 356960 67970 356969
rect 67914 356895 67970 356904
rect 67928 356114 67956 356895
rect 67916 356108 67968 356114
rect 67916 356050 67968 356056
rect 67730 355600 67786 355609
rect 67730 355535 67786 355544
rect 67640 355428 67692 355434
rect 67640 355370 67692 355376
rect 67652 355201 67680 355370
rect 67744 355366 67772 355535
rect 67732 355360 67784 355366
rect 67732 355302 67784 355308
rect 67638 355192 67694 355201
rect 67638 355127 67694 355136
rect 67638 352200 67694 352209
rect 67638 352135 67694 352144
rect 67652 351966 67680 352135
rect 67640 351960 67692 351966
rect 67640 351902 67692 351908
rect 67638 351112 67694 351121
rect 67638 351047 67694 351056
rect 67652 350606 67680 351047
rect 67640 350600 67692 350606
rect 67640 350542 67692 350548
rect 68006 350160 68062 350169
rect 68006 350095 68062 350104
rect 68020 349246 68048 350095
rect 68008 349240 68060 349246
rect 68008 349182 68060 349188
rect 67640 349104 67692 349110
rect 67638 349072 67640 349081
rect 67692 349072 67694 349081
rect 67638 349007 67694 349016
rect 68480 348242 68508 364306
rect 68560 359508 68612 359514
rect 68560 359450 68612 359456
rect 68572 353161 68600 359450
rect 68558 353152 68614 353161
rect 68558 353087 68614 353096
rect 68572 352646 68600 353087
rect 68560 352640 68612 352646
rect 68560 352582 68612 352588
rect 68480 348214 68692 348242
rect 67638 347032 67694 347041
rect 67638 346967 67640 346976
rect 67692 346967 67694 346976
rect 67640 346938 67692 346944
rect 68560 346384 68612 346390
rect 68560 346326 68612 346332
rect 67638 343768 67694 343777
rect 67638 343703 67640 343712
rect 67692 343703 67694 343712
rect 67640 343674 67692 343680
rect 67638 343632 67694 343641
rect 67638 343567 67640 343576
rect 67692 343567 67694 343576
rect 67640 343538 67692 343544
rect 67638 341048 67694 341057
rect 67638 340983 67694 340992
rect 67652 340950 67680 340983
rect 67640 340944 67692 340950
rect 67640 340886 67692 340892
rect 67638 340232 67694 340241
rect 67638 340167 67694 340176
rect 67652 339522 67680 340167
rect 67640 339516 67692 339522
rect 67640 339458 67692 339464
rect 68572 338910 68600 346326
rect 68664 345098 68692 348214
rect 68652 345092 68704 345098
rect 68652 345034 68704 345040
rect 68664 345001 68692 345034
rect 68650 344992 68706 345001
rect 68650 344927 68706 344936
rect 68652 342236 68704 342242
rect 68652 342178 68704 342184
rect 68664 342009 68692 342178
rect 68650 342000 68706 342009
rect 68650 341935 68706 341944
rect 68560 338904 68612 338910
rect 68560 338846 68612 338852
rect 68756 329118 68784 369407
rect 68848 346390 68876 444343
rect 68940 443873 68968 543895
rect 69018 541784 69074 541793
rect 69018 541719 69074 541728
rect 69032 525774 69060 541719
rect 69860 540110 70058 540138
rect 69860 536897 69888 540110
rect 69846 536888 69902 536897
rect 70228 536858 70256 582558
rect 70320 537742 70348 583850
rect 70952 583772 71004 583778
rect 70952 583714 71004 583720
rect 70964 581890 70992 583714
rect 71792 583030 71820 702986
rect 75184 702840 75236 702846
rect 75184 702782 75236 702788
rect 71872 596216 71924 596222
rect 71872 596158 71924 596164
rect 71780 583024 71832 583030
rect 71780 582966 71832 582972
rect 71884 582162 71912 596158
rect 74632 592068 74684 592074
rect 74632 592010 74684 592016
rect 73344 584112 73396 584118
rect 73344 584054 73396 584060
rect 72238 582448 72294 582457
rect 72238 582383 72294 582392
rect 71792 582134 71912 582162
rect 70964 581862 71300 581890
rect 71792 581754 71820 582134
rect 72252 581890 72280 582383
rect 73356 581890 73384 584054
rect 74644 581890 74672 592010
rect 75196 586514 75224 702782
rect 74920 586486 75224 586514
rect 74920 585342 74948 586486
rect 74908 585336 74960 585342
rect 74908 585278 74960 585284
rect 72252 581862 72588 581890
rect 73278 581862 73384 581890
rect 74566 581862 74672 581890
rect 74920 581890 74948 585278
rect 76576 583982 76604 702986
rect 77956 596174 77984 703258
rect 79324 702636 79376 702642
rect 79324 702578 79376 702584
rect 77956 596146 78076 596174
rect 78048 585206 78076 596146
rect 78036 585200 78088 585206
rect 78036 585142 78088 585148
rect 76564 583976 76616 583982
rect 76564 583918 76616 583924
rect 77852 583976 77904 583982
rect 77852 583918 77904 583924
rect 76576 581890 76604 583918
rect 77864 583846 77892 583918
rect 77852 583840 77904 583846
rect 77852 583782 77904 583788
rect 76748 582548 76800 582554
rect 76748 582490 76800 582496
rect 74920 581862 75164 581890
rect 76498 581862 76604 581890
rect 76760 581890 76788 582490
rect 77864 581890 77892 583782
rect 76760 581862 77096 581890
rect 77786 581862 77892 581890
rect 78048 581890 78076 585142
rect 78680 584044 78732 584050
rect 78680 583986 78732 583992
rect 78692 581890 78720 583986
rect 79336 583982 79364 702578
rect 89180 702434 89208 703520
rect 95148 703248 95200 703254
rect 95148 703190 95200 703196
rect 88352 702406 89208 702434
rect 87604 656940 87656 656946
rect 87604 656882 87656 656888
rect 85580 597576 85632 597582
rect 85580 597518 85632 597524
rect 85592 596174 85620 597518
rect 85592 596146 85712 596174
rect 81808 592680 81860 592686
rect 81808 592622 81860 592628
rect 80612 586560 80664 586566
rect 80612 586502 80664 586508
rect 79324 583976 79376 583982
rect 79324 583918 79376 583924
rect 80624 581890 80652 586502
rect 81820 583953 81848 592622
rect 85120 586764 85172 586770
rect 85120 586706 85172 586712
rect 81900 586696 81952 586702
rect 81900 586638 81952 586644
rect 81438 583944 81494 583953
rect 81438 583879 81494 583888
rect 81806 583944 81862 583953
rect 81806 583879 81862 583888
rect 81452 581890 81480 583879
rect 81912 581890 81940 586638
rect 84292 586628 84344 586634
rect 84292 586570 84344 586576
rect 83188 585268 83240 585274
rect 83188 585210 83240 585216
rect 83004 583908 83056 583914
rect 83004 583850 83056 583856
rect 83016 581890 83044 583850
rect 78048 581862 78384 581890
rect 78692 581862 79028 581890
rect 80624 581862 80960 581890
rect 81452 581862 81604 581890
rect 81912 581862 82248 581890
rect 82938 581862 83044 581890
rect 83200 581890 83228 585210
rect 84304 581890 84332 586570
rect 84476 582616 84528 582622
rect 84476 582558 84528 582564
rect 83200 581862 83536 581890
rect 84226 581862 84332 581890
rect 84488 581890 84516 582558
rect 85132 581890 85160 586706
rect 85684 581890 85712 596146
rect 87616 585410 87644 656882
rect 88352 588606 88380 702406
rect 88340 588600 88392 588606
rect 88340 588542 88392 588548
rect 92848 586696 92900 586702
rect 92848 586638 92900 586644
rect 89628 586560 89680 586566
rect 89628 586502 89680 586508
rect 87604 585404 87656 585410
rect 87604 585346 87656 585352
rect 87616 581890 87644 585346
rect 88984 584044 89036 584050
rect 88984 583986 89036 583992
rect 88246 583944 88302 583953
rect 88246 583879 88302 583888
rect 88260 581890 88288 583879
rect 88996 581890 89024 583986
rect 89640 581890 89668 586502
rect 91558 583808 91614 583817
rect 91558 583743 91614 583752
rect 91006 582584 91062 582593
rect 91006 582519 91062 582528
rect 91020 581890 91048 582519
rect 91572 581890 91600 583743
rect 92296 582684 92348 582690
rect 92296 582626 92348 582632
rect 92308 581890 92336 582626
rect 92860 581890 92888 586638
rect 94872 586628 94924 586634
rect 94872 586570 94924 586576
rect 94136 585336 94188 585342
rect 94136 585278 94188 585284
rect 94148 581890 94176 585278
rect 94884 581890 94912 586570
rect 95160 585177 95188 703190
rect 104808 702976 104860 702982
rect 104808 702918 104860 702924
rect 99288 698964 99340 698970
rect 99288 698906 99340 698912
rect 95424 587920 95476 587926
rect 95424 587862 95476 587868
rect 95146 585168 95202 585177
rect 84488 581862 84824 581890
rect 85132 581862 85468 581890
rect 85684 581862 86112 581890
rect 87446 581862 87644 581890
rect 88090 581862 88288 581890
rect 88734 581862 89024 581890
rect 89378 581862 89668 581890
rect 90666 581862 91048 581890
rect 91310 581862 91600 581890
rect 91954 581862 92336 581890
rect 92598 581862 92888 581890
rect 93886 581862 94176 581890
rect 94530 581862 94912 581890
rect 94976 585126 95146 585154
rect 94976 581754 95004 585126
rect 95146 585103 95202 585112
rect 95436 581890 95464 587862
rect 97908 586832 97960 586838
rect 97908 586774 97960 586780
rect 96528 583840 96580 583846
rect 96528 583782 96580 583788
rect 96540 581890 96568 583782
rect 97448 582616 97500 582622
rect 97448 582558 97500 582564
rect 97460 581890 97488 582558
rect 97920 581890 97948 586774
rect 99300 585478 99328 698906
rect 100576 586764 100628 586770
rect 100576 586706 100628 586712
rect 99288 585472 99340 585478
rect 99288 585414 99340 585420
rect 99300 585206 99328 585414
rect 98736 585200 98788 585206
rect 98736 585142 98788 585148
rect 99288 585200 99340 585206
rect 99288 585142 99340 585148
rect 98748 581890 98776 585142
rect 99288 582548 99340 582554
rect 99288 582490 99340 582496
rect 99300 581890 99328 582490
rect 100588 581890 100616 586706
rect 104820 584458 104848 702918
rect 105464 702434 105492 703520
rect 109684 703180 109736 703186
rect 109684 703122 109736 703128
rect 108948 702568 109000 702574
rect 108948 702510 109000 702516
rect 105464 702406 105584 702434
rect 105556 596174 105584 702406
rect 106280 697672 106332 697678
rect 106280 697614 106332 697620
rect 105556 596146 105676 596174
rect 103152 584452 103204 584458
rect 103152 584394 103204 584400
rect 104808 584452 104860 584458
rect 104808 584394 104860 584400
rect 101312 583976 101364 583982
rect 101312 583918 101364 583924
rect 101324 581890 101352 583918
rect 101862 582448 101918 582457
rect 101862 582383 101918 582392
rect 101876 581890 101904 582383
rect 103164 581890 103192 584394
rect 103888 583908 103940 583914
rect 103888 583850 103940 583856
rect 103900 581890 103928 583850
rect 105544 583772 105596 583778
rect 105544 583714 105596 583720
rect 105556 581890 105584 583714
rect 95436 581862 95772 581890
rect 96462 581862 96568 581890
rect 97106 581862 97488 581890
rect 97750 581862 97948 581890
rect 98394 581862 98776 581890
rect 99038 581862 99328 581890
rect 100326 581862 100616 581890
rect 100970 581862 101352 581890
rect 101614 581862 101904 581890
rect 102902 581862 103192 581890
rect 103546 581862 103928 581890
rect 105478 581862 105584 581890
rect 102598 581768 102654 581777
rect 71792 581726 71944 581754
rect 75472 581738 75808 581754
rect 79336 581738 79672 581754
rect 75460 581732 75808 581738
rect 75512 581726 75808 581732
rect 79324 581732 79672 581738
rect 75460 581674 75512 581680
rect 79376 581726 79672 581732
rect 90022 581738 90312 581754
rect 90022 581732 90324 581738
rect 90022 581726 90272 581732
rect 79324 581674 79376 581680
rect 94976 581726 95128 581754
rect 102258 581726 102598 581754
rect 104190 581738 104480 581754
rect 104834 581738 105032 581754
rect 104190 581732 104492 581738
rect 104190 581726 104440 581732
rect 102598 581703 102654 581712
rect 90272 581674 90324 581680
rect 104834 581732 105044 581738
rect 104834 581726 104992 581732
rect 104440 581674 104492 581680
rect 104992 581674 105044 581680
rect 70412 581318 70702 581346
rect 70412 581058 70440 581318
rect 70400 581052 70452 581058
rect 70400 580994 70452 581000
rect 105648 572014 105676 596146
rect 105636 572008 105688 572014
rect 105636 571950 105688 571956
rect 105634 561912 105690 561921
rect 105634 561847 105690 561856
rect 105648 557534 105676 561847
rect 106292 560425 106320 697614
rect 108960 586514 108988 702510
rect 108868 586486 108988 586514
rect 106922 583944 106978 583953
rect 106922 583879 106978 583888
rect 106936 567866 106964 583879
rect 107660 582480 107712 582486
rect 107660 582422 107712 582428
rect 107672 573345 107700 582422
rect 108868 577561 108896 586486
rect 109040 585472 109092 585478
rect 109040 585414 109092 585420
rect 108946 580816 109002 580825
rect 108946 580751 109002 580760
rect 108960 579766 108988 580751
rect 108948 579760 109000 579766
rect 108948 579702 109000 579708
rect 108946 579456 109002 579465
rect 108946 579391 109002 579400
rect 108960 578270 108988 579391
rect 108948 578264 109000 578270
rect 108948 578206 109000 578212
rect 108946 578096 109002 578105
rect 108946 578031 109002 578040
rect 108854 577552 108910 577561
rect 108854 577487 108910 577496
rect 108960 576910 108988 578031
rect 108948 576904 109000 576910
rect 108948 576846 109000 576852
rect 108762 576736 108818 576745
rect 108762 576671 108818 576680
rect 108776 575618 108804 576671
rect 108946 576056 109002 576065
rect 108946 575991 109002 576000
rect 108764 575612 108816 575618
rect 108764 575554 108816 575560
rect 108960 575550 108988 575991
rect 108948 575544 109000 575550
rect 108948 575486 109000 575492
rect 108946 574696 109002 574705
rect 108946 574631 109002 574640
rect 108960 574122 108988 574631
rect 108948 574116 109000 574122
rect 108948 574058 109000 574064
rect 108672 573368 108724 573374
rect 107658 573336 107714 573345
rect 107658 573271 107714 573280
rect 108670 573336 108672 573345
rect 108724 573336 108726 573345
rect 108670 573271 108726 573280
rect 107014 572792 107070 572801
rect 107014 572727 107070 572736
rect 106924 567860 106976 567866
rect 106924 567802 106976 567808
rect 106278 560416 106334 560425
rect 106278 560351 106334 560360
rect 105648 557506 105768 557534
rect 105478 540382 105676 540410
rect 70504 540110 70702 540138
rect 70308 537736 70360 537742
rect 70308 537678 70360 537684
rect 69846 536823 69902 536832
rect 70216 536852 70268 536858
rect 70216 536794 70268 536800
rect 70504 529310 70532 540110
rect 71332 538214 71360 540138
rect 70964 538186 71360 538214
rect 70492 529304 70544 529310
rect 70492 529246 70544 529252
rect 70964 528554 70992 538186
rect 71044 535424 71096 535430
rect 71044 535366 71096 535372
rect 70412 528526 70992 528554
rect 69020 525768 69072 525774
rect 69020 525710 69072 525716
rect 70412 497486 70440 528526
rect 70400 497480 70452 497486
rect 70400 497422 70452 497428
rect 70032 493332 70084 493338
rect 70032 493274 70084 493280
rect 70044 489940 70072 493274
rect 70400 491428 70452 491434
rect 70400 491370 70452 491376
rect 70412 489954 70440 491370
rect 71056 489977 71084 535366
rect 71976 526454 72004 540138
rect 72620 529378 72648 540138
rect 73160 539028 73212 539034
rect 73160 538970 73212 538976
rect 72608 529372 72660 529378
rect 72608 529314 72660 529320
rect 71964 526448 72016 526454
rect 71964 526390 72016 526396
rect 73172 499574 73200 538970
rect 73264 537606 73292 540138
rect 73908 538121 73936 540138
rect 73894 538112 73950 538121
rect 73894 538047 73950 538056
rect 73252 537600 73304 537606
rect 73252 537542 73304 537548
rect 74552 529242 74580 540138
rect 75092 536852 75144 536858
rect 75092 536794 75144 536800
rect 74540 529236 74592 529242
rect 74540 529178 74592 529184
rect 75104 528554 75132 536794
rect 75196 534886 75224 540138
rect 76467 540110 76512 540138
rect 75184 534880 75236 534886
rect 75184 534822 75236 534828
rect 76484 532166 76512 540110
rect 77128 535430 77156 540138
rect 77116 535424 77168 535430
rect 77116 535366 77168 535372
rect 76564 533384 76616 533390
rect 76564 533326 76616 533332
rect 76472 532160 76524 532166
rect 76472 532102 76524 532108
rect 75104 528526 75224 528554
rect 73172 499546 73292 499574
rect 71136 492720 71188 492726
rect 71136 492662 71188 492668
rect 71042 489968 71098 489977
rect 70412 489926 70656 489954
rect 71148 489954 71176 492662
rect 72240 492108 72292 492114
rect 72240 492050 72292 492056
rect 71780 491360 71832 491366
rect 71780 491302 71832 491308
rect 71792 489954 71820 491302
rect 72252 489954 72280 492050
rect 73264 489954 73292 499546
rect 74814 493368 74870 493377
rect 74814 493303 74870 493312
rect 74356 490000 74408 490006
rect 71148 489926 71300 489954
rect 71792 489926 71944 489954
rect 72252 489926 72588 489954
rect 73264 489940 73476 489954
rect 74828 489954 74856 493303
rect 75196 492658 75224 528526
rect 76576 499574 76604 533326
rect 77772 526425 77800 540138
rect 78416 534750 78444 540138
rect 78404 534744 78456 534750
rect 78404 534686 78456 534692
rect 77758 526416 77814 526425
rect 77758 526351 77814 526360
rect 76576 499546 76696 499574
rect 76472 496188 76524 496194
rect 76472 496130 76524 496136
rect 75460 494828 75512 494834
rect 75460 494770 75512 494776
rect 75184 492652 75236 492658
rect 75184 492594 75236 492600
rect 75472 489954 75500 494770
rect 74408 489948 74520 489954
rect 74356 489942 74520 489948
rect 73278 489938 73476 489940
rect 73278 489932 73488 489938
rect 73278 489926 73436 489932
rect 71042 489903 71098 489912
rect 74368 489926 74520 489942
rect 74828 489926 75164 489954
rect 75472 489926 75808 489954
rect 76484 489940 76512 496130
rect 76668 491638 76696 499546
rect 77392 494080 77444 494086
rect 77392 494022 77444 494028
rect 76656 491632 76708 491638
rect 76656 491574 76708 491580
rect 76668 489954 76696 491574
rect 77404 489954 77432 494022
rect 78404 492652 78456 492658
rect 78404 492594 78456 492600
rect 78416 491706 78444 492594
rect 78404 491700 78456 491706
rect 78404 491642 78456 491648
rect 76668 489926 77096 489954
rect 77404 489926 77740 489954
rect 78416 489940 78444 491642
rect 79060 490618 79088 540138
rect 79704 537606 79732 540138
rect 80348 538121 80376 540138
rect 80334 538112 80390 538121
rect 80334 538047 80390 538056
rect 79692 537600 79744 537606
rect 79692 537542 79744 537548
rect 79324 532092 79376 532098
rect 79324 532034 79376 532040
rect 79336 492833 79364 532034
rect 80992 494902 81020 540138
rect 81532 537736 81584 537742
rect 81532 537678 81584 537684
rect 81544 496194 81572 537678
rect 81636 537674 81664 540138
rect 82907 540110 82952 540138
rect 81624 537668 81676 537674
rect 81624 537610 81676 537616
rect 82924 537538 82952 540110
rect 83464 537668 83516 537674
rect 83464 537610 83516 537616
rect 82912 537532 82964 537538
rect 82912 537474 82964 537480
rect 81624 497480 81676 497486
rect 81624 497422 81676 497428
rect 81532 496188 81584 496194
rect 81532 496130 81584 496136
rect 80980 494896 81032 494902
rect 80980 494838 81032 494844
rect 80980 493332 81032 493338
rect 80980 493274 81032 493280
rect 79322 492824 79378 492833
rect 79322 492759 79378 492768
rect 79048 490612 79100 490618
rect 79048 490554 79100 490560
rect 79336 489954 79364 492759
rect 80060 492040 80112 492046
rect 80060 491982 80112 491988
rect 80072 489954 80100 491982
rect 79336 489926 79672 489954
rect 80072 489926 80316 489954
rect 80992 489940 81020 493274
rect 81636 489940 81664 497422
rect 82268 494896 82320 494902
rect 82268 494838 82320 494844
rect 82280 489940 82308 494838
rect 82912 494828 82964 494834
rect 82912 494770 82964 494776
rect 82820 494760 82872 494766
rect 82820 494702 82872 494708
rect 82832 494018 82860 494702
rect 82820 494012 82872 494018
rect 82820 493954 82872 493960
rect 82924 489940 82952 494770
rect 83476 491978 83504 537610
rect 83568 534818 83596 540138
rect 84212 537538 84240 540138
rect 84200 537532 84252 537538
rect 84200 537474 84252 537480
rect 84856 536858 84884 540138
rect 84108 536852 84160 536858
rect 84108 536794 84160 536800
rect 84844 536852 84896 536858
rect 84844 536794 84896 536800
rect 83556 534812 83608 534818
rect 83556 534754 83608 534760
rect 84120 497554 84148 536794
rect 85500 497622 85528 540138
rect 86144 532030 86172 540138
rect 86132 532024 86184 532030
rect 86132 531966 86184 531972
rect 85488 497616 85540 497622
rect 85488 497558 85540 497564
rect 84108 497548 84160 497554
rect 84108 497490 84160 497496
rect 86788 497457 86816 540138
rect 87052 537600 87104 537606
rect 87052 537542 87104 537548
rect 86774 497448 86830 497457
rect 86774 497383 86830 497392
rect 84842 496088 84898 496097
rect 84842 496023 84898 496032
rect 83556 494012 83608 494018
rect 83556 493954 83608 493960
rect 83464 491972 83516 491978
rect 83464 491914 83516 491920
rect 83568 489940 83596 493954
rect 84856 489940 84884 496023
rect 85488 493196 85540 493202
rect 85488 493138 85540 493144
rect 85500 489940 85528 493138
rect 86132 491972 86184 491978
rect 86132 491914 86184 491920
rect 86144 489940 86172 491914
rect 86776 491428 86828 491434
rect 86776 491370 86828 491376
rect 86788 489940 86816 491370
rect 87064 490521 87092 537542
rect 87432 532098 87460 540138
rect 88076 539034 88104 540138
rect 89347 540110 89392 540138
rect 88064 539028 88116 539034
rect 88064 538970 88116 538976
rect 87420 532092 87472 532098
rect 87420 532034 87472 532040
rect 88248 500336 88300 500342
rect 88248 500278 88300 500284
rect 88260 497486 88288 500278
rect 89364 498846 89392 540110
rect 90008 534750 90036 540138
rect 90364 538960 90416 538966
rect 90364 538902 90416 538908
rect 89996 534744 90048 534750
rect 89626 534712 89682 534721
rect 89996 534686 90048 534692
rect 89626 534647 89682 534656
rect 89640 499574 89668 534647
rect 89548 499546 89668 499574
rect 89352 498840 89404 498846
rect 89352 498782 89404 498788
rect 88248 497480 88300 497486
rect 88248 497422 88300 497428
rect 88064 496324 88116 496330
rect 88064 496266 88116 496272
rect 87420 490748 87472 490754
rect 87420 490690 87472 490696
rect 87050 490512 87106 490521
rect 87050 490447 87106 490456
rect 87432 489940 87460 490690
rect 88076 489940 88104 496266
rect 89548 493882 89576 499546
rect 89628 496256 89680 496262
rect 89628 496198 89680 496204
rect 88708 493876 88760 493882
rect 88708 493818 88760 493824
rect 89536 493876 89588 493882
rect 89536 493818 89588 493824
rect 88720 492726 88748 493818
rect 89640 493202 89668 496198
rect 89628 493196 89680 493202
rect 89628 493138 89680 493144
rect 88708 492720 88760 492726
rect 88708 492662 88760 492668
rect 88720 489940 88748 492662
rect 90376 491502 90404 538902
rect 90652 537674 90680 540138
rect 91296 538898 91324 540138
rect 91284 538892 91336 538898
rect 91284 538834 91336 538840
rect 90640 537668 90692 537674
rect 90640 537610 90692 537616
rect 91940 499574 91968 540138
rect 91940 499546 92060 499574
rect 91100 496120 91152 496126
rect 91100 496062 91152 496068
rect 91112 495514 91140 496062
rect 91100 495508 91152 495514
rect 91100 495450 91152 495456
rect 90640 494760 90692 494766
rect 90640 494702 90692 494708
rect 90364 491496 90416 491502
rect 90364 491438 90416 491444
rect 90376 489954 90404 491438
rect 90022 489926 90404 489954
rect 90652 489940 90680 494702
rect 91112 489954 91140 495450
rect 91928 492040 91980 492046
rect 91928 491982 91980 491988
rect 91112 489926 91264 489954
rect 91940 489940 91968 491982
rect 92032 490618 92060 499546
rect 92478 491464 92534 491473
rect 92478 491399 92480 491408
rect 92532 491399 92534 491408
rect 92480 491370 92532 491376
rect 92584 490657 92612 540138
rect 93228 495038 93256 540138
rect 93872 534818 93900 540138
rect 94516 537470 94544 540138
rect 95787 540110 95832 540138
rect 95148 539164 95200 539170
rect 95148 539106 95200 539112
rect 94504 537464 94556 537470
rect 94504 537406 94556 537412
rect 93860 534812 93912 534818
rect 93860 534754 93912 534760
rect 95056 532024 95108 532030
rect 95056 531966 95108 531972
rect 95068 499574 95096 531966
rect 94976 499546 95096 499574
rect 93216 495032 93268 495038
rect 93216 494974 93268 494980
rect 93216 493400 93268 493406
rect 93216 493342 93268 493348
rect 92848 490680 92900 490686
rect 92570 490648 92626 490657
rect 92020 490612 92072 490618
rect 92848 490622 92900 490628
rect 92570 490583 92626 490592
rect 92020 490554 92072 490560
rect 92860 489954 92888 490622
rect 92598 489926 92888 489954
rect 93228 489940 93256 493342
rect 94976 490521 95004 499546
rect 95160 493626 95188 539106
rect 95804 537606 95832 540110
rect 95792 537600 95844 537606
rect 95792 537542 95844 537548
rect 95240 500268 95292 500274
rect 95240 500210 95292 500216
rect 95252 499574 95280 500210
rect 95252 499546 96016 499574
rect 95068 493598 95188 493626
rect 95068 490754 95096 493598
rect 95148 493468 95200 493474
rect 95148 493410 95200 493416
rect 95056 490748 95108 490754
rect 95056 490690 95108 490696
rect 94134 490512 94190 490521
rect 94134 490447 94190 490456
rect 94962 490512 95018 490521
rect 94962 490447 95018 490456
rect 94148 489954 94176 490447
rect 93886 489926 94176 489954
rect 95160 489940 95188 493410
rect 95790 491872 95846 491881
rect 95790 491807 95846 491816
rect 95804 489940 95832 491807
rect 95988 489954 96016 499546
rect 96448 497486 96476 540138
rect 97092 532166 97120 540138
rect 97080 532160 97132 532166
rect 97080 532102 97132 532108
rect 96436 497480 96488 497486
rect 96436 497422 96488 497428
rect 97736 493542 97764 540138
rect 97908 539096 97960 539102
rect 97908 539038 97960 539044
rect 97816 536172 97868 536178
rect 97816 536114 97868 536120
rect 97724 493536 97776 493542
rect 97724 493478 97776 493484
rect 96988 491972 97040 491978
rect 96988 491914 97040 491920
rect 97000 491745 97028 491914
rect 97828 491745 97856 536114
rect 97920 492046 97948 539038
rect 98380 538218 98408 540138
rect 99024 539578 99052 540138
rect 99012 539572 99064 539578
rect 99012 539514 99064 539520
rect 98644 538960 98696 538966
rect 98644 538902 98696 538908
rect 98368 538212 98420 538218
rect 98368 538154 98420 538160
rect 98380 537674 98408 538154
rect 98368 537668 98420 537674
rect 98368 537610 98420 537616
rect 98552 537532 98604 537538
rect 98552 537474 98604 537480
rect 98564 529145 98592 537474
rect 98550 529136 98606 529145
rect 98550 529071 98606 529080
rect 97908 492040 97960 492046
rect 97908 491982 97960 491988
rect 98368 491972 98420 491978
rect 98368 491914 98420 491920
rect 96986 491736 97042 491745
rect 96986 491671 97042 491680
rect 97814 491736 97870 491745
rect 97814 491671 97870 491680
rect 97446 491192 97502 491201
rect 97446 491127 97502 491136
rect 97460 489954 97488 491127
rect 95988 489926 96416 489954
rect 97106 489926 97488 489954
rect 98380 489940 98408 491914
rect 73436 489874 73488 489880
rect 98656 489870 98684 538902
rect 99024 538898 99052 539514
rect 99012 538892 99064 538898
rect 99012 538834 99064 538840
rect 99668 538214 99696 540138
rect 99392 538186 99696 538214
rect 99288 534880 99340 534886
rect 99288 534822 99340 534828
rect 99300 491337 99328 534822
rect 99286 491328 99342 491337
rect 99286 491263 99342 491272
rect 99300 489954 99328 491263
rect 99038 489926 99328 489954
rect 69020 489864 69072 489870
rect 98000 489864 98052 489870
rect 69020 489806 69072 489812
rect 97750 489812 98000 489818
rect 97750 489806 98052 489812
rect 98644 489864 98696 489870
rect 98644 489806 98696 489812
rect 99196 489864 99248 489870
rect 99196 489806 99248 489812
rect 69032 489025 69060 489806
rect 97750 489790 98040 489806
rect 99208 489258 99236 489806
rect 99196 489252 99248 489258
rect 99196 489194 99248 489200
rect 69018 489016 69074 489025
rect 69018 488951 69074 488960
rect 68926 443864 68982 443873
rect 68926 443799 68982 443808
rect 69032 432614 69060 488951
rect 69846 485888 69902 485897
rect 69846 485823 69902 485832
rect 69860 482633 69888 485823
rect 69846 482624 69902 482633
rect 69846 482559 69902 482568
rect 69202 482488 69258 482497
rect 69860 482458 69888 482559
rect 69202 482423 69258 482432
rect 69848 482452 69900 482458
rect 69112 481636 69164 481642
rect 69112 481578 69164 481584
rect 69124 481545 69152 481578
rect 69110 481536 69166 481545
rect 69110 481471 69166 481480
rect 69020 432608 69072 432614
rect 69020 432550 69072 432556
rect 69124 431118 69152 481471
rect 69216 436966 69244 482423
rect 69848 482394 69900 482400
rect 69662 442232 69718 442241
rect 69662 442167 69718 442176
rect 69676 440065 69704 442167
rect 69754 440736 69810 440745
rect 69810 440694 70058 440722
rect 71056 440706 71346 440722
rect 71044 440700 71346 440706
rect 69754 440671 69810 440680
rect 71096 440694 71346 440700
rect 93886 440706 94176 440722
rect 93886 440700 94188 440706
rect 93886 440694 94136 440700
rect 71044 440642 71096 440648
rect 91744 440632 91796 440638
rect 91744 440574 91796 440580
rect 69662 440056 69718 440065
rect 69662 439991 69718 440000
rect 70398 440056 70454 440065
rect 70454 440014 70702 440042
rect 71792 440014 71990 440042
rect 70398 439991 70454 440000
rect 71792 437594 71820 440014
rect 71700 437566 71820 437594
rect 69204 436960 69256 436966
rect 69204 436902 69256 436908
rect 71700 436762 71728 437566
rect 72424 436960 72476 436966
rect 72424 436902 72476 436908
rect 71688 436756 71740 436762
rect 71688 436698 71740 436704
rect 71872 434648 71924 434654
rect 71872 434590 71924 434596
rect 69664 434036 69716 434042
rect 69664 433978 69716 433984
rect 69112 431112 69164 431118
rect 69112 431054 69164 431060
rect 68926 401432 68982 401441
rect 68982 401390 69244 401418
rect 68926 401367 68982 401376
rect 69216 400246 69244 401390
rect 69204 400240 69256 400246
rect 69204 400182 69256 400188
rect 69112 396024 69164 396030
rect 69112 395966 69164 395972
rect 69124 394738 69152 395966
rect 69112 394732 69164 394738
rect 69112 394674 69164 394680
rect 68928 394664 68980 394670
rect 68928 394606 68980 394612
rect 68940 393378 68968 394606
rect 68928 393372 68980 393378
rect 68928 393314 68980 393320
rect 68940 359514 68968 393314
rect 69124 380769 69152 394674
rect 69216 383489 69244 400182
rect 69296 398132 69348 398138
rect 69296 398074 69348 398080
rect 69308 397526 69336 398074
rect 69296 397520 69348 397526
rect 69296 397462 69348 397468
rect 69202 383480 69258 383489
rect 69202 383415 69258 383424
rect 69110 380760 69166 380769
rect 69110 380695 69166 380704
rect 69216 378826 69244 383415
rect 69204 378820 69256 378826
rect 69204 378762 69256 378768
rect 69308 373994 69336 397462
rect 69676 396030 69704 433978
rect 71884 396846 71912 434590
rect 71964 431112 72016 431118
rect 71964 431054 72016 431060
rect 71976 402974 72004 431054
rect 71976 402946 72096 402974
rect 71872 396840 71924 396846
rect 71872 396782 71924 396788
rect 69664 396024 69716 396030
rect 69664 395966 69716 395972
rect 70400 392624 70452 392630
rect 70400 392566 70452 392572
rect 69572 389904 69624 389910
rect 69572 389846 69624 389852
rect 69584 389434 69612 389846
rect 69572 389428 69624 389434
rect 69572 389370 69624 389376
rect 69584 383654 69612 389370
rect 69756 388612 69808 388618
rect 69756 388554 69808 388560
rect 69768 385914 69796 388554
rect 70412 387870 70440 392566
rect 70400 387864 70452 387870
rect 70400 387806 70452 387812
rect 70412 385914 70440 387806
rect 69768 385886 70058 385914
rect 70412 385886 70702 385914
rect 72068 385778 72096 402946
rect 72436 398886 72464 436902
rect 72620 434654 72648 440028
rect 73160 439544 73212 439550
rect 73160 439486 73212 439492
rect 73172 438802 73200 439486
rect 73160 438796 73212 438802
rect 73160 438738 73212 438744
rect 73264 438258 73292 440028
rect 73344 439136 73396 439142
rect 73344 439078 73396 439084
rect 73252 438252 73304 438258
rect 73252 438194 73304 438200
rect 72608 434648 72660 434654
rect 72608 434590 72660 434596
rect 73356 431954 73384 439078
rect 73908 439074 73936 440028
rect 73896 439068 73948 439074
rect 73896 439010 73948 439016
rect 74552 434722 74580 440028
rect 75840 438734 75868 440028
rect 75828 438728 75880 438734
rect 75828 438670 75880 438676
rect 75184 438320 75236 438326
rect 75184 438262 75236 438268
rect 74540 434716 74592 434722
rect 74540 434658 74592 434664
rect 73264 431926 73384 431954
rect 73264 402974 73292 431926
rect 74630 407552 74686 407561
rect 74630 407487 74686 407496
rect 74540 403028 74592 403034
rect 73264 402946 73384 402974
rect 74540 402970 74592 402976
rect 72424 398880 72476 398886
rect 72424 398822 72476 398828
rect 72436 388074 72464 398822
rect 72424 388068 72476 388074
rect 72424 388010 72476 388016
rect 72436 385914 72464 388010
rect 73356 387938 73384 402946
rect 73344 387932 73396 387938
rect 73344 387874 73396 387880
rect 72436 385886 72634 385914
rect 73356 385778 73384 387874
rect 74552 385948 74580 402970
rect 74506 385920 74580 385948
rect 74644 385948 74672 407487
rect 75196 403034 75224 438262
rect 75274 436792 75330 436801
rect 75274 436727 75330 436736
rect 75288 407561 75316 436727
rect 76010 435840 76066 435849
rect 76010 435775 76066 435784
rect 75274 407552 75330 407561
rect 75274 407487 75330 407496
rect 75288 407153 75316 407487
rect 75274 407144 75330 407153
rect 75274 407079 75330 407088
rect 75920 406292 75972 406298
rect 75920 406234 75972 406240
rect 75184 403028 75236 403034
rect 75184 402970 75236 402976
rect 75368 394120 75420 394126
rect 75368 394062 75420 394068
rect 75380 393446 75408 394062
rect 75368 393440 75420 393446
rect 75368 393382 75420 393388
rect 74644 385920 74856 385948
rect 74506 385914 74534 385920
rect 74828 385914 74856 385920
rect 75380 385914 75408 393382
rect 75932 386050 75960 406234
rect 76024 391338 76052 435775
rect 76484 433294 76512 440028
rect 76564 439612 76616 439618
rect 76564 439554 76616 439560
rect 76472 433288 76524 433294
rect 76472 433230 76524 433236
rect 76576 406298 76604 439554
rect 77128 435849 77156 440028
rect 77496 440014 77786 440042
rect 77496 438705 77524 440014
rect 77482 438696 77538 438705
rect 77482 438631 77538 438640
rect 77114 435840 77170 435849
rect 77114 435775 77170 435784
rect 77390 435296 77446 435305
rect 77390 435231 77446 435240
rect 76564 406292 76616 406298
rect 76564 406234 76616 406240
rect 76576 405822 76604 406234
rect 76564 405816 76616 405822
rect 76564 405758 76616 405764
rect 77404 393314 77432 435231
rect 77312 393286 77432 393314
rect 76012 391332 76064 391338
rect 76012 391274 76064 391280
rect 77312 388890 77340 393286
rect 77300 388884 77352 388890
rect 77300 388826 77352 388832
rect 75932 386022 76696 386050
rect 76668 385914 76696 386022
rect 74506 385886 74566 385914
rect 74828 385886 75210 385914
rect 75380 385886 75854 385914
rect 76668 385886 77142 385914
rect 71792 385750 72096 385778
rect 73278 385750 73384 385778
rect 71792 385354 71820 385750
rect 77496 385393 77524 438631
rect 78416 437374 78444 440028
rect 78784 440014 79074 440042
rect 78404 437368 78456 437374
rect 78404 437310 78456 437316
rect 78416 436490 78444 437310
rect 78404 436484 78456 436490
rect 78404 436426 78456 436432
rect 78784 436082 78812 440014
rect 78772 436076 78824 436082
rect 78772 436018 78824 436024
rect 78678 434616 78734 434625
rect 78678 434551 78734 434560
rect 78692 395418 78720 434551
rect 78680 395412 78732 395418
rect 78680 395354 78732 395360
rect 77576 388884 77628 388890
rect 77576 388826 77628 388832
rect 77588 388006 77616 388826
rect 78220 388476 78272 388482
rect 78220 388418 78272 388424
rect 77576 388000 77628 388006
rect 77576 387942 77628 387948
rect 77588 385914 77616 387942
rect 78232 386442 78260 388418
rect 78784 387122 78812 436018
rect 79704 434625 79732 440028
rect 80716 440014 81006 440042
rect 80716 438666 80744 440014
rect 80704 438660 80756 438666
rect 80704 438602 80756 438608
rect 79690 434616 79746 434625
rect 79690 434551 79746 434560
rect 80716 393990 80744 438602
rect 81636 437238 81664 440028
rect 82280 438802 82308 440028
rect 82268 438796 82320 438802
rect 82268 438738 82320 438744
rect 82924 437306 82952 440028
rect 83568 438870 83596 440028
rect 84226 440014 84608 440042
rect 83556 438864 83608 438870
rect 83556 438806 83608 438812
rect 83556 437980 83608 437986
rect 83556 437922 83608 437928
rect 82912 437300 82964 437306
rect 82912 437242 82964 437248
rect 81624 437232 81676 437238
rect 81624 437174 81676 437180
rect 80796 432608 80848 432614
rect 80796 432550 80848 432556
rect 80808 401674 80836 432550
rect 81636 431954 81664 437174
rect 82924 431954 82952 437242
rect 83464 436484 83516 436490
rect 83464 436426 83516 436432
rect 81544 431926 81664 431954
rect 82832 431926 82952 431954
rect 80796 401668 80848 401674
rect 80796 401610 80848 401616
rect 80704 393984 80756 393990
rect 80704 393926 80756 393932
rect 80808 393314 80836 401610
rect 80532 393286 80836 393314
rect 79324 390584 79376 390590
rect 79324 390526 79376 390532
rect 78772 387116 78824 387122
rect 78772 387058 78824 387064
rect 78220 386436 78272 386442
rect 78220 386378 78272 386384
rect 77588 385886 77786 385914
rect 78232 385778 78260 386378
rect 79336 385914 79364 390526
rect 80060 387864 80112 387870
rect 80060 387806 80112 387812
rect 80072 386073 80100 387806
rect 80532 386510 80560 393286
rect 80612 389360 80664 389366
rect 80612 389302 80664 389308
rect 80520 386504 80572 386510
rect 80520 386446 80572 386452
rect 80058 386064 80114 386073
rect 80058 385999 80114 386008
rect 80532 385914 80560 386446
rect 79336 385886 79718 385914
rect 80362 385886 80560 385914
rect 80624 385914 80652 389302
rect 81440 388544 81492 388550
rect 81440 388486 81492 388492
rect 81452 388074 81480 388486
rect 81440 388068 81492 388074
rect 81440 388010 81492 388016
rect 80624 385886 81006 385914
rect 78232 385750 78430 385778
rect 81544 385762 81572 431926
rect 82832 402974 82860 431926
rect 83476 431254 83504 436426
rect 83464 431248 83516 431254
rect 83464 431190 83516 431196
rect 82832 402946 82952 402974
rect 82820 395344 82872 395350
rect 82820 395286 82872 395292
rect 82832 394806 82860 395286
rect 82820 394800 82872 394806
rect 82820 394742 82872 394748
rect 82924 394058 82952 402946
rect 83004 394800 83056 394806
rect 83004 394742 83056 394748
rect 82912 394052 82964 394058
rect 82912 393994 82964 394000
rect 82820 393508 82872 393514
rect 82820 393450 82872 393456
rect 82832 393310 82860 393450
rect 82820 393304 82872 393310
rect 82820 393246 82872 393252
rect 82360 388068 82412 388074
rect 82360 388010 82412 388016
rect 82372 385778 82400 388010
rect 83016 385914 83044 394742
rect 83096 393508 83148 393514
rect 83096 393450 83148 393456
rect 82938 385886 83044 385914
rect 83108 385914 83136 393450
rect 83476 387190 83504 431190
rect 83568 396778 83596 437922
rect 84580 437345 84608 440014
rect 84856 439074 84884 440028
rect 86158 440014 86264 440042
rect 84844 439068 84896 439074
rect 84844 439010 84896 439016
rect 84856 437986 84884 439010
rect 84844 437980 84896 437986
rect 84844 437922 84896 437928
rect 85580 437436 85632 437442
rect 85580 437378 85632 437384
rect 84566 437336 84622 437345
rect 84566 437271 84622 437280
rect 84580 431954 84608 437271
rect 84580 431926 84884 431954
rect 84856 399634 84884 431926
rect 85488 402280 85540 402286
rect 85488 402222 85540 402228
rect 85500 401713 85528 402222
rect 85118 401704 85174 401713
rect 85118 401639 85174 401648
rect 85486 401704 85542 401713
rect 85486 401639 85542 401648
rect 84844 399628 84896 399634
rect 84844 399570 84896 399576
rect 83556 396772 83608 396778
rect 83556 396714 83608 396720
rect 84476 389428 84528 389434
rect 84476 389370 84528 389376
rect 83464 387184 83516 387190
rect 83464 387126 83516 387132
rect 84488 385914 84516 389370
rect 85132 385914 85160 401639
rect 85592 399566 85620 437378
rect 86236 437374 86264 440014
rect 86788 437442 86816 440028
rect 87432 437481 87460 440028
rect 87708 440014 88090 440042
rect 88734 440014 89024 440042
rect 87418 437472 87474 437481
rect 86776 437436 86828 437442
rect 87418 437407 87474 437416
rect 86776 437378 86828 437384
rect 86224 437368 86276 437374
rect 86224 437310 86276 437316
rect 85670 403608 85726 403617
rect 85670 403543 85726 403552
rect 85684 403073 85712 403543
rect 85670 403064 85726 403073
rect 85670 402999 85726 403008
rect 85580 399560 85632 399566
rect 85580 399502 85632 399508
rect 85684 385914 85712 402999
rect 86236 402974 86264 437310
rect 87432 436529 87460 437407
rect 87708 437238 87736 440014
rect 88996 438870 89024 440014
rect 88984 438864 89036 438870
rect 88984 438806 89036 438812
rect 87696 437232 87748 437238
rect 87696 437174 87748 437180
rect 87418 436520 87474 436529
rect 87418 436455 87474 436464
rect 87708 431954 87736 437174
rect 88246 436520 88302 436529
rect 88246 436455 88302 436464
rect 87616 431926 87736 431954
rect 86236 402946 86356 402974
rect 83108 385886 83582 385914
rect 84488 385886 84870 385914
rect 85132 385886 85514 385914
rect 85684 385886 86158 385914
rect 81532 385756 81584 385762
rect 82294 385750 82400 385778
rect 81532 385698 81584 385704
rect 86328 385694 86356 402946
rect 87512 399492 87564 399498
rect 87512 399434 87564 399440
rect 87524 388362 87552 399434
rect 87616 392698 87644 431926
rect 88260 405113 88288 436455
rect 88246 405104 88302 405113
rect 88246 405039 88302 405048
rect 88248 399492 88300 399498
rect 88248 399434 88300 399440
rect 88260 398954 88288 399434
rect 88248 398948 88300 398954
rect 88248 398890 88300 398896
rect 88340 398132 88392 398138
rect 88340 398074 88392 398080
rect 87604 392692 87656 392698
rect 87604 392634 87656 392640
rect 87524 388334 87736 388362
rect 87052 386572 87104 386578
rect 87052 386514 87104 386520
rect 87064 385914 87092 386514
rect 87708 385914 87736 388334
rect 88352 385914 88380 398074
rect 88996 391270 89024 438806
rect 89364 437782 89392 440028
rect 90008 438802 90036 440028
rect 89996 438796 90048 438802
rect 89996 438738 90048 438744
rect 91008 438796 91060 438802
rect 91008 438738 91060 438744
rect 89352 437776 89404 437782
rect 89352 437718 89404 437724
rect 89718 404968 89774 404977
rect 89718 404903 89774 404912
rect 89732 404433 89760 404903
rect 89718 404424 89774 404433
rect 89718 404359 89774 404368
rect 88984 391264 89036 391270
rect 88984 391206 89036 391212
rect 89732 389366 89760 404359
rect 89812 403640 89864 403646
rect 89812 403582 89864 403588
rect 89720 389360 89772 389366
rect 89720 389302 89772 389308
rect 89824 385914 89852 403582
rect 91020 391950 91048 438738
rect 91296 438190 91324 440028
rect 91652 439204 91704 439210
rect 91652 439146 91704 439152
rect 91664 439006 91692 439146
rect 91652 439000 91704 439006
rect 91652 438942 91704 438948
rect 91284 438184 91336 438190
rect 91284 438126 91336 438132
rect 91756 437782 91784 440574
rect 93964 440042 93992 440694
rect 94136 440642 94188 440648
rect 93886 440028 93992 440042
rect 91940 439210 91968 440028
rect 91928 439204 91980 439210
rect 91928 439146 91980 439152
rect 91940 438938 91968 439146
rect 91928 438932 91980 438938
rect 91928 438874 91980 438880
rect 91744 437776 91796 437782
rect 91744 437718 91796 437724
rect 91008 391944 91060 391950
rect 91008 391886 91060 391892
rect 90364 389360 90416 389366
rect 90364 389302 90416 389308
rect 90376 385914 90404 389302
rect 91560 387864 91612 387870
rect 91560 387806 91612 387812
rect 91572 385914 91600 387806
rect 87064 385886 87446 385914
rect 87708 385886 88090 385914
rect 88352 385886 88734 385914
rect 89824 385886 90022 385914
rect 90376 385886 90666 385914
rect 91310 385886 91600 385914
rect 91756 385694 91784 437718
rect 92584 436082 92612 440028
rect 93228 439249 93256 440028
rect 93872 440014 93992 440028
rect 94530 440014 94912 440042
rect 92846 439240 92902 439249
rect 92846 439175 92902 439184
rect 93214 439240 93270 439249
rect 93214 439175 93270 439184
rect 92572 436076 92624 436082
rect 92572 436018 92624 436024
rect 92860 431954 92888 439175
rect 93872 437474 93900 440014
rect 94044 439000 94096 439006
rect 94044 438942 94096 438948
rect 93780 437446 93900 437474
rect 93676 436076 93728 436082
rect 93676 436018 93728 436024
rect 92492 431926 92888 431954
rect 92492 407833 92520 431926
rect 92478 407824 92534 407833
rect 92478 407759 92534 407768
rect 92664 400988 92716 400994
rect 92664 400930 92716 400936
rect 92572 391944 92624 391950
rect 92572 391886 92624 391892
rect 92584 389978 92612 391886
rect 92572 389972 92624 389978
rect 92572 389914 92624 389920
rect 92676 385778 92704 400930
rect 93688 399537 93716 436018
rect 93674 399528 93730 399537
rect 93674 399463 93730 399472
rect 93780 396778 93808 437446
rect 94056 402286 94084 438942
rect 94884 437374 94912 440014
rect 95160 439006 95188 440028
rect 96448 439074 96476 440028
rect 95240 439068 95292 439074
rect 95240 439010 95292 439016
rect 96436 439068 96488 439074
rect 96436 439010 96488 439016
rect 95148 439000 95200 439006
rect 95148 438942 95200 438948
rect 94872 437368 94924 437374
rect 94872 437310 94924 437316
rect 94884 431954 94912 437310
rect 94884 431926 95188 431954
rect 94044 402280 94096 402286
rect 94044 402222 94096 402228
rect 95160 399498 95188 431926
rect 95148 399492 95200 399498
rect 95148 399434 95200 399440
rect 93768 396772 93820 396778
rect 93768 396714 93820 396720
rect 95252 393990 95280 439010
rect 96448 438938 96476 439010
rect 96618 438968 96674 438977
rect 95884 438932 95936 438938
rect 95884 438874 95936 438880
rect 96436 438932 96488 438938
rect 96618 438903 96674 438912
rect 96436 438874 96488 438880
rect 95896 405074 95924 438874
rect 95884 405068 95936 405074
rect 95884 405010 95936 405016
rect 96632 398041 96660 438903
rect 97092 437306 97120 440028
rect 97736 438977 97764 440028
rect 98090 439240 98146 439249
rect 98090 439175 98146 439184
rect 98104 438977 98132 439175
rect 97722 438968 97778 438977
rect 97722 438903 97778 438912
rect 98090 438968 98146 438977
rect 98090 438903 98146 438912
rect 98380 438598 98408 440028
rect 99024 438734 99052 440028
rect 99392 439793 99420 538186
rect 100312 537538 100340 540138
rect 100300 537532 100352 537538
rect 100300 537474 100352 537480
rect 100760 537464 100812 537470
rect 99470 537432 99526 537441
rect 100760 537406 100812 537412
rect 99470 537367 99526 537376
rect 99484 486713 99512 537367
rect 100772 536722 100800 537406
rect 100956 536897 100984 540138
rect 102227 540110 102272 540138
rect 102244 537810 102272 540110
rect 102232 537804 102284 537810
rect 102232 537746 102284 537752
rect 102888 537742 102916 540138
rect 103532 538218 103560 540138
rect 103520 538212 103572 538218
rect 103520 538154 103572 538160
rect 102876 537736 102928 537742
rect 102876 537678 102928 537684
rect 100942 536888 100998 536897
rect 104176 536858 104204 540138
rect 100942 536823 100998 536832
rect 102048 536852 102100 536858
rect 102048 536794 102100 536800
rect 104164 536852 104216 536858
rect 104164 536794 104216 536800
rect 100760 536716 100812 536722
rect 100760 536658 100812 536664
rect 101404 492040 101456 492046
rect 101404 491982 101456 491988
rect 99656 491564 99708 491570
rect 99656 491506 99708 491512
rect 99668 489940 99696 491506
rect 101218 491464 101274 491473
rect 101218 491399 101274 491408
rect 100024 490748 100076 490754
rect 100024 490690 100076 490696
rect 99470 486704 99526 486713
rect 99470 486639 99526 486648
rect 99484 485858 99512 486639
rect 99472 485852 99524 485858
rect 99472 485794 99524 485800
rect 99378 439784 99434 439793
rect 99378 439719 99434 439728
rect 99012 438728 99064 438734
rect 99012 438670 99064 438676
rect 99288 438728 99340 438734
rect 99288 438670 99340 438676
rect 98368 438592 98420 438598
rect 98368 438534 98420 438540
rect 99196 438592 99248 438598
rect 99196 438534 99248 438540
rect 97080 437300 97132 437306
rect 97080 437242 97132 437248
rect 97092 436422 97120 437242
rect 97080 436416 97132 436422
rect 97080 436358 97132 436364
rect 97908 436416 97960 436422
rect 97908 436358 97960 436364
rect 97920 405006 97948 436358
rect 97908 405000 97960 405006
rect 97908 404942 97960 404948
rect 99208 401062 99236 438534
rect 99196 401056 99248 401062
rect 99196 400998 99248 401004
rect 98000 400920 98052 400926
rect 98000 400862 98052 400868
rect 96618 398032 96674 398041
rect 96618 397967 96674 397976
rect 95976 395412 96028 395418
rect 95976 395354 96028 395360
rect 95240 393984 95292 393990
rect 95240 393926 95292 393932
rect 94136 392624 94188 392630
rect 94136 392566 94188 392572
rect 93308 388000 93360 388006
rect 93308 387942 93360 387948
rect 92598 385750 92704 385778
rect 86316 385688 86368 385694
rect 86316 385630 86368 385636
rect 91744 385688 91796 385694
rect 91744 385630 91796 385636
rect 77482 385384 77538 385393
rect 71780 385348 71832 385354
rect 93320 385370 93348 387942
rect 94148 385914 94176 392566
rect 95884 388272 95936 388278
rect 95884 388214 95936 388220
rect 94872 388136 94924 388142
rect 94872 388078 94924 388084
rect 94884 385914 94912 388078
rect 95896 385914 95924 388214
rect 93886 385886 94176 385914
rect 94530 385886 94912 385914
rect 95818 385886 95924 385914
rect 95988 385914 96016 395354
rect 96712 395344 96764 395350
rect 96712 395286 96764 395292
rect 96724 385914 96752 395286
rect 98012 385914 98040 400862
rect 98552 398200 98604 398206
rect 98552 398142 98604 398148
rect 98564 385914 98592 398142
rect 99300 396846 99328 438670
rect 99668 438190 99696 440028
rect 99656 438184 99708 438190
rect 99656 438126 99708 438132
rect 99380 406836 99432 406842
rect 99380 406778 99432 406784
rect 99392 405754 99420 406778
rect 99380 405748 99432 405754
rect 99380 405690 99432 405696
rect 99288 396840 99340 396846
rect 99288 396782 99340 396788
rect 99392 385914 99420 405690
rect 100036 388822 100064 490690
rect 101232 489870 101260 491399
rect 101220 489864 101272 489870
rect 101220 489806 101272 489812
rect 100114 484528 100170 484537
rect 100114 484463 100170 484472
rect 100128 406842 100156 484463
rect 101232 470594 101260 489806
rect 100956 470566 101260 470594
rect 100208 456204 100260 456210
rect 100208 456146 100260 456152
rect 100220 437442 100248 456146
rect 100668 440292 100720 440298
rect 100668 440234 100720 440240
rect 100680 439793 100708 440234
rect 100666 439784 100722 439793
rect 100666 439719 100722 439728
rect 100208 437436 100260 437442
rect 100208 437378 100260 437384
rect 100760 431316 100812 431322
rect 100760 431258 100812 431264
rect 100772 429894 100800 431258
rect 100760 429888 100812 429894
rect 100760 429830 100812 429836
rect 100116 406836 100168 406842
rect 100116 406778 100168 406784
rect 100956 402974 100984 470566
rect 100956 402946 101076 402974
rect 100024 388816 100076 388822
rect 100024 388758 100076 388764
rect 101048 385914 101076 402946
rect 101416 394058 101444 491982
rect 102060 445874 102088 536794
rect 102140 492720 102192 492726
rect 102140 492662 102192 492668
rect 102048 445868 102100 445874
rect 102048 445810 102100 445816
rect 102048 438184 102100 438190
rect 102048 438126 102100 438132
rect 101404 394052 101456 394058
rect 101404 393994 101456 394000
rect 102060 391270 102088 438126
rect 102152 396642 102180 492662
rect 103612 491700 103664 491706
rect 103612 491642 103664 491648
rect 102232 489320 102284 489326
rect 102230 489288 102232 489297
rect 102284 489288 102286 489297
rect 102230 489223 102286 489232
rect 102324 488504 102376 488510
rect 102324 488446 102376 488452
rect 102232 488096 102284 488102
rect 102336 488073 102364 488446
rect 102232 488038 102284 488044
rect 102322 488064 102378 488073
rect 102244 487937 102272 488038
rect 102322 487999 102378 488008
rect 102230 487928 102286 487937
rect 102230 487863 102286 487872
rect 102232 487144 102284 487150
rect 102232 487086 102284 487092
rect 102244 486713 102272 487086
rect 102230 486704 102286 486713
rect 102230 486639 102286 486648
rect 103518 486432 103574 486441
rect 103518 486367 103574 486376
rect 103426 485752 103482 485761
rect 103532 485738 103560 486367
rect 103482 485710 103560 485738
rect 103426 485687 103482 485696
rect 103426 485208 103482 485217
rect 103426 485143 103482 485152
rect 103440 485110 103468 485143
rect 103428 485104 103480 485110
rect 103428 485046 103480 485052
rect 103426 483848 103482 483857
rect 103426 483783 103482 483792
rect 103440 483682 103468 483783
rect 103428 483676 103480 483682
rect 103428 483618 103480 483624
rect 103334 482624 103390 482633
rect 103334 482559 103390 482568
rect 103348 481778 103376 482559
rect 103426 482488 103482 482497
rect 103426 482423 103482 482432
rect 103440 482322 103468 482423
rect 103428 482316 103480 482322
rect 103428 482258 103480 482264
rect 103336 481772 103388 481778
rect 103336 481714 103388 481720
rect 103428 481636 103480 481642
rect 103428 481578 103480 481584
rect 103336 481568 103388 481574
rect 103440 481545 103468 481578
rect 103336 481510 103388 481516
rect 103426 481536 103482 481545
rect 103348 481273 103376 481510
rect 103426 481471 103482 481480
rect 103334 481264 103390 481273
rect 103334 481199 103390 481208
rect 103426 479904 103482 479913
rect 103426 479839 103482 479848
rect 103334 479768 103390 479777
rect 103334 479703 103390 479712
rect 103348 479602 103376 479703
rect 103336 479596 103388 479602
rect 103336 479538 103388 479544
rect 103440 479534 103468 479839
rect 103428 479528 103480 479534
rect 103428 479470 103480 479476
rect 103426 477728 103482 477737
rect 103426 477663 103482 477672
rect 103440 477562 103468 477663
rect 103428 477556 103480 477562
rect 103428 477498 103480 477504
rect 103242 477048 103298 477057
rect 103242 476983 103298 476992
rect 103256 476066 103284 476983
rect 103336 476876 103388 476882
rect 103336 476818 103388 476824
rect 103348 476513 103376 476818
rect 103334 476504 103390 476513
rect 103334 476439 103390 476448
rect 103244 476060 103296 476066
rect 103244 476002 103296 476008
rect 102232 475992 102284 475998
rect 102232 475934 102284 475940
rect 102244 475697 102272 475934
rect 102324 475924 102376 475930
rect 102324 475866 102376 475872
rect 102230 475688 102286 475697
rect 102230 475623 102286 475632
rect 102336 475153 102364 475866
rect 102322 475144 102378 475153
rect 102322 475079 102378 475088
rect 102232 474700 102284 474706
rect 102232 474642 102284 474648
rect 102244 474337 102272 474642
rect 102230 474328 102286 474337
rect 102230 474263 102286 474272
rect 103256 473354 103284 476002
rect 103426 474736 103482 474745
rect 103426 474671 103482 474680
rect 102232 473340 102284 473346
rect 103256 473326 103376 473354
rect 102232 473282 102284 473288
rect 102244 472977 102272 473282
rect 102230 472968 102286 472977
rect 102230 472903 102286 472912
rect 102232 472660 102284 472666
rect 102232 472602 102284 472608
rect 102244 472297 102272 472602
rect 102230 472288 102286 472297
rect 102230 472223 102286 472232
rect 102324 472048 102376 472054
rect 102324 471990 102376 471996
rect 102230 470928 102286 470937
rect 102230 470863 102286 470872
rect 102244 470626 102272 470863
rect 102336 470665 102364 471990
rect 102322 470656 102378 470665
rect 102232 470620 102284 470626
rect 102322 470591 102378 470600
rect 103348 470594 103376 473326
rect 103440 472054 103468 474671
rect 103428 472048 103480 472054
rect 103428 471990 103480 471996
rect 103624 470594 103652 491642
rect 102232 470562 102284 470568
rect 103348 470566 103468 470594
rect 102230 470248 102286 470257
rect 102230 470183 102286 470192
rect 102244 469946 102272 470183
rect 102232 469940 102284 469946
rect 102232 469882 102284 469888
rect 102230 469568 102286 469577
rect 102230 469503 102286 469512
rect 102244 469266 102272 469503
rect 102232 469260 102284 469266
rect 102232 469202 102284 469208
rect 102230 466984 102286 466993
rect 102230 466919 102286 466928
rect 102244 466546 102272 466919
rect 102232 466540 102284 466546
rect 102232 466482 102284 466488
rect 102324 466404 102376 466410
rect 102324 466346 102376 466352
rect 102230 466168 102286 466177
rect 102230 466103 102286 466112
rect 102244 465730 102272 466103
rect 102232 465724 102284 465730
rect 102232 465666 102284 465672
rect 102336 465633 102364 466346
rect 102322 465624 102378 465633
rect 102322 465559 102378 465568
rect 102232 465044 102284 465050
rect 102232 464986 102284 464992
rect 102244 464817 102272 464986
rect 102230 464808 102286 464817
rect 102230 464743 102286 464752
rect 103334 464264 103390 464273
rect 103334 464199 103390 464208
rect 102232 463684 102284 463690
rect 102232 463626 102284 463632
rect 102244 463457 102272 463626
rect 102230 463448 102286 463457
rect 102230 463383 102286 463392
rect 102232 462324 102284 462330
rect 102232 462266 102284 462272
rect 102244 461553 102272 462266
rect 102322 462088 102378 462097
rect 102322 462023 102378 462032
rect 102230 461544 102286 461553
rect 102230 461479 102286 461488
rect 102336 461038 102364 462023
rect 102324 461032 102376 461038
rect 102324 460974 102376 460980
rect 102232 460896 102284 460902
rect 102232 460838 102284 460844
rect 102244 460193 102272 460838
rect 102414 460728 102470 460737
rect 102414 460663 102470 460672
rect 102324 460216 102376 460222
rect 102230 460184 102286 460193
rect 102324 460158 102376 460164
rect 102230 460119 102286 460128
rect 102230 459368 102286 459377
rect 102230 459303 102286 459312
rect 102244 458930 102272 459303
rect 102232 458924 102284 458930
rect 102232 458866 102284 458872
rect 102336 458833 102364 460158
rect 102428 459610 102456 460663
rect 102416 459604 102468 459610
rect 102416 459546 102468 459552
rect 102322 458824 102378 458833
rect 102322 458759 102378 458768
rect 102232 456748 102284 456754
rect 102232 456690 102284 456696
rect 102244 456113 102272 456690
rect 102322 456648 102378 456657
rect 102322 456583 102378 456592
rect 102336 456142 102364 456583
rect 102324 456136 102376 456142
rect 102230 456104 102286 456113
rect 102324 456078 102376 456084
rect 102230 456039 102286 456048
rect 102324 455388 102376 455394
rect 102324 455330 102376 455336
rect 102232 455320 102284 455326
rect 102230 455288 102232 455297
rect 102284 455288 102286 455297
rect 102230 455223 102286 455232
rect 102336 454753 102364 455330
rect 102322 454744 102378 454753
rect 102322 454679 102378 454688
rect 102232 454028 102284 454034
rect 102232 453970 102284 453976
rect 102244 453937 102272 453970
rect 102324 453960 102376 453966
rect 102230 453928 102286 453937
rect 102324 453902 102376 453908
rect 102230 453863 102286 453872
rect 102336 453393 102364 453902
rect 102322 453384 102378 453393
rect 102322 453319 102378 453328
rect 102232 452600 102284 452606
rect 102230 452568 102232 452577
rect 102284 452568 102286 452577
rect 102230 452503 102286 452512
rect 102784 451308 102836 451314
rect 102784 451250 102836 451256
rect 102230 450664 102286 450673
rect 102230 450599 102286 450608
rect 102244 450294 102272 450599
rect 102796 450537 102824 451250
rect 102782 450528 102838 450537
rect 102782 450463 102838 450472
rect 102232 450288 102284 450294
rect 102232 450230 102284 450236
rect 102232 448724 102284 448730
rect 102232 448666 102284 448672
rect 102244 448633 102272 448666
rect 102230 448624 102286 448633
rect 102230 448559 102286 448568
rect 102232 448520 102284 448526
rect 102230 448488 102232 448497
rect 102284 448488 102286 448497
rect 102230 448423 102286 448432
rect 102324 448452 102376 448458
rect 102324 448394 102376 448400
rect 102336 447953 102364 448394
rect 102322 447944 102378 447953
rect 102322 447879 102378 447888
rect 102322 446584 102378 446593
rect 102322 446519 102378 446528
rect 102336 445806 102364 446519
rect 102416 445868 102468 445874
rect 102416 445810 102468 445816
rect 102324 445800 102376 445806
rect 102230 445768 102286 445777
rect 102324 445742 102376 445748
rect 102230 445703 102232 445712
rect 102284 445703 102286 445712
rect 102232 445674 102284 445680
rect 102428 445233 102456 445810
rect 102414 445224 102470 445233
rect 102414 445159 102470 445168
rect 102232 444032 102284 444038
rect 102232 443974 102284 443980
rect 102244 443873 102272 443974
rect 102230 443864 102286 443873
rect 102230 443799 102286 443808
rect 102230 442504 102286 442513
rect 102230 442439 102286 442448
rect 102244 442270 102272 442439
rect 102232 442264 102284 442270
rect 102232 442206 102284 442212
rect 102232 441584 102284 441590
rect 102232 441526 102284 441532
rect 102244 441153 102272 441526
rect 102230 441144 102286 441153
rect 102230 441079 102286 441088
rect 102140 396636 102192 396642
rect 102140 396578 102192 396584
rect 102784 396636 102836 396642
rect 102784 396578 102836 396584
rect 102152 396098 102180 396578
rect 102140 396092 102192 396098
rect 102140 396034 102192 396040
rect 102048 391264 102100 391270
rect 102048 391206 102100 391212
rect 102138 391232 102194 391241
rect 102138 391167 102194 391176
rect 101404 388816 101456 388822
rect 101404 388758 101456 388764
rect 101416 387841 101444 388758
rect 102152 388278 102180 391167
rect 102600 389904 102652 389910
rect 102600 389846 102652 389852
rect 102140 388272 102192 388278
rect 102140 388214 102192 388220
rect 101402 387832 101458 387841
rect 101402 387767 101458 387776
rect 95988 385886 96462 385914
rect 96724 385886 97106 385914
rect 98012 385886 98394 385914
rect 98564 385886 99038 385914
rect 99392 385886 99682 385914
rect 100970 385886 101352 385914
rect 92952 385354 93348 385370
rect 101324 385354 101352 385886
rect 101416 385778 101444 387767
rect 102612 385914 102640 389846
rect 102796 389162 102824 396578
rect 103348 391338 103376 464199
rect 103440 392601 103468 470566
rect 103532 470566 103652 470594
rect 103426 392592 103482 392601
rect 103426 392527 103482 392536
rect 103336 391332 103388 391338
rect 103336 391274 103388 391280
rect 102784 389156 102836 389162
rect 102784 389098 102836 389104
rect 103532 387870 103560 470566
rect 103612 469872 103664 469878
rect 103612 469814 103664 469820
rect 103624 469033 103652 469814
rect 103610 469024 103666 469033
rect 103610 468959 103666 468968
rect 103612 468512 103664 468518
rect 103612 468454 103664 468460
rect 103624 466857 103652 468454
rect 104164 467152 104216 467158
rect 104164 467094 104216 467100
rect 103610 466848 103666 466857
rect 103610 466783 103666 466792
rect 103612 458856 103664 458862
rect 103612 458798 103664 458804
rect 103624 458153 103652 458798
rect 103610 458144 103666 458153
rect 103610 458079 103666 458088
rect 103610 441960 103666 441969
rect 103610 441895 103666 441904
rect 103624 439074 103652 441895
rect 103612 439068 103664 439074
rect 103612 439010 103664 439016
rect 104176 438666 104204 467094
rect 104716 447160 104768 447166
rect 104716 447102 104768 447108
rect 104164 438660 104216 438666
rect 104164 438602 104216 438608
rect 104728 393314 104756 447102
rect 104820 446162 104848 540138
rect 105648 536897 105676 540382
rect 105634 536888 105690 536897
rect 105634 536823 105690 536832
rect 105740 528554 105768 557506
rect 106922 548856 106978 548865
rect 106922 548791 106978 548800
rect 105910 543824 105966 543833
rect 105910 543759 105966 543768
rect 105556 528526 105768 528554
rect 105176 476808 105228 476814
rect 105174 476776 105176 476785
rect 105228 476776 105230 476785
rect 105174 476711 105230 476720
rect 105556 469946 105584 528526
rect 105636 478916 105688 478922
rect 105636 478858 105688 478864
rect 105544 469940 105596 469946
rect 105544 469882 105596 469888
rect 104992 450288 105044 450294
rect 104992 450230 105044 450236
rect 104820 446134 104940 446162
rect 104912 445738 104940 446134
rect 104900 445732 104952 445738
rect 104900 445674 104952 445680
rect 104808 444440 104860 444446
rect 104808 444382 104860 444388
rect 104820 444038 104848 444382
rect 104808 444032 104860 444038
rect 104808 443974 104860 443980
rect 105004 431322 105032 450230
rect 105544 445732 105596 445738
rect 105544 445674 105596 445680
rect 104992 431316 105044 431322
rect 104992 431258 105044 431264
rect 105004 430642 105032 431258
rect 104992 430636 105044 430642
rect 104992 430578 105044 430584
rect 104636 393286 104756 393314
rect 104532 392692 104584 392698
rect 104532 392634 104584 392640
rect 103612 389156 103664 389162
rect 103612 389098 103664 389104
rect 103520 387864 103572 387870
rect 103520 387806 103572 387812
rect 103624 385914 103652 389098
rect 104440 386572 104492 386578
rect 104440 386514 104492 386520
rect 104452 385914 104480 386514
rect 102258 385886 102640 385914
rect 103546 385886 103652 385914
rect 104190 385886 104480 385914
rect 104544 385778 104572 392634
rect 104636 386578 104664 393286
rect 104808 389156 104860 389162
rect 104808 389098 104860 389104
rect 104820 388278 104848 389098
rect 104808 388272 104860 388278
rect 104808 388214 104860 388220
rect 104808 387864 104860 387870
rect 104808 387806 104860 387812
rect 104820 387190 104848 387806
rect 104808 387184 104860 387190
rect 104808 387126 104860 387132
rect 104624 386572 104676 386578
rect 104624 386514 104676 386520
rect 105556 385801 105584 445674
rect 105648 437238 105676 478858
rect 105924 450294 105952 543759
rect 106278 540696 106334 540705
rect 106278 540631 106334 540640
rect 106292 536790 106320 540631
rect 106280 536784 106332 536790
rect 106280 536726 106332 536732
rect 106292 536110 106320 536726
rect 106280 536104 106332 536110
rect 106280 536046 106332 536052
rect 106188 489184 106240 489190
rect 106188 489126 106240 489132
rect 106200 488102 106228 489126
rect 106188 488096 106240 488102
rect 106188 488038 106240 488044
rect 106280 481840 106332 481846
rect 106280 481782 106332 481788
rect 106292 481574 106320 481782
rect 106280 481568 106332 481574
rect 106280 481510 106332 481516
rect 106188 469192 106240 469198
rect 106188 469134 106240 469140
rect 106096 456068 106148 456074
rect 106096 456010 106148 456016
rect 106108 455326 106136 456010
rect 106096 455320 106148 455326
rect 106096 455262 106148 455268
rect 105912 450288 105964 450294
rect 105912 450230 105964 450236
rect 105636 437232 105688 437238
rect 105636 437174 105688 437180
rect 106200 402354 106228 469134
rect 106936 456754 106964 548791
rect 107028 481846 107056 572727
rect 108946 571976 109002 571985
rect 108946 571911 109002 571920
rect 107658 571432 107714 571441
rect 108960 571402 108988 571911
rect 107658 571367 107714 571376
rect 108948 571396 109000 571402
rect 107476 540932 107528 540938
rect 107476 540874 107528 540880
rect 107488 540161 107516 540874
rect 107474 540152 107530 540161
rect 107474 540087 107530 540096
rect 107016 481840 107068 481846
rect 107016 481782 107068 481788
rect 106924 456748 106976 456754
rect 106924 456690 106976 456696
rect 107384 454708 107436 454714
rect 107384 454650 107436 454656
rect 107396 453966 107424 454650
rect 107384 453960 107436 453966
rect 107384 453902 107436 453908
rect 106278 451344 106334 451353
rect 106278 451279 106334 451288
rect 106292 449993 106320 451279
rect 107488 451274 107516 540087
rect 107568 491292 107620 491298
rect 107568 491234 107620 491240
rect 107580 490686 107608 491234
rect 107568 490680 107620 490686
rect 107568 490622 107620 490628
rect 107396 451246 107516 451274
rect 106278 449984 106334 449993
rect 106278 449919 106334 449928
rect 106832 448724 106884 448730
rect 106832 448666 106884 448672
rect 106844 447846 106872 448666
rect 107396 448662 107424 451246
rect 107384 448656 107436 448662
rect 107384 448598 107436 448604
rect 107396 448458 107424 448598
rect 107384 448452 107436 448458
rect 107384 448394 107436 448400
rect 106832 447840 106884 447846
rect 106832 447782 106884 447788
rect 106924 439068 106976 439074
rect 106924 439010 106976 439016
rect 106188 402348 106240 402354
rect 106188 402290 106240 402296
rect 106936 396030 106964 439010
rect 106924 396024 106976 396030
rect 106924 395966 106976 395972
rect 106280 394052 106332 394058
rect 106280 393994 106332 394000
rect 106292 392086 106320 393994
rect 106280 392080 106332 392086
rect 106280 392022 106332 392028
rect 106188 387864 106240 387870
rect 106188 387806 106240 387812
rect 106200 385914 106228 387806
rect 106122 385886 106228 385914
rect 106292 385914 106320 392022
rect 107580 386646 107608 490622
rect 107672 479602 107700 571367
rect 108948 571338 109000 571344
rect 108854 570616 108910 570625
rect 108854 570551 108910 570560
rect 108868 569974 108896 570551
rect 108946 570072 109002 570081
rect 108946 570007 108948 570016
rect 109000 570007 109002 570016
rect 108948 569978 109000 569984
rect 108856 569968 108908 569974
rect 108856 569910 108908 569916
rect 108946 569256 109002 569265
rect 108946 569191 109002 569200
rect 108960 568614 108988 569191
rect 108948 568608 109000 568614
rect 108948 568550 109000 568556
rect 108854 567896 108910 567905
rect 108854 567831 108910 567840
rect 108868 567254 108896 567831
rect 108946 567352 109002 567361
rect 108946 567287 108948 567296
rect 109000 567287 109002 567296
rect 108948 567258 109000 567264
rect 108856 567248 108908 567254
rect 108856 567190 108908 567196
rect 108394 566536 108450 566545
rect 108394 566471 108450 566480
rect 108408 565894 108436 566471
rect 108946 565992 109002 566001
rect 108946 565927 108948 565936
rect 109000 565927 109002 565936
rect 108948 565898 109000 565904
rect 108396 565888 108448 565894
rect 108396 565830 108448 565836
rect 108854 565176 108910 565185
rect 108854 565111 108910 565120
rect 108868 564466 108896 565111
rect 108948 564528 109000 564534
rect 108946 564496 108948 564505
rect 109000 564496 109002 564505
rect 108856 564460 108908 564466
rect 108946 564431 109002 564440
rect 108856 564402 108908 564408
rect 108948 564392 109000 564398
rect 108948 564334 109000 564340
rect 108960 563961 108988 564334
rect 108946 563952 109002 563961
rect 108946 563887 109002 563896
rect 108946 561096 109002 561105
rect 108946 561031 109002 561040
rect 108210 560416 108266 560425
rect 108960 560386 108988 561031
rect 108210 560351 108266 560360
rect 108948 560380 109000 560386
rect 108224 560318 108252 560351
rect 108948 560322 109000 560328
rect 108212 560312 108264 560318
rect 108212 560254 108264 560260
rect 108854 559736 108910 559745
rect 108854 559671 108910 559680
rect 108868 558958 108896 559671
rect 108946 559056 109002 559065
rect 108946 558991 108948 559000
rect 109000 558991 109002 559000
rect 108948 558962 109000 558968
rect 108856 558952 108908 558958
rect 108856 558894 108908 558900
rect 108946 558376 109002 558385
rect 108946 558311 109002 558320
rect 108302 557696 108358 557705
rect 108302 557631 108358 557640
rect 107842 551576 107898 551585
rect 107842 551511 107844 551520
rect 107896 551511 107898 551520
rect 107844 551482 107896 551488
rect 107660 479596 107712 479602
rect 107660 479538 107712 479544
rect 108316 466410 108344 557631
rect 108960 557598 108988 558311
rect 108948 557592 109000 557598
rect 108948 557534 109000 557540
rect 108946 557016 109002 557025
rect 108946 556951 109002 556960
rect 108960 556578 108988 556951
rect 108948 556572 109000 556578
rect 108948 556514 109000 556520
rect 108948 556164 109000 556170
rect 108948 556106 109000 556112
rect 108960 555801 108988 556106
rect 108946 555792 109002 555801
rect 108946 555727 109002 555736
rect 108854 554296 108910 554305
rect 108854 554231 108910 554240
rect 108868 553518 108896 554231
rect 108946 553616 109002 553625
rect 108946 553551 109002 553560
rect 108856 553512 108908 553518
rect 108856 553454 108908 553460
rect 108960 553450 108988 553551
rect 108948 553444 109000 553450
rect 108948 553386 109000 553392
rect 108946 552936 109002 552945
rect 108946 552871 109002 552880
rect 108394 552256 108450 552265
rect 108394 552191 108450 552200
rect 108304 466404 108356 466410
rect 108304 466346 108356 466352
rect 108304 464364 108356 464370
rect 108304 464306 108356 464312
rect 108316 442270 108344 464306
rect 108408 460902 108436 552191
rect 108960 552090 108988 552871
rect 108948 552084 109000 552090
rect 108948 552026 109000 552032
rect 108946 550896 109002 550905
rect 108946 550831 109002 550840
rect 108960 550662 108988 550831
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108854 550216 108910 550225
rect 108854 550151 108910 550160
rect 108868 549302 108896 550151
rect 108946 549536 109002 549545
rect 108946 549471 109002 549480
rect 108960 549370 108988 549471
rect 108948 549364 109000 549370
rect 108948 549306 109000 549312
rect 108856 549296 108908 549302
rect 108856 549238 108908 549244
rect 108946 547496 109002 547505
rect 108946 547431 109002 547440
rect 108486 546816 108542 546825
rect 108486 546751 108542 546760
rect 108396 460896 108448 460902
rect 108396 460838 108448 460844
rect 108396 460284 108448 460290
rect 108396 460226 108448 460232
rect 108408 459610 108436 460226
rect 108396 459604 108448 459610
rect 108396 459546 108448 459552
rect 108500 458250 108528 546751
rect 108960 546514 108988 547431
rect 108948 546508 109000 546514
rect 108948 546450 109000 546456
rect 108946 546136 109002 546145
rect 108946 546071 109002 546080
rect 108960 545766 108988 546071
rect 108948 545760 109000 545766
rect 108948 545702 109000 545708
rect 108946 545456 109002 545465
rect 108946 545391 109002 545400
rect 108960 545154 108988 545391
rect 108948 545148 109000 545154
rect 108948 545090 109000 545096
rect 108856 545080 108908 545086
rect 108856 545022 108908 545028
rect 108868 544921 108896 545022
rect 108854 544912 108910 544921
rect 108854 544847 108910 544856
rect 108946 543416 109002 543425
rect 108946 543351 109002 543360
rect 108960 542434 108988 543351
rect 108948 542428 109000 542434
rect 108948 542370 109000 542376
rect 108946 542056 109002 542065
rect 108946 541991 109002 542000
rect 108960 541006 108988 541991
rect 108948 541000 109000 541006
rect 108948 540942 109000 540948
rect 109052 491298 109080 585414
rect 109130 580136 109186 580145
rect 109130 580071 109186 580080
rect 109040 491292 109092 491298
rect 109040 491234 109092 491240
rect 109144 488510 109172 580071
rect 109696 540938 109724 703122
rect 115204 703112 115256 703118
rect 115204 703054 115256 703060
rect 111708 702908 111760 702914
rect 111708 702850 111760 702856
rect 110696 585404 110748 585410
rect 110696 585346 110748 585352
rect 110512 582684 110564 582690
rect 110512 582626 110564 582632
rect 110420 545216 110472 545222
rect 110420 545158 110472 545164
rect 110432 545086 110460 545158
rect 110420 545080 110472 545086
rect 110420 545022 110472 545028
rect 109776 541068 109828 541074
rect 109776 541010 109828 541016
rect 109684 540932 109736 540938
rect 109684 540874 109736 540880
rect 109788 538218 109816 541010
rect 109776 538212 109828 538218
rect 109776 538154 109828 538160
rect 110524 536178 110552 582626
rect 110604 572008 110656 572014
rect 110604 571950 110656 571956
rect 110616 556170 110644 571950
rect 110604 556164 110656 556170
rect 110604 556106 110656 556112
rect 110616 555490 110644 556106
rect 110604 555484 110656 555490
rect 110604 555426 110656 555432
rect 110604 551540 110656 551546
rect 110604 551482 110656 551488
rect 110512 536172 110564 536178
rect 110512 536114 110564 536120
rect 109224 532092 109276 532098
rect 109224 532034 109276 532040
rect 109132 488504 109184 488510
rect 109132 488446 109184 488452
rect 109144 487830 109172 488446
rect 109132 487824 109184 487830
rect 109132 487766 109184 487772
rect 109236 478922 109264 532034
rect 110616 529242 110644 551482
rect 110420 529236 110472 529242
rect 110420 529178 110472 529184
rect 110604 529236 110656 529242
rect 110604 529178 110656 529184
rect 110432 528630 110460 529178
rect 110420 528624 110472 528630
rect 110420 528566 110472 528572
rect 109316 497616 109368 497622
rect 109316 497558 109368 497564
rect 109224 478916 109276 478922
rect 109224 478858 109276 478864
rect 108948 477488 109000 477494
rect 108948 477430 109000 477436
rect 108856 459604 108908 459610
rect 108856 459546 108908 459552
rect 108488 458244 108540 458250
rect 108488 458186 108540 458192
rect 108500 455394 108528 458186
rect 108488 455388 108540 455394
rect 108488 455330 108540 455336
rect 108304 442264 108356 442270
rect 108304 442206 108356 442212
rect 108316 394058 108344 442206
rect 108868 396914 108896 459546
rect 108960 399673 108988 477430
rect 109328 456210 109356 497558
rect 110420 497548 110472 497554
rect 110420 497490 110472 497496
rect 109408 490612 109460 490618
rect 109408 490554 109460 490560
rect 109316 456204 109368 456210
rect 109316 456146 109368 456152
rect 109420 436082 109448 490554
rect 110328 481772 110380 481778
rect 110328 481714 110380 481720
rect 110340 481574 110368 481714
rect 110328 481568 110380 481574
rect 110328 481510 110380 481516
rect 109408 436076 109460 436082
rect 109408 436018 109460 436024
rect 108946 399664 109002 399673
rect 108946 399599 109002 399608
rect 108856 396908 108908 396914
rect 108856 396850 108908 396856
rect 108304 394052 108356 394058
rect 108304 393994 108356 394000
rect 110340 389881 110368 481510
rect 110432 439142 110460 497490
rect 110708 493610 110736 585346
rect 111720 545222 111748 702850
rect 113088 702704 113140 702710
rect 113088 702646 113140 702652
rect 112076 584452 112128 584458
rect 112076 584394 112128 584400
rect 111984 584044 112036 584050
rect 111984 583986 112036 583992
rect 111892 565888 111944 565894
rect 111892 565830 111944 565836
rect 111708 545216 111760 545222
rect 111708 545158 111760 545164
rect 110788 537804 110840 537810
rect 110788 537746 110840 537752
rect 110512 493604 110564 493610
rect 110512 493546 110564 493552
rect 110696 493604 110748 493610
rect 110696 493546 110748 493552
rect 110524 493338 110552 493546
rect 110512 493332 110564 493338
rect 110512 493274 110564 493280
rect 110604 491496 110656 491502
rect 110604 491438 110656 491444
rect 110616 447166 110644 491438
rect 110800 464370 110828 537746
rect 111800 498840 111852 498846
rect 111800 498782 111852 498788
rect 111062 491328 111118 491337
rect 111062 491263 111118 491272
rect 110788 464364 110840 464370
rect 110788 464306 110840 464312
rect 110604 447160 110656 447166
rect 110604 447102 110656 447108
rect 110420 439136 110472 439142
rect 110420 439078 110472 439084
rect 110880 392828 110932 392834
rect 110880 392770 110932 392776
rect 110892 392154 110920 392770
rect 110880 392148 110932 392154
rect 110880 392090 110932 392096
rect 109038 389872 109094 389881
rect 109038 389807 109040 389816
rect 109092 389807 109094 389816
rect 110326 389872 110382 389881
rect 110326 389807 110382 389816
rect 109040 389778 109092 389784
rect 110328 389360 110380 389366
rect 110328 389302 110380 389308
rect 109130 388920 109186 388929
rect 109130 388855 109186 388864
rect 109144 388210 109172 388855
rect 109132 388204 109184 388210
rect 109132 388146 109184 388152
rect 109040 388136 109092 388142
rect 109040 388078 109092 388084
rect 108948 387932 109000 387938
rect 108948 387874 109000 387880
rect 107568 386640 107620 386646
rect 107568 386582 107620 386588
rect 107580 385914 107608 386582
rect 108960 385914 108988 387874
rect 109052 386374 109080 388078
rect 109040 386368 109092 386374
rect 109040 386310 109092 386316
rect 106292 385886 106766 385914
rect 107410 385886 107608 385914
rect 108698 385886 108988 385914
rect 105542 385792 105598 385801
rect 101416 385750 101614 385778
rect 104544 385750 104834 385778
rect 109144 385778 109172 388146
rect 110340 385914 110368 389302
rect 109986 385886 110368 385914
rect 110892 385914 110920 392090
rect 111076 390114 111104 491263
rect 111706 459640 111762 459649
rect 111706 459575 111762 459584
rect 111156 430636 111208 430642
rect 111156 430578 111208 430584
rect 111064 390108 111116 390114
rect 111064 390050 111116 390056
rect 111168 387122 111196 430578
rect 111720 400994 111748 459575
rect 111812 440638 111840 498782
rect 111904 475930 111932 565830
rect 111996 494902 112024 583986
rect 112088 499574 112116 584394
rect 113100 545766 113128 702646
rect 113364 586832 113416 586838
rect 113364 586774 113416 586780
rect 113272 583976 113324 583982
rect 113272 583918 113324 583924
rect 113180 565956 113232 565962
rect 113180 565898 113232 565904
rect 113088 545760 113140 545766
rect 113088 545702 113140 545708
rect 112088 499546 112484 499574
rect 112168 495032 112220 495038
rect 112168 494974 112220 494980
rect 111984 494896 112036 494902
rect 111984 494838 112036 494844
rect 111984 485104 112036 485110
rect 111982 485072 111984 485081
rect 112036 485072 112038 485081
rect 111982 485007 112038 485016
rect 111892 475924 111944 475930
rect 111892 475866 111944 475872
rect 112180 440978 112208 494974
rect 112456 491201 112484 499546
rect 112442 491192 112498 491201
rect 112442 491127 112498 491136
rect 112168 440972 112220 440978
rect 112168 440914 112220 440920
rect 111800 440632 111852 440638
rect 111800 440574 111852 440580
rect 111708 400988 111760 400994
rect 111708 400930 111760 400936
rect 112456 393314 112484 491127
rect 112628 475924 112680 475930
rect 112628 475866 112680 475872
rect 112640 475386 112668 475866
rect 112628 475380 112680 475386
rect 112628 475322 112680 475328
rect 113192 474706 113220 565898
rect 113284 493474 113312 583918
rect 113376 539102 113404 586774
rect 114560 583772 114612 583778
rect 114560 583714 114612 583720
rect 113916 556572 113968 556578
rect 113916 556514 113968 556520
rect 113364 539096 113416 539102
rect 113364 539038 113416 539044
rect 113272 493468 113324 493474
rect 113272 493410 113324 493416
rect 113272 491632 113324 491638
rect 113272 491574 113324 491580
rect 113180 474700 113232 474706
rect 113180 474642 113232 474648
rect 113180 422340 113232 422346
rect 113180 422282 113232 422288
rect 113192 421598 113220 422282
rect 113180 421592 113232 421598
rect 113180 421534 113232 421540
rect 113284 403646 113312 491574
rect 113824 489252 113876 489258
rect 113824 489194 113876 489200
rect 113272 403640 113324 403646
rect 113272 403582 113324 403588
rect 113836 402974 113864 489194
rect 113928 465118 113956 556514
rect 114572 491570 114600 583714
rect 114652 581188 114704 581194
rect 114652 581130 114704 581136
rect 114664 534886 114692 581130
rect 115216 538214 115244 703054
rect 117228 702772 117280 702778
rect 117228 702714 117280 702720
rect 116032 582616 116084 582622
rect 116032 582558 116084 582564
rect 115940 557592 115992 557598
rect 115940 557534 115992 557540
rect 114848 538186 115244 538214
rect 114848 538121 114876 538186
rect 114834 538112 114890 538121
rect 114834 538047 114890 538056
rect 114652 534880 114704 534886
rect 114652 534822 114704 534828
rect 114744 493536 114796 493542
rect 114744 493478 114796 493484
rect 114560 491564 114612 491570
rect 114560 491506 114612 491512
rect 114558 482352 114614 482361
rect 114558 482287 114560 482296
rect 114612 482287 114614 482296
rect 114560 482258 114612 482264
rect 113916 465112 113968 465118
rect 113916 465054 113968 465060
rect 114756 438598 114784 493478
rect 114848 467158 114876 538047
rect 115204 534880 115256 534886
rect 115204 534822 115256 534828
rect 115216 489326 115244 534822
rect 115204 489320 115256 489326
rect 115204 489262 115256 489268
rect 115216 483002 115244 489262
rect 115204 482996 115256 483002
rect 115204 482938 115256 482944
rect 115204 479596 115256 479602
rect 115204 479538 115256 479544
rect 114836 467152 114888 467158
rect 114836 467094 114888 467100
rect 114744 438592 114796 438598
rect 114744 438534 114796 438540
rect 115216 402974 115244 479538
rect 115480 474700 115532 474706
rect 115480 474642 115532 474648
rect 113836 402946 113956 402974
rect 115216 402946 115336 402974
rect 112364 393286 112484 393314
rect 112168 388136 112220 388142
rect 112168 388078 112220 388084
rect 111800 387864 111852 387870
rect 111800 387806 111852 387812
rect 111156 387116 111208 387122
rect 111156 387058 111208 387064
rect 111812 387025 111840 387806
rect 111798 387016 111854 387025
rect 111798 386951 111854 386960
rect 112180 385914 112208 388078
rect 112364 386617 112392 393286
rect 113928 390726 113956 402946
rect 114284 392760 114336 392766
rect 114284 392702 114336 392708
rect 113916 390720 113968 390726
rect 113916 390662 113968 390668
rect 112350 386608 112406 386617
rect 112350 386543 112406 386552
rect 110892 385886 111274 385914
rect 111918 385886 112208 385914
rect 112364 385778 112392 386543
rect 113928 385914 113956 390662
rect 113850 385886 113956 385914
rect 114296 385778 114324 392702
rect 114928 390108 114980 390114
rect 114928 390050 114980 390056
rect 114940 387870 114968 390050
rect 114928 387864 114980 387870
rect 114928 387806 114980 387812
rect 114940 385778 114968 387806
rect 109144 385750 109342 385778
rect 112364 385750 112562 385778
rect 114296 385750 114494 385778
rect 114940 385750 115138 385778
rect 105542 385727 105598 385736
rect 77482 385319 77538 385328
rect 92940 385348 93348 385354
rect 71780 385290 71832 385296
rect 92992 385342 93348 385348
rect 101312 385348 101364 385354
rect 92940 385290 92992 385296
rect 101312 385290 101364 385296
rect 69032 373966 69336 373994
rect 69400 383626 69612 383654
rect 69032 364410 69060 373966
rect 69296 371204 69348 371210
rect 69296 371146 69348 371152
rect 69308 370161 69336 371146
rect 69294 370152 69350 370161
rect 69294 370087 69350 370096
rect 69020 364404 69072 364410
rect 69020 364346 69072 364352
rect 69032 363633 69060 364346
rect 69018 363624 69074 363633
rect 69018 363559 69074 363568
rect 69110 360632 69166 360641
rect 69110 360567 69166 360576
rect 68928 359508 68980 359514
rect 68928 359450 68980 359456
rect 68836 346384 68888 346390
rect 68834 346352 68836 346361
rect 68888 346352 68890 346361
rect 68834 346287 68890 346296
rect 68744 329112 68796 329118
rect 68744 329054 68796 329060
rect 67456 319660 67508 319666
rect 67456 319602 67508 319608
rect 69124 302326 69152 360567
rect 69308 354674 69336 370087
rect 69400 363730 69428 383626
rect 69662 380760 69718 380769
rect 69662 380695 69718 380704
rect 69676 379574 69704 380695
rect 115308 380322 115336 402946
rect 115492 383654 115520 474642
rect 115952 465730 115980 557534
rect 116044 495514 116072 582558
rect 117240 564398 117268 702714
rect 137284 700460 137336 700466
rect 137284 700402 137336 700408
rect 126244 616888 126296 616894
rect 126244 616830 126296 616836
rect 118884 588600 118936 588606
rect 118884 588542 118936 588548
rect 117320 586696 117372 586702
rect 117320 586638 117372 586644
rect 117228 564392 117280 564398
rect 117228 564334 117280 564340
rect 117240 563718 117268 564334
rect 117228 563712 117280 563718
rect 117228 563654 117280 563660
rect 116124 560380 116176 560386
rect 116124 560322 116176 560328
rect 116032 495508 116084 495514
rect 116032 495450 116084 495456
rect 116032 487824 116084 487830
rect 116032 487766 116084 487772
rect 115940 465724 115992 465730
rect 115940 465666 115992 465672
rect 115940 461032 115992 461038
rect 115940 460974 115992 460980
rect 115952 460902 115980 460974
rect 115940 460896 115992 460902
rect 115940 460838 115992 460844
rect 115848 389496 115900 389502
rect 115848 389438 115900 389444
rect 115754 387968 115810 387977
rect 115754 387903 115756 387912
rect 115808 387903 115810 387912
rect 115756 387874 115808 387880
rect 115860 385914 115888 389438
rect 115782 385886 115888 385914
rect 115492 383626 115612 383654
rect 115296 380316 115348 380322
rect 115296 380258 115348 380264
rect 69664 379568 69716 379574
rect 69664 379510 69716 379516
rect 69848 379432 69900 379438
rect 69848 379374 69900 379380
rect 69860 378321 69888 379374
rect 69478 378312 69534 378321
rect 69478 378247 69534 378256
rect 69846 378312 69902 378321
rect 69846 378247 69902 378256
rect 69388 363724 69440 363730
rect 69388 363666 69440 363672
rect 69216 354646 69336 354674
rect 69216 340202 69244 354646
rect 69204 340196 69256 340202
rect 69204 340138 69256 340144
rect 69492 316810 69520 378247
rect 115478 376408 115534 376417
rect 115478 376343 115534 376352
rect 115492 371929 115520 376343
rect 115478 371920 115534 371929
rect 115478 371855 115534 371864
rect 115584 367713 115612 383626
rect 115570 367704 115626 367713
rect 115570 367639 115626 367648
rect 115294 364848 115350 364857
rect 115294 364783 115350 364792
rect 115308 345014 115336 364783
rect 115308 344986 115428 345014
rect 69754 340096 69810 340105
rect 69810 340068 70058 340082
rect 69810 340054 70072 340068
rect 69754 340031 69810 340040
rect 70044 337550 70072 340054
rect 70400 339652 70452 339658
rect 70400 339594 70452 339600
rect 70032 337544 70084 337550
rect 70032 337486 70084 337492
rect 70412 322250 70440 339594
rect 70688 339590 70716 340068
rect 71332 339658 71360 340068
rect 71320 339652 71372 339658
rect 71320 339594 71372 339600
rect 70492 339584 70544 339590
rect 70492 339526 70544 339532
rect 70676 339584 70728 339590
rect 70676 339526 70728 339532
rect 70504 327826 70532 339526
rect 71976 336462 72004 340068
rect 73218 339930 73246 340068
rect 73068 339924 73120 339930
rect 73068 339866 73120 339872
rect 73206 339924 73258 339930
rect 73206 339866 73258 339872
rect 71964 336456 72016 336462
rect 71964 336398 72016 336404
rect 72424 336456 72476 336462
rect 72424 336398 72476 336404
rect 70492 327820 70544 327826
rect 70492 327762 70544 327768
rect 71780 325032 71832 325038
rect 71780 324974 71832 324980
rect 70400 322244 70452 322250
rect 70400 322186 70452 322192
rect 69480 316804 69532 316810
rect 69480 316746 69532 316752
rect 70400 306536 70452 306542
rect 70400 306478 70452 306484
rect 69204 303680 69256 303686
rect 69204 303622 69256 303628
rect 69112 302320 69164 302326
rect 69112 302262 69164 302268
rect 68836 301368 68888 301374
rect 68836 301310 68888 301316
rect 68848 300898 68876 301310
rect 68836 300892 68888 300898
rect 68836 300834 68888 300840
rect 67546 298208 67602 298217
rect 67546 298143 67602 298152
rect 67560 297566 67588 298143
rect 67548 297560 67600 297566
rect 67548 297502 67600 297508
rect 68744 292596 68796 292602
rect 68744 292538 68796 292544
rect 67640 291168 67692 291174
rect 67640 291110 67692 291116
rect 67652 290873 67680 291110
rect 67638 290864 67694 290873
rect 67638 290799 67694 290808
rect 67638 289912 67694 289921
rect 67638 289847 67640 289856
rect 67692 289847 67694 289856
rect 67640 289818 67692 289824
rect 67454 288552 67510 288561
rect 67454 288487 67510 288496
rect 67362 246392 67418 246401
rect 67362 246327 67418 246336
rect 67376 245546 67404 246327
rect 67364 245540 67416 245546
rect 67364 245482 67416 245488
rect 67362 244352 67418 244361
rect 67362 244287 67418 244296
rect 67376 235278 67404 244287
rect 67364 235272 67416 235278
rect 67364 235214 67416 235220
rect 67468 224262 67496 288487
rect 67638 287192 67694 287201
rect 67638 287127 67694 287136
rect 67652 287094 67680 287127
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67822 287056 67878 287065
rect 67732 287020 67784 287026
rect 67822 286991 67878 287000
rect 67732 286962 67784 286968
rect 67744 286793 67772 286962
rect 67730 286784 67786 286793
rect 67730 286719 67786 286728
rect 67836 285734 67864 286991
rect 68192 286340 68244 286346
rect 68192 286282 68244 286288
rect 68204 286113 68232 286282
rect 68190 286104 68246 286113
rect 68190 286039 68246 286048
rect 67824 285728 67876 285734
rect 67824 285670 67876 285676
rect 67640 285660 67692 285666
rect 67640 285602 67692 285608
rect 67652 285433 67680 285602
rect 67638 285424 67694 285433
rect 67638 285359 67694 285368
rect 67638 284472 67694 284481
rect 67638 284407 67694 284416
rect 67652 284374 67680 284407
rect 67640 284368 67692 284374
rect 67640 284310 67692 284316
rect 67732 284300 67784 284306
rect 67732 284242 67784 284248
rect 67744 283393 67772 284242
rect 67730 283384 67786 283393
rect 67730 283319 67786 283328
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 282169 67680 282814
rect 67638 282160 67694 282169
rect 67638 282095 67694 282104
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67640 280084 67692 280090
rect 67640 280026 67692 280032
rect 67652 279313 67680 280026
rect 67744 279993 67772 280094
rect 67730 279984 67786 279993
rect 67730 279919 67786 279928
rect 67638 279304 67694 279313
rect 67638 279239 67694 279248
rect 67640 278724 67692 278730
rect 67640 278666 67692 278672
rect 67652 278633 67680 278666
rect 67638 278624 67694 278633
rect 67638 278559 67694 278568
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277438 67680 277607
rect 67640 277432 67692 277438
rect 67640 277374 67692 277380
rect 67730 276448 67786 276457
rect 67730 276383 67786 276392
rect 67744 276078 67772 276383
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 67640 276004 67692 276010
rect 67640 275946 67692 275952
rect 67652 275913 67680 275946
rect 67638 275904 67694 275913
rect 67638 275839 67694 275848
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274718 67680 274887
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 67732 274644 67784 274650
rect 67732 274586 67784 274592
rect 67744 274553 67772 274586
rect 67730 274544 67786 274553
rect 67730 274479 67786 274488
rect 67638 273592 67694 273601
rect 67638 273527 67694 273536
rect 67652 273290 67680 273527
rect 67640 273284 67692 273290
rect 67640 273226 67692 273232
rect 67638 272368 67694 272377
rect 67638 272303 67694 272312
rect 67652 271930 67680 272303
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67744 271153 67772 271798
rect 68098 271552 68154 271561
rect 68098 271487 68154 271496
rect 67730 271144 67786 271153
rect 67730 271079 67786 271088
rect 68112 270570 68140 271487
rect 68100 270564 68152 270570
rect 68100 270506 68152 270512
rect 67638 269648 67694 269657
rect 67638 269583 67694 269592
rect 67652 269142 67680 269583
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67640 268388 67692 268394
rect 67640 268330 67692 268336
rect 67652 268161 67680 268330
rect 67638 268152 67694 268161
rect 67638 268087 67694 268096
rect 67732 267708 67784 267714
rect 67732 267650 67784 267656
rect 67638 267064 67694 267073
rect 67638 266999 67640 267008
rect 67692 266999 67694 267008
rect 67640 266970 67692 266976
rect 67744 266937 67772 267650
rect 67730 266928 67786 266937
rect 67730 266863 67786 266872
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265713 67680 266290
rect 68756 266257 68784 292538
rect 68848 288153 68876 300834
rect 68928 295452 68980 295458
rect 68928 295394 68980 295400
rect 68834 288144 68890 288153
rect 68834 288079 68890 288088
rect 68834 272232 68890 272241
rect 68834 272167 68890 272176
rect 68742 266248 68798 266257
rect 68742 266183 68798 266192
rect 67638 265704 67694 265713
rect 67638 265639 67694 265648
rect 67730 264208 67786 264217
rect 67730 264143 67786 264152
rect 67640 263696 67692 263702
rect 67638 263664 67640 263673
rect 67692 263664 67694 263673
rect 67744 263634 67772 264143
rect 67638 263599 67694 263608
rect 67732 263628 67784 263634
rect 68848 263594 68876 272167
rect 67732 263570 67784 263576
rect 68756 263566 68876 263594
rect 67640 263560 67692 263566
rect 67638 263528 67640 263537
rect 67692 263528 67694 263537
rect 67638 263463 67694 263472
rect 67638 262304 67694 262313
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67824 262200 67876 262206
rect 67824 262142 67876 262148
rect 67730 261488 67786 261497
rect 67730 261423 67786 261432
rect 67744 260914 67772 261423
rect 67836 261361 67864 262142
rect 67822 261352 67878 261361
rect 67822 261287 67878 261296
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 258632 67694 258641
rect 67638 258567 67694 258576
rect 67652 258194 67680 258567
rect 67730 258224 67786 258233
rect 67640 258188 67692 258194
rect 67730 258159 67786 258168
rect 67640 258130 67692 258136
rect 67744 258126 67772 258159
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257961 67680 257994
rect 67638 257952 67694 257961
rect 67638 257887 67694 257896
rect 67638 256864 67694 256873
rect 67638 256799 67694 256808
rect 67652 256766 67680 256799
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 68756 256034 68784 263566
rect 68756 256006 68876 256034
rect 68742 255912 68798 255921
rect 68742 255847 68798 255856
rect 67638 255368 67694 255377
rect 67638 255303 67640 255312
rect 67692 255303 67694 255312
rect 67640 255274 67692 255280
rect 67732 255264 67784 255270
rect 67638 255232 67694 255241
rect 67732 255206 67784 255212
rect 67638 255167 67640 255176
rect 67692 255167 67694 255176
rect 67640 255138 67692 255144
rect 67744 254833 67772 255206
rect 67730 254824 67786 254833
rect 67730 254759 67786 254768
rect 67640 253904 67692 253910
rect 67638 253872 67640 253881
rect 67692 253872 67694 253881
rect 67638 253807 67694 253816
rect 67732 253836 67784 253842
rect 67732 253778 67784 253784
rect 67744 253473 67772 253778
rect 67730 253464 67786 253473
rect 67730 253399 67786 253408
rect 67640 251184 67692 251190
rect 67638 251152 67640 251161
rect 67692 251152 67694 251161
rect 67638 251087 67694 251096
rect 68558 249928 68614 249937
rect 68558 249863 68614 249872
rect 67638 249112 67694 249121
rect 67638 249047 67694 249056
rect 67652 248470 67680 249047
rect 68374 248704 68430 248713
rect 68374 248639 68430 248648
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67638 247752 67694 247761
rect 67638 247687 67694 247696
rect 67652 247110 67680 247687
rect 67640 247104 67692 247110
rect 67640 247046 67692 247052
rect 67546 245712 67602 245721
rect 67546 245647 67602 245656
rect 67560 238066 67588 245647
rect 67640 245608 67692 245614
rect 67640 245550 67692 245556
rect 67652 245313 67680 245550
rect 67638 245304 67694 245313
rect 67638 245239 67694 245248
rect 67732 244248 67784 244254
rect 67732 244190 67784 244196
rect 67640 244180 67692 244186
rect 67640 244122 67692 244128
rect 67652 243817 67680 244122
rect 67638 243808 67694 243817
rect 67638 243743 67694 243752
rect 67744 243681 67772 244190
rect 67730 243672 67786 243681
rect 67730 243607 67786 243616
rect 68388 238754 68416 248639
rect 68572 243574 68600 249863
rect 68560 243568 68612 243574
rect 68560 243510 68612 243516
rect 68388 238726 68692 238754
rect 67548 238060 67600 238066
rect 67548 238002 67600 238008
rect 68664 236706 68692 238726
rect 68652 236700 68704 236706
rect 68652 236642 68704 236648
rect 67456 224256 67508 224262
rect 67456 224198 67508 224204
rect 68756 222970 68784 255847
rect 68848 231169 68876 256006
rect 68940 251433 68968 295394
rect 69112 295384 69164 295390
rect 69112 295326 69164 295332
rect 69020 289196 69072 289202
rect 69020 289138 69072 289144
rect 68926 251424 68982 251433
rect 68926 251359 68982 251368
rect 68928 243568 68980 243574
rect 68928 243510 68980 243516
rect 68834 231160 68890 231169
rect 68834 231095 68890 231104
rect 68744 222964 68796 222970
rect 68744 222906 68796 222912
rect 68940 198121 68968 243510
rect 68926 198112 68982 198121
rect 68926 198047 68982 198056
rect 69032 186969 69060 289138
rect 69124 281353 69152 295326
rect 69110 281344 69166 281353
rect 69110 281279 69166 281288
rect 69110 268288 69166 268297
rect 69110 268223 69166 268232
rect 69124 191214 69152 268223
rect 69216 260273 69244 303622
rect 69480 302320 69532 302326
rect 69480 302262 69532 302268
rect 69492 301510 69520 302262
rect 69480 301504 69532 301510
rect 69480 301446 69532 301452
rect 70412 291977 70440 306478
rect 71320 295316 71372 295322
rect 71320 295258 71372 295264
rect 70412 291949 70702 291977
rect 71332 291963 71360 295258
rect 71688 292528 71740 292534
rect 71688 292470 71740 292476
rect 71700 292369 71728 292470
rect 71686 292360 71742 292369
rect 71686 292295 71742 292304
rect 71792 291977 71820 324974
rect 72436 311166 72464 336398
rect 72424 311160 72476 311166
rect 72424 311102 72476 311108
rect 73080 307154 73108 339866
rect 73908 339386 73936 340068
rect 73896 339380 73948 339386
rect 73896 339322 73948 339328
rect 73908 335354 73936 339322
rect 74552 337958 74580 340068
rect 75840 339425 75868 340068
rect 76500 339810 76528 340068
rect 76500 339782 76604 339810
rect 75826 339416 75882 339425
rect 75826 339351 75882 339360
rect 74540 337952 74592 337958
rect 74540 337894 74592 337900
rect 75276 337952 75328 337958
rect 75276 337894 75328 337900
rect 73816 335326 73936 335354
rect 73160 323604 73212 323610
rect 73160 323546 73212 323552
rect 73068 307148 73120 307154
rect 73068 307090 73120 307096
rect 72608 294772 72660 294778
rect 72608 294714 72660 294720
rect 71792 291949 71990 291977
rect 72620 291963 72648 294714
rect 73172 291977 73200 323546
rect 73816 308514 73844 335326
rect 74632 332648 74684 332654
rect 74632 332590 74684 332596
rect 73896 309188 73948 309194
rect 73896 309130 73948 309136
rect 73804 308508 73856 308514
rect 73804 308450 73856 308456
rect 73908 296002 73936 309130
rect 73896 295996 73948 296002
rect 73896 295938 73948 295944
rect 74644 294370 74672 332590
rect 75184 319524 75236 319530
rect 75184 319466 75236 319472
rect 75196 295322 75224 319466
rect 75288 315994 75316 337894
rect 75840 336802 75868 339351
rect 75828 336796 75880 336802
rect 75828 336738 75880 336744
rect 76576 336530 76604 339782
rect 76564 336524 76616 336530
rect 76564 336466 76616 336472
rect 75920 335164 75972 335170
rect 75920 335106 75972 335112
rect 75932 334422 75960 335106
rect 75920 334416 75972 334422
rect 75920 334358 75972 334364
rect 75276 315988 75328 315994
rect 75276 315930 75328 315936
rect 75276 298172 75328 298178
rect 75276 298114 75328 298120
rect 75184 295316 75236 295322
rect 75184 295258 75236 295264
rect 74632 294364 74684 294370
rect 74632 294306 74684 294312
rect 74540 294160 74592 294166
rect 74540 294102 74592 294108
rect 73896 292732 73948 292738
rect 73896 292674 73948 292680
rect 73172 291949 73278 291977
rect 73908 291963 73936 292674
rect 74552 291963 74580 294102
rect 75288 291977 75316 298114
rect 75460 294364 75512 294370
rect 75460 294306 75512 294312
rect 75210 291949 75316 291977
rect 75472 291938 75500 294306
rect 75932 293282 75960 334358
rect 76472 296744 76524 296750
rect 76472 296686 76524 296692
rect 75920 293276 75972 293282
rect 75920 293218 75972 293224
rect 76484 291963 76512 296686
rect 76576 296041 76604 336466
rect 77128 334422 77156 340068
rect 77298 338736 77354 338745
rect 77298 338671 77354 338680
rect 77116 334416 77168 334422
rect 77116 334358 77168 334364
rect 76562 296032 76618 296041
rect 76562 295967 76618 295976
rect 77312 294370 77340 338671
rect 77390 336016 77446 336025
rect 77390 335951 77446 335960
rect 77300 294364 77352 294370
rect 77300 294306 77352 294312
rect 77116 294296 77168 294302
rect 77116 294238 77168 294244
rect 77128 291963 77156 294238
rect 77404 291977 77432 335951
rect 78416 332586 78444 340068
rect 79076 339810 79104 340068
rect 79076 339782 79364 339810
rect 79336 337929 79364 339782
rect 79704 339318 79732 340068
rect 80946 339810 80974 340068
rect 80716 339782 80974 339810
rect 79692 339312 79744 339318
rect 79692 339254 79744 339260
rect 79704 338230 79732 339254
rect 79692 338224 79744 338230
rect 79692 338166 79744 338172
rect 79322 337920 79378 337929
rect 79322 337855 79378 337864
rect 78404 332580 78456 332586
rect 78404 332522 78456 332528
rect 78416 331294 78444 332522
rect 77944 331288 77996 331294
rect 77944 331230 77996 331236
rect 78404 331288 78456 331294
rect 78404 331230 78456 331236
rect 77956 320958 77984 331230
rect 77944 320952 77996 320958
rect 77944 320894 77996 320900
rect 79336 305726 79364 337855
rect 80716 335238 80744 339782
rect 80704 335232 80756 335238
rect 80704 335174 80756 335180
rect 80716 316742 80744 335174
rect 81636 333946 81664 340068
rect 82280 337482 82308 340068
rect 83464 338224 83516 338230
rect 83464 338166 83516 338172
rect 82268 337476 82320 337482
rect 82268 337418 82320 337424
rect 81624 333940 81676 333946
rect 81624 333882 81676 333888
rect 81636 332722 81664 333882
rect 81624 332716 81676 332722
rect 81624 332658 81676 332664
rect 82084 332716 82136 332722
rect 82084 332658 82136 332664
rect 80704 316736 80756 316742
rect 80704 316678 80756 316684
rect 79416 315308 79468 315314
rect 79416 315250 79468 315256
rect 79324 305720 79376 305726
rect 79324 305662 79376 305668
rect 79324 302932 79376 302938
rect 79324 302874 79376 302880
rect 78036 294364 78088 294370
rect 78036 294306 78088 294312
rect 77404 291949 77786 291977
rect 78048 291938 78076 294306
rect 79336 294302 79364 302874
rect 79324 294296 79376 294302
rect 79324 294238 79376 294244
rect 79428 294030 79456 315250
rect 82096 314090 82124 332658
rect 82084 314084 82136 314090
rect 82084 314026 82136 314032
rect 81440 312588 81492 312594
rect 81440 312530 81492 312536
rect 80336 295316 80388 295322
rect 80336 295258 80388 295264
rect 79692 294092 79744 294098
rect 79692 294034 79744 294040
rect 79416 294024 79468 294030
rect 79416 293966 79468 293972
rect 79428 291977 79456 293966
rect 79074 291949 79456 291977
rect 79704 291963 79732 294034
rect 80348 291963 80376 295258
rect 80980 292800 81032 292806
rect 80980 292742 81032 292748
rect 80992 291963 81020 292742
rect 81452 291977 81480 312530
rect 82820 299736 82872 299742
rect 82820 299678 82872 299684
rect 81900 299600 81952 299606
rect 81900 299542 81952 299548
rect 81452 291949 81650 291977
rect 81912 291938 81940 299542
rect 82832 291977 82860 299678
rect 83476 298790 83504 338166
rect 83568 333810 83596 340068
rect 84212 337414 84240 340068
rect 84856 339114 84884 340068
rect 84844 339108 84896 339114
rect 84844 339050 84896 339056
rect 84200 337408 84252 337414
rect 84200 337350 84252 337356
rect 84856 335102 84884 339050
rect 86144 337890 86172 340068
rect 86742 339810 86770 340068
rect 86420 339782 86770 339810
rect 86132 337884 86184 337890
rect 86132 337826 86184 337832
rect 86420 336598 86448 339782
rect 87432 339386 87460 340068
rect 87420 339380 87472 339386
rect 87420 339322 87472 339328
rect 87604 339380 87656 339386
rect 87604 339322 87656 339328
rect 86868 337884 86920 337890
rect 86868 337826 86920 337832
rect 86880 337414 86908 337826
rect 86868 337408 86920 337414
rect 86868 337350 86920 337356
rect 86408 336592 86460 336598
rect 86408 336534 86460 336540
rect 86224 336116 86276 336122
rect 86224 336058 86276 336064
rect 84844 335096 84896 335102
rect 84844 335038 84896 335044
rect 83556 333804 83608 333810
rect 83556 333746 83608 333752
rect 83568 308446 83596 333746
rect 84292 329248 84344 329254
rect 84292 329190 84344 329196
rect 83556 308440 83608 308446
rect 83556 308382 83608 308388
rect 83464 298784 83516 298790
rect 83464 298726 83516 298732
rect 83556 296880 83608 296886
rect 83556 296822 83608 296828
rect 82832 291949 82938 291977
rect 83568 291963 83596 296822
rect 84200 294024 84252 294030
rect 84200 293966 84252 293972
rect 84212 291963 84240 293966
rect 84304 291938 84332 329190
rect 84384 318164 84436 318170
rect 84384 318106 84436 318112
rect 84396 306374 84424 318106
rect 85580 307080 85632 307086
rect 85580 307022 85632 307028
rect 84396 306346 84976 306374
rect 84948 291977 84976 306346
rect 85592 294386 85620 307022
rect 86236 295322 86264 336058
rect 86316 327956 86368 327962
rect 86316 327898 86368 327904
rect 86328 306374 86356 327898
rect 86420 320793 86448 336534
rect 87616 333878 87644 339322
rect 88720 335306 88748 340068
rect 89318 339810 89346 340068
rect 89088 339782 89346 339810
rect 89088 336666 89116 339782
rect 90008 337793 90036 340068
rect 91008 338836 91060 338842
rect 91008 338778 91060 338784
rect 89994 337784 90050 337793
rect 89994 337719 90050 337728
rect 90914 337784 90970 337793
rect 90914 337719 90970 337728
rect 89076 336660 89128 336666
rect 89076 336602 89128 336608
rect 88708 335300 88760 335306
rect 88708 335242 88760 335248
rect 88720 334014 88748 335242
rect 88708 334008 88760 334014
rect 88708 333950 88760 333956
rect 87604 333872 87656 333878
rect 87604 333814 87656 333820
rect 88340 327752 88392 327758
rect 88340 327694 88392 327700
rect 86406 320784 86462 320793
rect 86406 320719 86462 320728
rect 87604 306468 87656 306474
rect 87604 306410 87656 306416
rect 86328 306346 86448 306374
rect 86224 295316 86276 295322
rect 86224 295258 86276 295264
rect 85592 294358 86264 294386
rect 86132 294296 86184 294302
rect 86132 294238 86184 294244
rect 84948 291949 85514 291977
rect 86144 291963 86172 294238
rect 86236 291977 86264 294358
rect 86420 292534 86448 306346
rect 86960 302320 87012 302326
rect 86960 302262 87012 302268
rect 86408 292528 86460 292534
rect 86408 292470 86460 292476
rect 86236 291949 86802 291977
rect 86972 291938 87000 302262
rect 87616 294302 87644 306410
rect 88352 306374 88380 327694
rect 88984 326392 89036 326398
rect 88984 326334 89036 326340
rect 88996 306374 89024 326334
rect 89088 309806 89116 336602
rect 89168 334008 89220 334014
rect 89168 333950 89220 333956
rect 89180 323678 89208 333950
rect 89168 323672 89220 323678
rect 89168 323614 89220 323620
rect 90928 314022 90956 337719
rect 90916 314016 90968 314022
rect 90916 313958 90968 313964
rect 89720 310616 89772 310622
rect 89720 310558 89772 310564
rect 89076 309800 89128 309806
rect 89076 309742 89128 309748
rect 88352 306346 88932 306374
rect 88996 306346 89116 306374
rect 87696 301572 87748 301578
rect 87696 301514 87748 301520
rect 87708 294778 87736 301514
rect 87696 294772 87748 294778
rect 87696 294714 87748 294720
rect 88708 294772 88760 294778
rect 88708 294714 88760 294720
rect 88064 294636 88116 294642
rect 88064 294578 88116 294584
rect 87604 294296 87656 294302
rect 87604 294238 87656 294244
rect 88076 291963 88104 294578
rect 88720 291963 88748 294714
rect 88904 291977 88932 306346
rect 89088 292126 89116 306346
rect 89076 292120 89128 292126
rect 89076 292062 89128 292068
rect 89732 291977 89760 310558
rect 91020 305794 91048 338778
rect 91296 338026 91324 340068
rect 91940 338842 91968 340068
rect 91928 338836 91980 338842
rect 91928 338778 91980 338784
rect 91284 338020 91336 338026
rect 91284 337962 91336 337968
rect 91744 338020 91796 338026
rect 91744 337962 91796 337968
rect 91100 336864 91152 336870
rect 91100 336806 91152 336812
rect 91112 336734 91140 336806
rect 91100 336728 91152 336734
rect 91100 336670 91152 336676
rect 91008 305788 91060 305794
rect 91008 305730 91060 305736
rect 91756 304366 91784 337962
rect 92584 335306 92612 340068
rect 92572 335300 92624 335306
rect 92572 335242 92624 335248
rect 93228 331226 93256 340068
rect 94516 336870 94544 340068
rect 94504 336864 94556 336870
rect 94504 336806 94556 336812
rect 93768 335300 93820 335306
rect 93768 335242 93820 335248
rect 93216 331220 93268 331226
rect 93216 331162 93268 331168
rect 93124 326596 93176 326602
rect 93124 326538 93176 326544
rect 91744 304360 91796 304366
rect 91744 304302 91796 304308
rect 91282 297392 91338 297401
rect 91282 297327 91338 297336
rect 91296 296857 91324 297327
rect 91282 296848 91338 296857
rect 90640 296812 90692 296818
rect 91282 296783 91338 296792
rect 90640 296754 90692 296760
rect 88904 291949 89378 291977
rect 89732 291949 90022 291977
rect 90652 291963 90680 296754
rect 91296 291963 91324 296783
rect 93136 296714 93164 326538
rect 93780 301646 93808 335242
rect 95160 333946 95188 340068
rect 95148 333940 95200 333946
rect 95148 333882 95200 333888
rect 95160 330698 95188 333882
rect 95804 330721 95832 340068
rect 97092 334558 97120 340068
rect 97736 339182 97764 340068
rect 97724 339176 97776 339182
rect 97724 339118 97776 339124
rect 97908 339176 97960 339182
rect 97908 339118 97960 339124
rect 97264 336796 97316 336802
rect 97264 336738 97316 336744
rect 97080 334552 97132 334558
rect 97080 334494 97132 334500
rect 96526 331120 96582 331129
rect 96526 331055 96582 331064
rect 96540 330721 96568 331055
rect 95068 330670 95188 330698
rect 95790 330712 95846 330721
rect 95068 330614 95096 330670
rect 95790 330647 95846 330656
rect 96526 330712 96582 330721
rect 96526 330647 96582 330656
rect 95056 330608 95108 330614
rect 95056 330550 95108 330556
rect 95148 330608 95200 330614
rect 95148 330550 95200 330556
rect 93952 316872 94004 316878
rect 93952 316814 94004 316820
rect 93964 306374 93992 316814
rect 93964 306346 94636 306374
rect 93768 301640 93820 301646
rect 93768 301582 93820 301588
rect 94504 299124 94556 299130
rect 94504 299066 94556 299072
rect 94516 298382 94544 299066
rect 94504 298376 94556 298382
rect 94504 298318 94556 298324
rect 92952 296686 93164 296714
rect 92952 292874 92980 296686
rect 93216 292936 93268 292942
rect 93216 292878 93268 292884
rect 92572 292868 92624 292874
rect 92572 292810 92624 292816
rect 92940 292868 92992 292874
rect 92940 292810 92992 292816
rect 92584 291963 92612 292810
rect 93228 291963 93256 292878
rect 93860 292868 93912 292874
rect 93860 292810 93912 292816
rect 93872 291963 93900 292810
rect 94516 291963 94544 298318
rect 94608 291938 94636 306346
rect 95160 299130 95188 330550
rect 95332 319456 95384 319462
rect 95332 319398 95384 319404
rect 95148 299124 95200 299130
rect 95148 299066 95200 299072
rect 95344 291977 95372 319398
rect 96540 308582 96568 330647
rect 96620 324964 96672 324970
rect 96620 324906 96672 324912
rect 96528 308576 96580 308582
rect 96528 308518 96580 308524
rect 96632 306374 96660 324906
rect 97276 312662 97304 336738
rect 97816 335096 97868 335102
rect 97816 335038 97868 335044
rect 97828 334558 97856 335038
rect 97816 334552 97868 334558
rect 97816 334494 97868 334500
rect 97264 312656 97316 312662
rect 97264 312598 97316 312604
rect 97828 311234 97856 334494
rect 97816 311228 97868 311234
rect 97816 311170 97868 311176
rect 96632 306346 97396 306374
rect 97080 297424 97132 297430
rect 97080 297366 97132 297372
rect 96436 292664 96488 292670
rect 97092 292641 97120 297366
rect 96436 292606 96488 292612
rect 97078 292632 97134 292641
rect 95344 291949 95818 291977
rect 96448 291963 96476 292606
rect 97078 292567 97134 292576
rect 97092 291963 97120 292567
rect 97368 291938 97396 306346
rect 97920 297430 97948 339118
rect 98380 335238 98408 340068
rect 98644 338904 98696 338910
rect 98644 338846 98696 338852
rect 98368 335232 98420 335238
rect 98368 335174 98420 335180
rect 98656 306374 98684 338846
rect 99286 338192 99342 338201
rect 99286 338127 99342 338136
rect 98656 306346 98776 306374
rect 98552 300688 98604 300694
rect 98552 300630 98604 300636
rect 97908 297424 97960 297430
rect 97908 297366 97960 297372
rect 98368 292664 98420 292670
rect 98368 292606 98420 292612
rect 98380 291963 98408 292606
rect 98564 291938 98592 300630
rect 98748 292670 98776 306346
rect 99300 303074 99328 338127
rect 99668 337754 99696 340068
rect 99656 337748 99708 337754
rect 99656 337690 99708 337696
rect 100312 336734 100340 340068
rect 100668 337748 100720 337754
rect 100668 337690 100720 337696
rect 100300 336728 100352 336734
rect 100300 336670 100352 336676
rect 99288 303068 99340 303074
rect 99288 303010 99340 303016
rect 99656 298308 99708 298314
rect 99656 298250 99708 298256
rect 98736 292664 98788 292670
rect 98736 292606 98788 292612
rect 99668 291963 99696 298250
rect 100680 296954 100708 337690
rect 100956 333878 100984 340068
rect 102244 339289 102272 340068
rect 102230 339280 102286 339289
rect 102230 339215 102286 339224
rect 102244 338201 102272 339215
rect 102230 338192 102286 338201
rect 102230 338127 102286 338136
rect 101404 337544 101456 337550
rect 101404 337486 101456 337492
rect 100944 333872 100996 333878
rect 100944 333814 100996 333820
rect 101416 301714 101444 337486
rect 102888 337482 102916 340068
rect 103532 338094 103560 340068
rect 104820 339318 104848 340068
rect 104808 339312 104860 339318
rect 104808 339254 104860 339260
rect 104820 338774 104848 339254
rect 104808 338768 104860 338774
rect 104808 338710 104860 338716
rect 103520 338088 103572 338094
rect 103520 338030 103572 338036
rect 101956 337476 102008 337482
rect 101956 337418 102008 337424
rect 102876 337476 102928 337482
rect 102876 337418 102928 337424
rect 101968 317422 101996 337418
rect 102048 333872 102100 333878
rect 102048 333814 102100 333820
rect 101956 317416 102008 317422
rect 101956 317358 102008 317364
rect 102060 305658 102088 333814
rect 104900 332036 104952 332042
rect 104900 331978 104952 331984
rect 103520 329180 103572 329186
rect 103520 329122 103572 329128
rect 102784 314696 102836 314702
rect 102784 314638 102836 314644
rect 102048 305652 102100 305658
rect 102048 305594 102100 305600
rect 101404 301708 101456 301714
rect 101404 301650 101456 301656
rect 102140 300960 102192 300966
rect 102140 300902 102192 300908
rect 100760 300076 100812 300082
rect 100760 300018 100812 300024
rect 101220 300076 101272 300082
rect 101220 300018 101272 300024
rect 100772 299674 100800 300018
rect 100760 299668 100812 299674
rect 100760 299610 100812 299616
rect 100668 296948 100720 296954
rect 100668 296890 100720 296896
rect 100944 295656 100996 295662
rect 100944 295598 100996 295604
rect 100956 291963 100984 295598
rect 101232 291938 101260 300018
rect 102152 291977 102180 300902
rect 102796 300694 102824 314638
rect 102784 300688 102836 300694
rect 102784 300630 102836 300636
rect 102152 291949 102258 291977
rect 103532 291963 103560 329122
rect 104808 296948 104860 296954
rect 104808 296890 104860 296896
rect 104162 294536 104218 294545
rect 104162 294471 104218 294480
rect 104176 291963 104204 294471
rect 104820 291963 104848 296890
rect 104912 294370 104940 331978
rect 105464 314634 105492 340068
rect 106124 339810 106152 340068
rect 106124 339782 106228 339810
rect 106200 336666 106228 339782
rect 106924 339516 106976 339522
rect 106924 339458 106976 339464
rect 106188 336660 106240 336666
rect 106188 336602 106240 336608
rect 106200 325106 106228 336602
rect 106936 326534 106964 339458
rect 107396 332586 107424 340068
rect 107568 337340 107620 337346
rect 107568 337282 107620 337288
rect 107384 332580 107436 332586
rect 107384 332522 107436 332528
rect 107476 327140 107528 327146
rect 107476 327082 107528 327088
rect 106924 326528 106976 326534
rect 106924 326470 106976 326476
rect 106188 325100 106240 325106
rect 106188 325042 106240 325048
rect 107108 316804 107160 316810
rect 107108 316746 107160 316752
rect 105452 314628 105504 314634
rect 105452 314570 105504 314576
rect 107120 310486 107148 316746
rect 107108 310480 107160 310486
rect 107108 310422 107160 310428
rect 104992 300212 105044 300218
rect 104992 300154 105044 300160
rect 104900 294364 104952 294370
rect 104900 294306 104952 294312
rect 103150 291952 103206 291961
rect 75472 291910 75842 291938
rect 78048 291910 78418 291938
rect 81912 291910 82282 291938
rect 84304 291910 84858 291938
rect 86972 291910 87434 291938
rect 92296 291916 92348 291922
rect 91954 291864 92296 291870
rect 94608 291910 95162 291938
rect 97368 291910 97738 291938
rect 98564 291910 99026 291938
rect 101232 291910 101602 291938
rect 102902 291910 103150 291938
rect 105004 291938 105032 300154
rect 107488 296714 107516 327082
rect 107396 296686 107516 296714
rect 107396 295361 107424 296686
rect 107580 295882 107608 337282
rect 108040 335170 108068 340068
rect 108028 335164 108080 335170
rect 108028 335106 108080 335112
rect 108040 331906 108068 335106
rect 108028 331900 108080 331906
rect 108028 331842 108080 331848
rect 107658 331800 107714 331809
rect 107658 331735 107714 331744
rect 107672 306374 107700 331735
rect 108684 327078 108712 340068
rect 109972 337822 110000 340068
rect 110616 339046 110644 340068
rect 110604 339040 110656 339046
rect 110604 338982 110656 338988
rect 111260 337929 111288 340068
rect 111708 339040 111760 339046
rect 111708 338982 111760 338988
rect 111246 337920 111302 337929
rect 111246 337855 111302 337864
rect 111614 337920 111670 337929
rect 111614 337855 111670 337864
rect 109960 337816 110012 337822
rect 109960 337758 110012 337764
rect 108672 327072 108724 327078
rect 108672 327014 108724 327020
rect 108684 319530 108712 327014
rect 108672 319524 108724 319530
rect 108672 319466 108724 319472
rect 111064 319524 111116 319530
rect 111064 319466 111116 319472
rect 107672 306346 108436 306374
rect 107488 295854 107608 295882
rect 107382 295352 107438 295361
rect 107382 295287 107438 295296
rect 106740 294840 106792 294846
rect 106740 294782 106792 294788
rect 105820 294364 105872 294370
rect 105820 294306 105872 294312
rect 105832 291977 105860 294306
rect 105832 291949 106122 291977
rect 106752 291963 106780 294782
rect 107396 291963 107424 295287
rect 107488 293185 107516 295854
rect 107568 295724 107620 295730
rect 107568 295666 107620 295672
rect 107580 294642 107608 295666
rect 107568 294636 107620 294642
rect 107568 294578 107620 294584
rect 108028 294636 108080 294642
rect 108028 294578 108080 294584
rect 107474 293176 107530 293185
rect 107474 293111 107530 293120
rect 108040 291963 108068 294578
rect 108408 291977 108436 306346
rect 109684 299668 109736 299674
rect 109684 299610 109736 299616
rect 109316 294908 109368 294914
rect 109316 294850 109368 294856
rect 108408 291949 108698 291977
rect 109328 291963 109356 294850
rect 109696 291977 109724 299610
rect 111076 294914 111104 319466
rect 111628 316810 111656 337855
rect 111616 316804 111668 316810
rect 111616 316746 111668 316752
rect 111156 305040 111208 305046
rect 111156 304982 111208 304988
rect 111064 294908 111116 294914
rect 111064 294850 111116 294856
rect 111168 294710 111196 304982
rect 111720 298858 111748 338982
rect 111800 327888 111852 327894
rect 111800 327830 111852 327836
rect 111708 298852 111760 298858
rect 111708 298794 111760 298800
rect 111248 294908 111300 294914
rect 111248 294850 111300 294856
rect 111156 294704 111208 294710
rect 111156 294646 111208 294652
rect 110604 294092 110656 294098
rect 110604 294034 110656 294040
rect 109696 291949 109986 291977
rect 110616 291963 110644 294034
rect 111260 291963 111288 294850
rect 111812 291977 111840 327830
rect 112548 318782 112576 340068
rect 113192 339454 113220 340068
rect 113180 339448 113232 339454
rect 113180 339390 113232 339396
rect 113836 336598 113864 340068
rect 115138 340054 115244 340082
rect 115110 339552 115166 339561
rect 115110 339487 115166 339496
rect 113916 339448 113968 339454
rect 113916 339390 113968 339396
rect 113824 336592 113876 336598
rect 113824 336534 113876 336540
rect 113836 330614 113864 336534
rect 113824 330608 113876 330614
rect 113824 330550 113876 330556
rect 113824 325100 113876 325106
rect 113824 325042 113876 325048
rect 112536 318776 112588 318782
rect 112536 318718 112588 318724
rect 113272 302388 113324 302394
rect 113272 302330 113324 302336
rect 112536 297016 112588 297022
rect 112536 296958 112588 296964
rect 111812 291949 111918 291977
rect 112548 291963 112576 296958
rect 113180 295588 113232 295594
rect 113180 295530 113232 295536
rect 113192 291963 113220 295530
rect 113284 294794 113312 302330
rect 113836 295594 113864 325042
rect 113928 318170 113956 339390
rect 115124 337482 115152 339487
rect 115216 337958 115244 340054
rect 115400 339946 115428 344986
rect 115308 339918 115428 339946
rect 115204 337952 115256 337958
rect 115204 337894 115256 337900
rect 115216 337754 115244 337894
rect 115204 337748 115256 337754
rect 115204 337690 115256 337696
rect 115112 337476 115164 337482
rect 115112 337418 115164 337424
rect 115308 327146 115336 339918
rect 115388 337748 115440 337754
rect 115388 337690 115440 337696
rect 115296 327140 115348 327146
rect 115296 327082 115348 327088
rect 115400 326602 115428 337690
rect 115388 326596 115440 326602
rect 115388 326538 115440 326544
rect 115296 326528 115348 326534
rect 115296 326470 115348 326476
rect 113916 318164 113968 318170
rect 113916 318106 113968 318112
rect 115204 318096 115256 318102
rect 115204 318038 115256 318044
rect 114652 315988 114704 315994
rect 114652 315930 114704 315936
rect 114664 315382 114692 315930
rect 114652 315376 114704 315382
rect 114652 315318 114704 315324
rect 113824 295588 113876 295594
rect 113824 295530 113876 295536
rect 113284 294766 114324 294794
rect 114190 294672 114246 294681
rect 114190 294607 114246 294616
rect 105004 291910 105466 291938
rect 103150 291887 103206 291896
rect 114204 291870 114232 294607
rect 114296 291977 114324 294766
rect 114664 291977 114692 315318
rect 115216 295526 115244 318038
rect 115308 315382 115336 326470
rect 115296 315376 115348 315382
rect 115296 315318 115348 315324
rect 115584 299674 115612 367639
rect 115952 354006 115980 460838
rect 116044 384713 116072 487766
rect 116136 469198 116164 560322
rect 116584 555484 116636 555490
rect 116584 555426 116636 555432
rect 116400 495508 116452 495514
rect 116400 495450 116452 495456
rect 116412 491298 116440 495450
rect 116400 491292 116452 491298
rect 116400 491234 116452 491240
rect 116124 469192 116176 469198
rect 116124 469134 116176 469140
rect 116596 463690 116624 555426
rect 117332 489870 117360 586638
rect 118792 585200 118844 585206
rect 118792 585142 118844 585148
rect 118700 583840 118752 583846
rect 118700 583782 118752 583788
rect 117412 567860 117464 567866
rect 117412 567802 117464 567808
rect 117424 500342 117452 567802
rect 117964 567316 118016 567322
rect 117964 567258 118016 567264
rect 117412 500336 117464 500342
rect 117412 500278 117464 500284
rect 117502 496088 117558 496097
rect 117502 496023 117558 496032
rect 117320 489864 117372 489870
rect 117320 489806 117372 489812
rect 117412 482996 117464 483002
rect 117412 482938 117464 482944
rect 116860 465724 116912 465730
rect 116860 465666 116912 465672
rect 116872 465050 116900 465666
rect 116860 465044 116912 465050
rect 116860 464986 116912 464992
rect 116584 463684 116636 463690
rect 116584 463626 116636 463632
rect 117228 398268 117280 398274
rect 117228 398210 117280 398216
rect 117240 397594 117268 398210
rect 116584 397588 116636 397594
rect 116584 397530 116636 397536
rect 117228 397588 117280 397594
rect 117228 397530 117280 397536
rect 116124 391332 116176 391338
rect 116124 391274 116176 391280
rect 116030 384704 116086 384713
rect 116030 384639 116086 384648
rect 116030 360632 116086 360641
rect 116030 360567 116086 360576
rect 115940 354000 115992 354006
rect 115938 353968 115940 353977
rect 115992 353968 115994 353977
rect 115938 353903 115994 353912
rect 115768 338026 115796 340068
rect 115756 338020 115808 338026
rect 115756 337962 115808 337968
rect 116044 329254 116072 360567
rect 116136 355745 116164 391274
rect 116596 370025 116624 397530
rect 117424 384985 117452 482938
rect 117516 400926 117544 496023
rect 117686 480856 117742 480865
rect 117686 480791 117742 480800
rect 117596 402348 117648 402354
rect 117596 402290 117648 402296
rect 117504 400920 117556 400926
rect 117504 400862 117556 400868
rect 117504 396908 117556 396914
rect 117504 396850 117556 396856
rect 117410 384976 117466 384985
rect 117410 384911 117466 384920
rect 117320 380316 117372 380322
rect 117320 380258 117372 380264
rect 117332 373425 117360 380258
rect 117318 373416 117374 373425
rect 117318 373351 117374 373360
rect 117332 373318 117360 373351
rect 117320 373312 117372 373318
rect 117320 373254 117372 373260
rect 116582 370016 116638 370025
rect 116582 369951 116638 369960
rect 117410 365256 117466 365265
rect 117410 365191 117466 365200
rect 117424 365022 117452 365191
rect 117412 365016 117464 365022
rect 117412 364958 117464 364964
rect 116122 355736 116178 355745
rect 116122 355671 116178 355680
rect 117516 351665 117544 396850
rect 117608 361865 117636 402290
rect 117700 380186 117728 480791
rect 117976 476134 118004 567258
rect 118712 494766 118740 583782
rect 118804 539170 118832 585142
rect 118792 539164 118844 539170
rect 118792 539106 118844 539112
rect 118792 539028 118844 539034
rect 118792 538970 118844 538976
rect 118700 494760 118752 494766
rect 118700 494702 118752 494708
rect 117964 476128 118016 476134
rect 117964 476070 118016 476076
rect 117976 475998 118004 476070
rect 117964 475992 118016 475998
rect 117964 475934 118016 475940
rect 118804 438870 118832 538970
rect 118896 536722 118924 588542
rect 121644 586764 121696 586770
rect 121644 586706 121696 586712
rect 120172 583908 120224 583914
rect 120172 583850 120224 583856
rect 120080 582548 120132 582554
rect 120080 582490 120132 582496
rect 118976 553512 119028 553518
rect 118976 553454 119028 553460
rect 118884 536716 118936 536722
rect 118884 536658 118936 536664
rect 118896 536178 118924 536658
rect 118884 536172 118936 536178
rect 118884 536114 118936 536120
rect 118884 534744 118936 534750
rect 118884 534686 118936 534692
rect 118792 438864 118844 438870
rect 118792 438806 118844 438812
rect 118896 438802 118924 534686
rect 118988 460902 119016 553454
rect 119068 494896 119120 494902
rect 119068 494838 119120 494844
rect 118976 460896 119028 460902
rect 118976 460838 119028 460844
rect 118884 438796 118936 438802
rect 118884 438738 118936 438744
rect 119080 391241 119108 494838
rect 120092 493950 120120 582490
rect 120184 538966 120212 583850
rect 121460 581052 121512 581058
rect 121460 580994 121512 581000
rect 120264 570036 120316 570042
rect 120264 569978 120316 569984
rect 120172 538960 120224 538966
rect 120172 538902 120224 538908
rect 120172 534812 120224 534818
rect 120172 534754 120224 534760
rect 120080 493944 120132 493950
rect 120080 493886 120132 493892
rect 120092 493270 120120 493886
rect 120080 493264 120132 493270
rect 120080 493206 120132 493212
rect 120080 491292 120132 491298
rect 120080 491234 120132 491240
rect 119344 448656 119396 448662
rect 119344 448598 119396 448604
rect 119066 391232 119122 391241
rect 119066 391167 119122 391176
rect 117964 388204 118016 388210
rect 117964 388146 118016 388152
rect 117976 387938 118004 388146
rect 117964 387932 118016 387938
rect 117964 387874 118016 387880
rect 118700 387184 118752 387190
rect 118700 387126 118752 387132
rect 118712 386510 118740 387126
rect 118700 386504 118752 386510
rect 118700 386446 118752 386452
rect 118514 384976 118570 384985
rect 118514 384911 118570 384920
rect 118528 384334 118556 384911
rect 118516 384328 118568 384334
rect 118054 384296 118110 384305
rect 118516 384270 118568 384276
rect 118054 384231 118110 384240
rect 118068 383722 118096 384231
rect 118056 383716 118108 383722
rect 118056 383658 118108 383664
rect 118146 383616 118202 383625
rect 118146 383551 118202 383560
rect 118160 382294 118188 383551
rect 118148 382288 118200 382294
rect 118148 382230 118200 382236
rect 118606 382256 118662 382265
rect 118606 382191 118608 382200
rect 118660 382191 118662 382200
rect 118608 382162 118660 382168
rect 118606 381576 118662 381585
rect 118606 381511 118608 381520
rect 118660 381511 118662 381520
rect 118608 381482 118660 381488
rect 118606 380896 118662 380905
rect 118606 380831 118662 380840
rect 118620 380390 118648 380831
rect 118608 380384 118660 380390
rect 118608 380326 118660 380332
rect 117688 380180 117740 380186
rect 117688 380122 117740 380128
rect 118332 380180 118384 380186
rect 118332 380122 118384 380128
rect 118344 379545 118372 380122
rect 118330 379536 118386 379545
rect 118330 379471 118386 379480
rect 118606 378856 118662 378865
rect 118606 378791 118662 378800
rect 118620 378758 118648 378791
rect 118608 378752 118660 378758
rect 118608 378694 118660 378700
rect 118056 378276 118108 378282
rect 118056 378218 118108 378224
rect 118068 378185 118096 378218
rect 118054 378176 118110 378185
rect 118054 378111 118110 378120
rect 117870 376816 117926 376825
rect 117870 376751 117872 376760
rect 117924 376751 117926 376760
rect 117872 376722 117924 376728
rect 118608 376712 118660 376718
rect 118608 376654 118660 376660
rect 118514 376136 118570 376145
rect 118514 376071 118570 376080
rect 118528 375426 118556 376071
rect 118620 375465 118648 376654
rect 118606 375456 118662 375465
rect 118516 375420 118568 375426
rect 118606 375391 118662 375400
rect 118516 375362 118568 375368
rect 118608 375352 118660 375358
rect 118608 375294 118660 375300
rect 118620 374105 118648 375294
rect 118606 374096 118662 374105
rect 118606 374031 118662 374040
rect 118054 372736 118110 372745
rect 118054 372671 118110 372680
rect 118068 372638 118096 372671
rect 118056 372632 118108 372638
rect 118056 372574 118108 372580
rect 117870 371376 117926 371385
rect 117870 371311 117926 371320
rect 117884 371278 117912 371311
rect 117872 371272 117924 371278
rect 117872 371214 117924 371220
rect 118606 370696 118662 370705
rect 118606 370631 118662 370640
rect 118620 370598 118648 370631
rect 118608 370592 118660 370598
rect 118608 370534 118660 370540
rect 118238 370016 118294 370025
rect 118238 369951 118240 369960
rect 118292 369951 118294 369960
rect 118240 369922 118292 369928
rect 118608 369844 118660 369850
rect 118608 369786 118660 369792
rect 118620 368665 118648 369786
rect 118606 368656 118662 368665
rect 118606 368591 118662 368600
rect 118606 367976 118662 367985
rect 118606 367911 118608 367920
rect 118660 367911 118662 367920
rect 118608 367882 118660 367888
rect 118608 367056 118660 367062
rect 118608 366998 118660 367004
rect 118620 365945 118648 366998
rect 118606 365936 118662 365945
rect 118606 365871 118662 365880
rect 117872 365696 117924 365702
rect 117872 365638 117924 365644
rect 117884 364585 117912 365638
rect 117870 364576 117926 364585
rect 117870 364511 117926 364520
rect 118148 364336 118200 364342
rect 118148 364278 118200 364284
rect 118160 363225 118188 364278
rect 118146 363216 118202 363225
rect 118146 363151 118202 363160
rect 118608 362908 118660 362914
rect 118608 362850 118660 362856
rect 118620 362545 118648 362850
rect 118606 362536 118662 362545
rect 118606 362471 118662 362480
rect 117594 361856 117650 361865
rect 117594 361791 117650 361800
rect 118606 361856 118662 361865
rect 118606 361791 118608 361800
rect 118660 361791 118662 361800
rect 118608 361762 118660 361768
rect 118056 361480 118108 361486
rect 118056 361422 118108 361428
rect 118068 361185 118096 361422
rect 118054 361176 118110 361185
rect 118054 361111 118110 361120
rect 118516 360188 118568 360194
rect 118516 360130 118568 360136
rect 118528 359145 118556 360130
rect 118608 360120 118660 360126
rect 118608 360062 118660 360068
rect 118620 359825 118648 360062
rect 118606 359816 118662 359825
rect 118606 359751 118662 359760
rect 118514 359136 118570 359145
rect 118514 359071 118570 359080
rect 118606 358456 118662 358465
rect 118606 358391 118662 358400
rect 118620 358086 118648 358391
rect 118608 358080 118660 358086
rect 118608 358022 118660 358028
rect 118608 357400 118660 357406
rect 118608 357342 118660 357348
rect 118620 357105 118648 357342
rect 118606 357096 118662 357105
rect 118606 357031 118662 357040
rect 118608 356720 118660 356726
rect 118608 356662 118660 356668
rect 118620 356425 118648 356662
rect 118606 356416 118662 356425
rect 118606 356351 118662 356360
rect 118146 355736 118202 355745
rect 118146 355671 118202 355680
rect 118160 354754 118188 355671
rect 118148 354748 118200 354754
rect 118148 354690 118200 354696
rect 117780 354680 117832 354686
rect 117780 354622 117832 354628
rect 117792 354385 117820 354622
rect 117778 354376 117834 354385
rect 117778 354311 117834 354320
rect 118606 353016 118662 353025
rect 118606 352951 118662 352960
rect 118620 352578 118648 352951
rect 118608 352572 118660 352578
rect 118608 352514 118660 352520
rect 118056 351892 118108 351898
rect 118056 351834 118108 351840
rect 117502 351656 117558 351665
rect 117502 351591 117558 351600
rect 118068 350985 118096 351834
rect 118606 351656 118662 351665
rect 118606 351591 118662 351600
rect 118620 351218 118648 351591
rect 118608 351212 118660 351218
rect 118608 351154 118660 351160
rect 118054 350976 118110 350985
rect 118054 350911 118110 350920
rect 118608 350328 118660 350334
rect 118606 350296 118608 350305
rect 118660 350296 118662 350305
rect 118606 350231 118662 350240
rect 118712 349858 118740 386446
rect 119356 368626 119384 448598
rect 119436 421592 119488 421598
rect 119436 421534 119488 421540
rect 119448 389842 119476 421534
rect 119436 389836 119488 389842
rect 119436 389778 119488 389784
rect 119448 389502 119476 389778
rect 119436 389496 119488 389502
rect 119436 389438 119488 389444
rect 119436 388068 119488 388074
rect 119436 388010 119488 388016
rect 119448 376106 119476 388010
rect 119528 388000 119580 388006
rect 119528 387942 119580 387948
rect 119540 382974 119568 387942
rect 120092 387705 120120 491234
rect 120184 437374 120212 534754
rect 120276 476066 120304 569978
rect 121472 494018 121500 580994
rect 121552 537600 121604 537606
rect 121552 537542 121604 537548
rect 121460 494012 121512 494018
rect 121460 493954 121512 493960
rect 121472 493406 121500 493954
rect 121460 493400 121512 493406
rect 121460 493342 121512 493348
rect 120356 491224 120408 491230
rect 120356 491166 120408 491172
rect 120264 476060 120316 476066
rect 120264 476002 120316 476008
rect 120172 437368 120224 437374
rect 120172 437310 120224 437316
rect 120368 421598 120396 491166
rect 121564 438938 121592 537542
rect 121656 532030 121684 586706
rect 123116 586628 123168 586634
rect 123116 586570 123168 586576
rect 123024 586560 123076 586566
rect 123024 586502 123076 586508
rect 122748 575544 122800 575550
rect 122748 575486 122800 575492
rect 121736 532160 121788 532166
rect 121736 532102 121788 532108
rect 121644 532024 121696 532030
rect 121644 531966 121696 531972
rect 121644 465044 121696 465050
rect 121644 464986 121696 464992
rect 121552 438932 121604 438938
rect 121552 438874 121604 438880
rect 120356 421592 120408 421598
rect 120356 421534 120408 421540
rect 120264 402280 120316 402286
rect 120264 402222 120316 402228
rect 120078 387696 120134 387705
rect 120078 387631 120134 387640
rect 119528 382968 119580 382974
rect 119528 382910 119580 382916
rect 119436 376100 119488 376106
rect 119436 376042 119488 376048
rect 120172 376032 120224 376038
rect 120172 375974 120224 375980
rect 120184 375426 120212 375974
rect 120172 375420 120224 375426
rect 120172 375362 120224 375368
rect 119436 368824 119488 368830
rect 119436 368766 119488 368772
rect 119344 368620 119396 368626
rect 119344 368562 119396 368568
rect 117964 349852 118016 349858
rect 117964 349794 118016 349800
rect 118700 349852 118752 349858
rect 118700 349794 118752 349800
rect 117688 349036 117740 349042
rect 117688 348978 117740 348984
rect 117700 348265 117728 348978
rect 117686 348256 117742 348265
rect 117686 348191 117742 348200
rect 117412 347744 117464 347750
rect 117412 347686 117464 347692
rect 117424 347585 117452 347686
rect 117410 347576 117466 347585
rect 117410 347511 117466 347520
rect 117872 343596 117924 343602
rect 117872 343538 117924 343544
rect 117502 343496 117558 343505
rect 117502 343431 117558 343440
rect 117516 342990 117544 343431
rect 117504 342984 117556 342990
rect 117504 342926 117556 342932
rect 117688 342916 117740 342922
rect 117688 342858 117740 342864
rect 117412 340876 117464 340882
rect 117412 340818 117464 340824
rect 117320 340808 117372 340814
rect 117318 340776 117320 340785
rect 117372 340776 117374 340785
rect 117318 340711 117374 340720
rect 117332 339522 117360 340711
rect 117424 340105 117452 340818
rect 117410 340096 117466 340105
rect 117410 340031 117466 340040
rect 117320 339516 117372 339522
rect 117320 339458 117372 339464
rect 117700 339182 117728 342858
rect 117884 342825 117912 343538
rect 117870 342816 117926 342825
rect 117870 342751 117926 342760
rect 117688 339176 117740 339182
rect 117688 339118 117740 339124
rect 117976 336122 118004 349794
rect 118608 349104 118660 349110
rect 118608 349046 118660 349052
rect 118620 348945 118648 349046
rect 118606 348936 118662 348945
rect 118606 348871 118662 348880
rect 118608 346384 118660 346390
rect 118608 346326 118660 346332
rect 118514 346216 118570 346225
rect 118514 346151 118570 346160
rect 118528 345642 118556 346151
rect 118516 345636 118568 345642
rect 118516 345578 118568 345584
rect 118620 345545 118648 346326
rect 118606 345536 118662 345545
rect 118606 345471 118662 345480
rect 118608 345024 118660 345030
rect 118608 344966 118660 344972
rect 118620 344865 118648 344966
rect 118606 344856 118662 344865
rect 118606 344791 118662 344800
rect 118608 342236 118660 342242
rect 118608 342178 118660 342184
rect 118620 342145 118648 342178
rect 118606 342136 118662 342145
rect 118606 342071 118662 342080
rect 119356 339454 119384 368562
rect 119344 339448 119396 339454
rect 119344 339390 119396 339396
rect 117964 336116 118016 336122
rect 117964 336058 118016 336064
rect 116032 329248 116084 329254
rect 116032 329190 116084 329196
rect 117964 323740 118016 323746
rect 117964 323682 118016 323688
rect 117320 319592 117372 319598
rect 117320 319534 117372 319540
rect 115848 317552 115900 317558
rect 115848 317494 115900 317500
rect 115860 316878 115888 317494
rect 116676 317484 116728 317490
rect 116676 317426 116728 317432
rect 115848 316872 115900 316878
rect 115848 316814 115900 316820
rect 116584 313948 116636 313954
rect 116584 313890 116636 313896
rect 115572 299668 115624 299674
rect 115572 299610 115624 299616
rect 116596 296954 116624 313890
rect 116688 302394 116716 317426
rect 116676 302388 116728 302394
rect 116676 302330 116728 302336
rect 116584 296948 116636 296954
rect 116584 296890 116636 296896
rect 115204 295520 115256 295526
rect 115204 295462 115256 295468
rect 115756 295520 115808 295526
rect 115756 295462 115808 295468
rect 114296 291949 114494 291977
rect 114664 291949 115138 291977
rect 115768 291963 115796 295462
rect 116596 291977 116624 296890
rect 117044 295316 117096 295322
rect 117044 295258 117096 295264
rect 116426 291949 116624 291977
rect 117056 291963 117084 295258
rect 117228 294092 117280 294098
rect 117228 294034 117280 294040
rect 117240 291922 117268 294034
rect 117332 291977 117360 319534
rect 117976 306374 118004 323682
rect 117976 306346 118096 306374
rect 117872 300280 117924 300286
rect 117872 300222 117924 300228
rect 117884 299538 117912 300222
rect 117872 299532 117924 299538
rect 117872 299474 117924 299480
rect 117332 291949 117714 291977
rect 117884 291938 117912 299474
rect 118068 292466 118096 306346
rect 118974 295216 119030 295225
rect 118974 295151 119030 295160
rect 118056 292460 118108 292466
rect 118056 292402 118108 292408
rect 118988 291963 119016 295151
rect 119448 294778 119476 368766
rect 120080 361820 120132 361826
rect 120080 361762 120132 361768
rect 119528 361004 119580 361010
rect 119528 360946 119580 360952
rect 119540 337890 119568 360946
rect 119712 345636 119764 345642
rect 119712 345578 119764 345584
rect 119528 337884 119580 337890
rect 119528 337826 119580 337832
rect 119436 294772 119488 294778
rect 119436 294714 119488 294720
rect 119620 294704 119672 294710
rect 119620 294646 119672 294652
rect 91954 291858 92348 291864
rect 91954 291842 92336 291858
rect 113850 291842 114232 291870
rect 117228 291916 117280 291922
rect 117884 291910 118346 291938
rect 119632 291924 119660 294646
rect 117228 291858 117280 291864
rect 69768 291230 70058 291258
rect 69768 289202 69796 291230
rect 69756 289196 69808 289202
rect 69756 289138 69808 289144
rect 119724 267734 119752 345578
rect 119896 308508 119948 308514
rect 119896 308450 119948 308456
rect 119908 304026 119936 308450
rect 119896 304020 119948 304026
rect 119896 303962 119948 303968
rect 119724 267706 119844 267734
rect 69202 260264 69258 260273
rect 69202 260199 69258 260208
rect 69202 251832 69258 251841
rect 69202 251767 69258 251776
rect 69216 222154 69244 251767
rect 119816 251161 119844 267706
rect 119802 251152 119858 251161
rect 119802 251087 119858 251096
rect 69846 247072 69902 247081
rect 69846 247007 69902 247016
rect 69860 239426 69888 247007
rect 120092 241505 120120 361762
rect 120184 326466 120212 375362
rect 120276 361010 120304 402222
rect 121460 389972 121512 389978
rect 121460 389914 121512 389920
rect 120724 389428 120776 389434
rect 120724 389370 120776 389376
rect 120736 389298 120764 389370
rect 121472 389298 121500 389914
rect 121656 389434 121684 464986
rect 121748 462913 121776 532102
rect 121828 493944 121880 493950
rect 121828 493886 121880 493892
rect 121734 462904 121790 462913
rect 121734 462839 121790 462848
rect 121840 402974 121868 493886
rect 122760 484378 122788 575486
rect 122932 537668 122984 537674
rect 122932 537610 122984 537616
rect 122760 484350 122880 484378
rect 122852 483682 122880 484350
rect 122840 483676 122892 483682
rect 122840 483618 122892 483624
rect 122840 475380 122892 475386
rect 122840 475322 122892 475328
rect 121840 402946 122328 402974
rect 121644 389428 121696 389434
rect 121644 389370 121696 389376
rect 120724 389292 120776 389298
rect 120724 389234 120776 389240
rect 121460 389292 121512 389298
rect 121460 389234 121512 389240
rect 122104 389292 122156 389298
rect 122104 389234 122156 389240
rect 120264 361004 120316 361010
rect 120264 360946 120316 360952
rect 120262 358728 120318 358737
rect 120262 358663 120318 358672
rect 120276 335102 120304 358663
rect 120736 358086 120764 389234
rect 121460 376780 121512 376786
rect 121460 376722 121512 376728
rect 121472 374678 121500 376722
rect 121460 374672 121512 374678
rect 121460 374614 121512 374620
rect 121460 372632 121512 372638
rect 121460 372574 121512 372580
rect 121472 370530 121500 372574
rect 121460 370524 121512 370530
rect 121460 370466 121512 370472
rect 121460 369980 121512 369986
rect 121460 369922 121512 369928
rect 121472 369170 121500 369922
rect 121460 369164 121512 369170
rect 121460 369106 121512 369112
rect 120724 358080 120776 358086
rect 120724 358022 120776 358028
rect 121460 336048 121512 336054
rect 121460 335990 121512 335996
rect 120264 335096 120316 335102
rect 120264 335038 120316 335044
rect 121472 334626 121500 335990
rect 121460 334620 121512 334626
rect 121460 334562 121512 334568
rect 122116 331226 122144 389234
rect 122300 387977 122328 402946
rect 122286 387968 122342 387977
rect 122286 387903 122342 387912
rect 122194 386608 122250 386617
rect 122194 386543 122250 386552
rect 122208 376825 122236 386543
rect 122300 385150 122328 387903
rect 122288 385144 122340 385150
rect 122288 385086 122340 385092
rect 122472 380384 122524 380390
rect 122472 380326 122524 380332
rect 122484 380225 122512 380326
rect 122470 380216 122526 380225
rect 122470 380151 122526 380160
rect 122194 376816 122250 376825
rect 122194 376751 122250 376760
rect 122656 369844 122708 369850
rect 122656 369786 122708 369792
rect 122194 359272 122250 359281
rect 122194 359207 122250 359216
rect 122208 337346 122236 359207
rect 122668 358154 122696 369786
rect 122852 367946 122880 475322
rect 122944 438734 122972 537610
rect 123036 494834 123064 586502
rect 123128 496330 123156 586570
rect 125690 583808 125746 583817
rect 125690 583743 125746 583752
rect 124220 574116 124272 574122
rect 124220 574058 124272 574064
rect 123208 564528 123260 564534
rect 123208 564470 123260 564476
rect 123116 496324 123168 496330
rect 123116 496266 123168 496272
rect 123024 494828 123076 494834
rect 123024 494770 123076 494776
rect 123220 472666 123248 564470
rect 123300 496188 123352 496194
rect 123300 496130 123352 496136
rect 123208 472660 123260 472666
rect 123208 472602 123260 472608
rect 122932 438728 122984 438734
rect 122932 438670 122984 438676
rect 123312 398138 123340 496130
rect 123392 483676 123444 483682
rect 123392 483618 123444 483624
rect 123404 483177 123432 483618
rect 123390 483168 123446 483177
rect 123390 483103 123446 483112
rect 124232 481574 124260 574058
rect 124588 552084 124640 552090
rect 124588 552026 124640 552032
rect 124496 538892 124548 538898
rect 124496 538834 124548 538840
rect 124404 493604 124456 493610
rect 124404 493546 124456 493552
rect 124220 481568 124272 481574
rect 124220 481510 124272 481516
rect 124312 476128 124364 476134
rect 124312 476070 124364 476076
rect 124128 472660 124180 472666
rect 124128 472602 124180 472608
rect 124140 471306 124168 472602
rect 124128 471300 124180 471306
rect 124128 471242 124180 471248
rect 124220 458924 124272 458930
rect 124220 458866 124272 458872
rect 123300 398132 123352 398138
rect 123300 398074 123352 398080
rect 123760 385144 123812 385150
rect 123760 385086 123812 385092
rect 123484 372700 123536 372706
rect 123484 372642 123536 372648
rect 122840 367940 122892 367946
rect 122840 367882 122892 367888
rect 122852 367094 122880 367882
rect 122760 367066 122880 367094
rect 122656 358148 122708 358154
rect 122656 358090 122708 358096
rect 122760 340270 122788 367066
rect 122748 340264 122800 340270
rect 122748 340206 122800 340212
rect 122196 337340 122248 337346
rect 122196 337282 122248 337288
rect 122196 331900 122248 331906
rect 122196 331842 122248 331848
rect 122104 331220 122156 331226
rect 122104 331162 122156 331168
rect 120172 326460 120224 326466
rect 120172 326402 120224 326408
rect 122104 319660 122156 319666
rect 122104 319602 122156 319608
rect 120170 296032 120226 296041
rect 120170 295967 120226 295976
rect 120184 275505 120212 295967
rect 121460 292528 121512 292534
rect 121460 292470 121512 292476
rect 121472 291825 121500 292470
rect 121458 291816 121514 291825
rect 121458 291751 121514 291760
rect 121550 291136 121606 291145
rect 121550 291071 121606 291080
rect 121458 290456 121514 290465
rect 121458 290391 121514 290400
rect 121472 289950 121500 290391
rect 121564 290018 121592 291071
rect 121552 290012 121604 290018
rect 121552 289954 121604 289960
rect 121460 289944 121512 289950
rect 121460 289886 121512 289892
rect 121552 289808 121604 289814
rect 121458 289776 121514 289785
rect 121552 289750 121604 289756
rect 121458 289711 121460 289720
rect 121512 289711 121514 289720
rect 121460 289682 121512 289688
rect 121564 289105 121592 289750
rect 121550 289096 121606 289105
rect 121550 289031 121606 289040
rect 121458 288416 121514 288425
rect 121458 288351 121460 288360
rect 121512 288351 121514 288360
rect 121460 288322 121512 288328
rect 121552 288312 121604 288318
rect 121552 288254 121604 288260
rect 121564 287745 121592 288254
rect 121550 287736 121606 287745
rect 121550 287671 121606 287680
rect 121458 287056 121514 287065
rect 121458 286991 121514 287000
rect 121552 287020 121604 287026
rect 121472 286890 121500 286991
rect 121552 286962 121604 286968
rect 121460 286884 121512 286890
rect 121460 286826 121512 286832
rect 121564 286385 121592 286962
rect 121644 286952 121696 286958
rect 121644 286894 121696 286900
rect 121550 286376 121606 286385
rect 121550 286311 121606 286320
rect 121656 285705 121684 286894
rect 121642 285696 121698 285705
rect 121460 285660 121512 285666
rect 121642 285631 121698 285640
rect 121460 285602 121512 285608
rect 121472 285025 121500 285602
rect 121552 285592 121604 285598
rect 121552 285534 121604 285540
rect 121458 285016 121514 285025
rect 121458 284951 121514 284960
rect 121564 284345 121592 285534
rect 121644 285048 121696 285054
rect 121644 284990 121696 284996
rect 121550 284336 121606 284345
rect 121460 284300 121512 284306
rect 121550 284271 121606 284280
rect 121460 284242 121512 284248
rect 121472 283665 121500 284242
rect 121458 283656 121514 283665
rect 121458 283591 121514 283600
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121458 281616 121514 281625
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121552 281512 121604 281518
rect 121552 281454 121604 281460
rect 121564 280945 121592 281454
rect 121550 280936 121606 280945
rect 121550 280871 121606 280880
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121656 279585 121684 284990
rect 121642 279576 121698 279585
rect 121642 279511 121698 279520
rect 121458 278896 121514 278905
rect 121458 278831 121514 278840
rect 121472 278798 121500 278831
rect 121460 278792 121512 278798
rect 121460 278734 121512 278740
rect 121458 277536 121514 277545
rect 121458 277471 121514 277480
rect 121472 277438 121500 277471
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 121460 277296 121512 277302
rect 121460 277238 121512 277244
rect 121472 276865 121500 277238
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121458 276176 121514 276185
rect 121458 276111 121514 276120
rect 121472 276078 121500 276111
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 120170 275496 120226 275505
rect 120170 275431 120226 275440
rect 120722 275496 120778 275505
rect 120722 275431 120778 275440
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120078 241496 120134 241505
rect 120078 241431 120134 241440
rect 119988 240168 120040 240174
rect 69952 240094 70058 240122
rect 119646 240094 119752 240122
rect 119988 240110 120040 240116
rect 69848 239420 69900 239426
rect 69848 239362 69900 239368
rect 69952 238338 69980 240094
rect 70400 239828 70452 239834
rect 70400 239770 70452 239776
rect 69940 238332 69992 238338
rect 69940 238274 69992 238280
rect 69204 222148 69256 222154
rect 69204 222090 69256 222096
rect 70412 192574 70440 239770
rect 70688 238754 70716 240037
rect 71320 239834 71348 240037
rect 71308 239828 71360 239834
rect 71308 239770 71360 239776
rect 70504 238726 70716 238754
rect 70504 226098 70532 238726
rect 71976 238202 72004 240037
rect 72422 239864 72478 239873
rect 72422 239799 72478 239808
rect 71964 238196 72016 238202
rect 71964 238138 72016 238144
rect 70492 226092 70544 226098
rect 70492 226034 70544 226040
rect 72436 213926 72464 239799
rect 72620 238678 72648 240037
rect 72608 238672 72660 238678
rect 72608 238614 72660 238620
rect 73264 238134 73292 240037
rect 73804 239624 73856 239630
rect 73804 239566 73856 239572
rect 73252 238128 73304 238134
rect 73252 238070 73304 238076
rect 73816 230314 73844 239566
rect 73908 235822 73936 240037
rect 74552 238754 74580 240037
rect 74552 238726 74672 238754
rect 73896 235816 73948 235822
rect 73896 235758 73948 235764
rect 74540 233912 74592 233918
rect 74540 233854 74592 233860
rect 73804 230308 73856 230314
rect 73804 230250 73856 230256
rect 72424 213920 72476 213926
rect 72424 213862 72476 213868
rect 74552 206378 74580 233854
rect 74644 222018 74672 238726
rect 75196 233918 75224 240037
rect 75184 233912 75236 233918
rect 75184 233854 75236 233860
rect 75840 233073 75868 240037
rect 76012 239828 76064 239834
rect 76012 239770 76064 239776
rect 75826 233064 75882 233073
rect 75826 232999 75882 233008
rect 76024 224874 76052 239770
rect 76380 239556 76432 239562
rect 76380 239498 76432 239504
rect 76392 238754 76420 239498
rect 76484 239442 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 76484 239414 76696 239442
rect 76392 238726 76604 238754
rect 76012 224868 76064 224874
rect 76012 224810 76064 224816
rect 74632 222012 74684 222018
rect 74632 221954 74684 221960
rect 74540 206372 74592 206378
rect 74540 206314 74592 206320
rect 76576 205018 76604 238726
rect 76668 237250 76696 239414
rect 77772 239086 77800 240037
rect 78404 239816 78432 240037
rect 78324 239788 78432 239816
rect 77760 239080 77812 239086
rect 77760 239022 77812 239028
rect 76656 237244 76708 237250
rect 76656 237186 76708 237192
rect 76668 230382 76696 237186
rect 76656 230376 76708 230382
rect 76656 230318 76708 230324
rect 78324 219434 78352 239788
rect 79060 238754 79088 240037
rect 79692 239816 79720 240037
rect 77312 219406 78352 219434
rect 78692 238726 79088 238754
rect 79612 239788 79720 239816
rect 77312 207806 77340 219406
rect 77300 207800 77352 207806
rect 77300 207742 77352 207748
rect 76564 205012 76616 205018
rect 76564 204954 76616 204960
rect 78692 200705 78720 238726
rect 79232 238196 79284 238202
rect 79232 238138 79284 238144
rect 79244 233918 79272 238138
rect 79232 233912 79284 233918
rect 79232 233854 79284 233860
rect 79612 219434 79640 239788
rect 80348 238754 80376 240037
rect 78784 219406 79640 219434
rect 80072 238726 80376 238754
rect 78784 217938 78812 219406
rect 78772 217932 78824 217938
rect 78772 217874 78824 217880
rect 80072 213790 80100 238726
rect 80992 238202 81020 240037
rect 80980 238196 81032 238202
rect 80980 238138 81032 238144
rect 81636 233102 81664 240037
rect 82280 238746 82308 240037
rect 82912 239816 82940 240037
rect 82832 239788 82940 239816
rect 82268 238740 82320 238746
rect 82268 238682 82320 238688
rect 81624 233096 81676 233102
rect 81624 233038 81676 233044
rect 82832 231742 82860 239788
rect 83464 239420 83516 239426
rect 83464 239362 83516 239368
rect 82820 231736 82872 231742
rect 82820 231678 82872 231684
rect 80060 213784 80112 213790
rect 80060 213726 80112 213732
rect 78678 200696 78734 200705
rect 78678 200631 78734 200640
rect 83476 198082 83504 239362
rect 83568 238678 83596 240037
rect 83556 238672 83608 238678
rect 83556 238614 83608 238620
rect 83568 229770 83596 238614
rect 84212 233866 84240 240037
rect 84292 239828 84344 239834
rect 84292 239770 84344 239776
rect 84304 233986 84332 239770
rect 84856 238754 84884 240037
rect 85488 239834 85516 240037
rect 85476 239828 85528 239834
rect 85476 239770 85528 239776
rect 85580 238944 85632 238950
rect 85580 238886 85632 238892
rect 84396 238726 84884 238754
rect 84292 233980 84344 233986
rect 84292 233922 84344 233928
rect 84212 233838 84332 233866
rect 84200 233776 84252 233782
rect 84200 233718 84252 233724
rect 83556 229764 83608 229770
rect 83556 229706 83608 229712
rect 83464 198076 83516 198082
rect 83464 198018 83516 198024
rect 70400 192568 70452 192574
rect 70400 192510 70452 192516
rect 69112 191208 69164 191214
rect 69112 191150 69164 191156
rect 84212 188494 84240 233718
rect 84304 219366 84332 233838
rect 84396 227594 84424 238726
rect 85592 234462 85620 238886
rect 86144 237318 86172 240037
rect 86788 238950 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86776 238944 86828 238950
rect 86776 238886 86828 238892
rect 86224 238128 86276 238134
rect 86224 238070 86276 238076
rect 86132 237312 86184 237318
rect 86132 237254 86184 237260
rect 86144 234569 86172 237254
rect 86130 234560 86186 234569
rect 86130 234495 86186 234504
rect 85580 234456 85632 234462
rect 85580 234398 85632 234404
rect 84384 227588 84436 227594
rect 84384 227530 84436 227536
rect 84292 219360 84344 219366
rect 84292 219302 84344 219308
rect 86236 219298 86264 238070
rect 86224 219292 86276 219298
rect 86224 219234 86276 219240
rect 86972 199442 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 87064 238726 87460 238754
rect 87064 231674 87092 238726
rect 88720 238610 88748 240037
rect 88708 238604 88760 238610
rect 88708 238546 88760 238552
rect 88984 238196 89036 238202
rect 88984 238138 89036 238144
rect 87052 231668 87104 231674
rect 87052 231610 87104 231616
rect 88996 212430 89024 238138
rect 89364 235958 89392 240037
rect 89720 239828 89772 239834
rect 89720 239770 89772 239776
rect 89352 235952 89404 235958
rect 89352 235894 89404 235900
rect 88984 212424 89036 212430
rect 88984 212366 89036 212372
rect 86960 199436 87012 199442
rect 86960 199378 87012 199384
rect 89732 195362 89760 239770
rect 90008 238754 90036 240037
rect 90640 239834 90668 240037
rect 90628 239828 90680 239834
rect 90628 239770 90680 239776
rect 89824 238726 90036 238754
rect 89824 205086 89852 238726
rect 91296 235890 91324 240037
rect 91940 238754 91968 240037
rect 92572 239850 92600 240037
rect 93216 239850 93244 240037
rect 91756 238726 91968 238754
rect 92492 239822 92600 239850
rect 93136 239822 93244 239850
rect 91284 235884 91336 235890
rect 91284 235826 91336 235832
rect 91756 235754 91784 238726
rect 91744 235748 91796 235754
rect 91744 235690 91796 235696
rect 91756 227730 91784 235690
rect 91744 227724 91796 227730
rect 91744 227666 91796 227672
rect 89812 205080 89864 205086
rect 89812 205022 89864 205028
rect 89720 195356 89772 195362
rect 89720 195298 89772 195304
rect 92492 192710 92520 239822
rect 93136 219434 93164 239822
rect 92584 219406 93164 219434
rect 92584 216578 92612 219406
rect 92572 216572 92624 216578
rect 92572 216514 92624 216520
rect 93872 214810 93900 240037
rect 94516 238754 94544 240037
rect 95148 239850 95176 240037
rect 93964 238726 94544 238754
rect 95068 239822 95176 239850
rect 95240 239828 95292 239834
rect 93964 223514 93992 238726
rect 95068 227526 95096 239822
rect 95240 239770 95292 239776
rect 95056 227520 95108 227526
rect 95056 227462 95108 227468
rect 95252 224942 95280 239770
rect 95804 237318 95832 240037
rect 96436 239834 96464 240037
rect 96424 239828 96476 239834
rect 96424 239770 96476 239776
rect 97092 238754 97120 240037
rect 97724 239850 97752 240037
rect 96632 238726 97120 238754
rect 97644 239822 97752 239850
rect 95792 237312 95844 237318
rect 95792 237254 95844 237260
rect 95240 224936 95292 224942
rect 95240 224878 95292 224884
rect 93952 223508 94004 223514
rect 93952 223450 94004 223456
rect 93860 214804 93912 214810
rect 93860 214746 93912 214752
rect 96632 203726 96660 238726
rect 97644 228954 97672 239822
rect 98380 235929 98408 240037
rect 99012 239850 99040 240037
rect 98932 239822 99040 239850
rect 98366 235920 98422 235929
rect 98366 235855 98422 235864
rect 97632 228948 97684 228954
rect 97632 228890 97684 228896
rect 98932 219434 98960 239822
rect 99668 238754 99696 240037
rect 100300 239850 100328 240037
rect 98012 219406 98960 219434
rect 99392 238726 99696 238754
rect 100220 239822 100328 239850
rect 98012 204270 98040 219406
rect 99392 208350 99420 238726
rect 100220 229906 100248 239822
rect 100956 238754 100984 240037
rect 101588 239850 101616 240037
rect 100772 238726 100984 238754
rect 101508 239822 101616 239850
rect 102140 239828 102192 239834
rect 100208 229900 100260 229906
rect 100208 229842 100260 229848
rect 99380 208344 99432 208350
rect 99380 208286 99432 208292
rect 98000 204264 98052 204270
rect 98000 204206 98052 204212
rect 96620 203720 96672 203726
rect 96620 203662 96672 203668
rect 100772 194002 100800 238726
rect 101508 220250 101536 239822
rect 102140 239770 102192 239776
rect 101496 220244 101548 220250
rect 101496 220186 101548 220192
rect 102152 211954 102180 239770
rect 102244 223582 102272 240037
rect 102876 239834 102904 240037
rect 102864 239828 102916 239834
rect 102864 239770 102916 239776
rect 103532 237386 103560 240037
rect 104176 239018 104204 240037
rect 104808 239850 104836 240037
rect 104728 239822 104836 239850
rect 104164 239012 104216 239018
rect 104164 238954 104216 238960
rect 103520 237380 103572 237386
rect 103520 237322 103572 237328
rect 102232 223576 102284 223582
rect 102232 223518 102284 223524
rect 104728 219434 104756 239822
rect 105464 238406 105492 240037
rect 105452 238400 105504 238406
rect 105452 238342 105504 238348
rect 105544 238060 105596 238066
rect 105544 238002 105596 238008
rect 103716 219406 104756 219434
rect 103716 213858 103744 219406
rect 103704 213852 103756 213858
rect 103704 213794 103756 213800
rect 102140 211948 102192 211954
rect 102140 211890 102192 211896
rect 105556 209778 105584 238002
rect 106108 235346 106136 240037
rect 106752 235929 106780 240037
rect 107396 237153 107424 240037
rect 107660 239828 107712 239834
rect 107660 239770 107712 239776
rect 107382 237144 107438 237153
rect 107382 237079 107438 237088
rect 106738 235920 106794 235929
rect 106738 235855 106794 235864
rect 106096 235340 106148 235346
rect 106096 235282 106148 235288
rect 105544 209772 105596 209778
rect 105544 209714 105596 209720
rect 107672 205630 107700 239770
rect 108040 238754 108068 240037
rect 108672 239834 108700 240037
rect 108660 239828 108712 239834
rect 108660 239770 108712 239776
rect 107764 238726 108068 238754
rect 107764 211138 107792 238726
rect 109040 234592 109092 234598
rect 109040 234534 109092 234540
rect 109052 234190 109080 234534
rect 109972 234190 110000 240037
rect 110604 239850 110632 240037
rect 110420 239828 110472 239834
rect 110420 239770 110472 239776
rect 110524 239822 110632 239850
rect 111248 239834 111276 240037
rect 111892 239850 111920 240037
rect 111236 239828 111288 239834
rect 109040 234184 109092 234190
rect 109040 234126 109092 234132
rect 109960 234184 110012 234190
rect 109960 234126 110012 234132
rect 107752 211132 107804 211138
rect 107752 211074 107804 211080
rect 107660 205624 107712 205630
rect 107660 205566 107712 205572
rect 100760 193996 100812 194002
rect 100760 193938 100812 193944
rect 92480 192704 92532 192710
rect 92480 192646 92532 192652
rect 84200 188488 84252 188494
rect 84200 188430 84252 188436
rect 69018 186960 69074 186969
rect 69018 186895 69074 186904
rect 102048 184952 102100 184958
rect 102048 184894 102100 184900
rect 100666 183696 100722 183705
rect 100666 183631 100722 183640
rect 97816 179444 97868 179450
rect 97816 179386 97868 179392
rect 97828 177041 97856 179386
rect 98736 178424 98788 178430
rect 98736 178366 98788 178372
rect 97814 177032 97870 177041
rect 97814 176967 97870 176976
rect 98748 176769 98776 178366
rect 100680 176769 100708 183631
rect 102060 177721 102088 184894
rect 107568 183660 107620 183666
rect 107568 183602 107620 183608
rect 105726 180840 105782 180849
rect 105726 180775 105782 180784
rect 105740 177721 105768 180775
rect 107580 177721 107608 183602
rect 109052 182850 109080 234126
rect 110432 187134 110460 239770
rect 110524 218006 110552 239822
rect 111236 239770 111288 239776
rect 111812 239822 111920 239850
rect 110512 218000 110564 218006
rect 110512 217942 110564 217948
rect 110524 210458 110552 217942
rect 110512 210452 110564 210458
rect 110512 210394 110564 210400
rect 111812 203658 111840 239822
rect 112548 238882 112576 240037
rect 111892 238876 111944 238882
rect 111892 238818 111944 238824
rect 112536 238876 112588 238882
rect 112536 238818 112588 238824
rect 111904 229838 111932 238818
rect 113192 237386 113220 240037
rect 113180 237380 113232 237386
rect 113180 237322 113232 237328
rect 113836 237250 113864 240037
rect 114480 238882 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 238876 114520 238882
rect 114468 238818 114520 238824
rect 114468 237380 114520 237386
rect 114468 237322 114520 237328
rect 113824 237244 113876 237250
rect 113824 237186 113876 237192
rect 111892 229832 111944 229838
rect 111892 229774 111944 229780
rect 111800 203652 111852 203658
rect 111800 203594 111852 203600
rect 114480 188426 114508 237322
rect 114572 212498 114600 239770
rect 115124 238474 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 116412 238754 116440 240037
rect 117056 239737 117084 240037
rect 117042 239728 117098 239737
rect 117042 239663 117098 239672
rect 115952 238726 116440 238754
rect 115112 238468 115164 238474
rect 115112 238410 115164 238416
rect 114560 212492 114612 212498
rect 114560 212434 114612 212440
rect 115952 202366 115980 238726
rect 117700 235006 117728 240037
rect 118344 238542 118372 240037
rect 118988 238746 119016 240037
rect 118976 238740 119028 238746
rect 118976 238682 119028 238688
rect 118332 238536 118384 238542
rect 118332 238478 118384 238484
rect 118608 235748 118660 235754
rect 118608 235690 118660 235696
rect 118620 235006 118648 235690
rect 117688 235000 117740 235006
rect 117688 234942 117740 234948
rect 118608 235000 118660 235006
rect 118608 234942 118660 234948
rect 115940 202360 115992 202366
rect 115940 202302 115992 202308
rect 118620 191146 118648 234942
rect 119724 219434 119752 240094
rect 120000 238338 120028 240110
rect 119988 238332 120040 238338
rect 119988 238274 120040 238280
rect 118712 219406 119752 219434
rect 118712 215286 118740 219406
rect 118700 215280 118752 215286
rect 118700 215222 118752 215228
rect 120184 202842 120212 250951
rect 120632 240236 120684 240242
rect 120632 240178 120684 240184
rect 120644 235822 120672 240178
rect 120736 239873 120764 275431
rect 121458 274816 121514 274825
rect 122116 274786 122144 319602
rect 122208 312730 122236 331842
rect 122196 312724 122248 312730
rect 122196 312666 122248 312672
rect 123496 294681 123524 372642
rect 123576 367124 123628 367130
rect 123576 367066 123628 367072
rect 123588 295322 123616 367066
rect 123668 364608 123720 364614
rect 123668 364550 123720 364556
rect 123576 295316 123628 295322
rect 123576 295258 123628 295264
rect 123680 295225 123708 364550
rect 123772 328506 123800 385086
rect 124128 378752 124180 378758
rect 124126 378720 124128 378729
rect 124180 378720 124182 378729
rect 124126 378655 124182 378664
rect 124232 350334 124260 458866
rect 124324 369850 124352 476070
rect 124416 392630 124444 493546
rect 124508 438190 124536 538834
rect 124600 460290 124628 552026
rect 125600 500336 125652 500342
rect 125600 500278 125652 500284
rect 124588 460284 124640 460290
rect 124588 460226 124640 460232
rect 125140 459604 125192 459610
rect 125140 459546 125192 459552
rect 125152 458930 125180 459546
rect 125140 458924 125192 458930
rect 125140 458866 125192 458872
rect 124496 438184 124548 438190
rect 124496 438126 124548 438132
rect 124404 392624 124456 392630
rect 124404 392566 124456 392572
rect 124404 386572 124456 386578
rect 124404 386514 124456 386520
rect 124312 369844 124364 369850
rect 124312 369786 124364 369792
rect 124220 350328 124272 350334
rect 124220 350270 124272 350276
rect 124232 345014 124260 350270
rect 124232 344986 124352 345014
rect 124324 331974 124352 344986
rect 124312 331968 124364 331974
rect 124312 331910 124364 331916
rect 124416 331906 124444 386514
rect 125612 386374 125640 500278
rect 125704 496262 125732 583743
rect 125876 567248 125928 567254
rect 125876 567190 125928 567196
rect 125784 545760 125836 545766
rect 125784 545702 125836 545708
rect 125692 496256 125744 496262
rect 125692 496198 125744 496204
rect 125690 491872 125746 491881
rect 125690 491807 125746 491816
rect 125704 392834 125732 491807
rect 125796 454034 125824 545702
rect 125888 476882 125916 567190
rect 126256 539034 126284 616830
rect 137296 585818 137324 700402
rect 137848 700398 137876 703520
rect 154132 700398 154160 703520
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 170324 697610 170352 703520
rect 202800 703390 202828 703520
rect 201500 703384 201552 703390
rect 201500 703326 201552 703332
rect 202788 703384 202840 703390
rect 202788 703326 202840 703332
rect 170312 697604 170364 697610
rect 170312 697546 170364 697552
rect 159364 643136 159416 643142
rect 159364 643078 159416 643084
rect 137284 585812 137336 585818
rect 137284 585754 137336 585760
rect 136822 581768 136878 581777
rect 136822 581703 136878 581712
rect 126980 581120 127032 581126
rect 126980 581062 127032 581068
rect 126244 539028 126296 539034
rect 126244 538970 126296 538976
rect 126992 491978 127020 581062
rect 128360 579760 128412 579766
rect 128360 579702 128412 579708
rect 127624 537736 127676 537742
rect 127624 537678 127676 537684
rect 127072 496256 127124 496262
rect 127072 496198 127124 496204
rect 126980 491972 127032 491978
rect 126980 491914 127032 491920
rect 125876 476876 125928 476882
rect 125876 476818 125928 476824
rect 125784 454028 125836 454034
rect 125784 453970 125836 453976
rect 125796 453937 125824 453970
rect 125782 453928 125838 453937
rect 125782 453863 125838 453872
rect 125888 398274 125916 476818
rect 125876 398268 125928 398274
rect 125876 398210 125928 398216
rect 127084 398206 127112 496198
rect 127256 494828 127308 494834
rect 127256 494770 127308 494776
rect 127072 398200 127124 398206
rect 127072 398142 127124 398148
rect 127164 396772 127216 396778
rect 127164 396714 127216 396720
rect 126336 394800 126388 394806
rect 126336 394742 126388 394748
rect 125692 392828 125744 392834
rect 125692 392770 125744 392776
rect 126244 386640 126296 386646
rect 126244 386582 126296 386588
rect 125600 386368 125652 386374
rect 125600 386310 125652 386316
rect 125692 385688 125744 385694
rect 125692 385630 125744 385636
rect 125600 381540 125652 381546
rect 125600 381482 125652 381488
rect 124956 368756 125008 368762
rect 124956 368698 125008 368704
rect 124404 331900 124456 331906
rect 124404 331842 124456 331848
rect 124312 331220 124364 331226
rect 124312 331162 124364 331168
rect 123760 328500 123812 328506
rect 123760 328442 123812 328448
rect 124128 328500 124180 328506
rect 124128 328442 124180 328448
rect 124140 327962 124168 328442
rect 124128 327956 124180 327962
rect 124128 327898 124180 327904
rect 123760 304020 123812 304026
rect 123760 303962 123812 303968
rect 123666 295216 123722 295225
rect 123666 295151 123722 295160
rect 123482 294672 123538 294681
rect 123482 294607 123538 294616
rect 123484 292800 123536 292806
rect 123484 292742 123536 292748
rect 122194 282296 122250 282305
rect 122194 282231 122250 282240
rect 121458 274751 121514 274760
rect 121552 274780 121604 274786
rect 121472 274718 121500 274751
rect 121552 274722 121604 274728
rect 122104 274780 122156 274786
rect 122104 274722 122156 274728
rect 121460 274712 121512 274718
rect 121460 274654 121512 274660
rect 121564 274145 121592 274722
rect 121550 274136 121606 274145
rect 121550 274071 121606 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273358 121500 273391
rect 121460 273352 121512 273358
rect 121460 273294 121512 273300
rect 121460 273216 121512 273222
rect 121460 273158 121512 273164
rect 121472 272785 121500 273158
rect 121458 272776 121514 272785
rect 121458 272711 121514 272720
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121458 270056 121514 270065
rect 121458 269991 121514 270000
rect 121472 269686 121500 269991
rect 121460 269680 121512 269686
rect 121460 269622 121512 269628
rect 121458 269376 121514 269385
rect 121458 269311 121514 269320
rect 121472 269142 121500 269311
rect 121460 269136 121512 269142
rect 121460 269078 121512 269084
rect 121552 269068 121604 269074
rect 121552 269010 121604 269016
rect 121564 268705 121592 269010
rect 121550 268696 121606 268705
rect 121550 268631 121606 268640
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267782 121500 267951
rect 121460 267776 121512 267782
rect 121460 267718 121512 267724
rect 121550 267336 121606 267345
rect 121550 267271 121606 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266490 121500 266591
rect 121460 266484 121512 266490
rect 121460 266426 121512 266432
rect 121564 266422 121592 267271
rect 121552 266416 121604 266422
rect 121552 266358 121604 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121460 264920 121512 264926
rect 121460 264862 121512 264868
rect 121472 264625 121500 264862
rect 121458 264616 121514 264625
rect 121458 264551 121514 264560
rect 121458 263936 121514 263945
rect 121458 263871 121514 263880
rect 121472 263634 121500 263871
rect 121460 263628 121512 263634
rect 121460 263570 121512 263576
rect 121552 263560 121604 263566
rect 121552 263502 121604 263508
rect 121460 263492 121512 263498
rect 121460 263434 121512 263440
rect 121472 263265 121500 263434
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121564 262585 121592 263502
rect 121550 262576 121606 262585
rect 121550 262511 121606 262520
rect 121552 262200 121604 262206
rect 121552 262142 121604 262148
rect 121460 262064 121512 262070
rect 121460 262006 121512 262012
rect 121472 261905 121500 262006
rect 121458 261896 121514 261905
rect 121458 261831 121514 261840
rect 121564 261225 121592 262142
rect 121550 261216 121606 261225
rect 121550 261151 121606 261160
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121552 259412 121604 259418
rect 121552 259354 121604 259360
rect 121564 258505 121592 259354
rect 121642 259176 121698 259185
rect 121642 259111 121698 259120
rect 121550 258496 121606 258505
rect 121550 258431 121606 258440
rect 121656 258126 121684 259111
rect 121644 258120 121696 258126
rect 122208 258074 122236 282231
rect 122746 278216 122802 278225
rect 122746 278151 122802 278160
rect 122760 277370 122788 278151
rect 122748 277364 122800 277370
rect 122748 277306 122800 277312
rect 122286 272096 122342 272105
rect 122286 272031 122342 272040
rect 122300 267734 122328 272031
rect 122300 267706 122512 267734
rect 121644 258062 121696 258068
rect 121460 258052 121512 258058
rect 121460 257994 121512 258000
rect 122116 258046 122236 258074
rect 121472 257145 121500 257994
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121460 256692 121512 256698
rect 121460 256634 121512 256640
rect 121472 255785 121500 256634
rect 121458 255776 121514 255785
rect 121458 255711 121514 255720
rect 121458 255096 121514 255105
rect 121458 255031 121514 255040
rect 121472 253978 121500 255031
rect 122116 254658 122144 258046
rect 122104 254652 122156 254658
rect 122104 254594 122156 254600
rect 122484 254590 122512 267706
rect 122472 254584 122524 254590
rect 122472 254526 122524 254532
rect 122102 254416 122158 254425
rect 122102 254351 122158 254360
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252686 121500 252991
rect 121460 252680 121512 252686
rect 121460 252622 121512 252628
rect 120816 252612 120868 252618
rect 120816 252554 120868 252560
rect 120722 239864 120778 239873
rect 120722 239799 120778 239808
rect 120828 239018 120856 252554
rect 121460 252544 121512 252550
rect 121460 252486 121512 252492
rect 121472 252385 121500 252486
rect 121458 252376 121514 252385
rect 121458 252311 121514 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121552 249756 121604 249762
rect 121552 249698 121604 249704
rect 121460 249688 121512 249694
rect 121564 249665 121592 249698
rect 121460 249630 121512 249636
rect 121550 249656 121606 249665
rect 121472 248985 121500 249630
rect 121550 249591 121606 249600
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247178 121500 248231
rect 121550 247616 121606 247625
rect 121550 247551 121606 247560
rect 121460 247172 121512 247178
rect 121460 247114 121512 247120
rect 121564 247110 121592 247551
rect 121552 247104 121604 247110
rect 121552 247046 121604 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121460 246200
rect 121512 246191 121514 246200
rect 121460 246162 121512 246168
rect 121564 245750 121592 246871
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121550 245576 121606 245585
rect 121550 245511 121606 245520
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121550 244216 121606 244225
rect 121472 243545 121500 244190
rect 121550 244151 121606 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121564 242962 121592 244151
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121458 242791 121514 242800
rect 121458 242176 121514 242185
rect 121458 242111 121514 242120
rect 121472 241534 121500 242111
rect 121460 241528 121512 241534
rect 121460 241470 121512 241476
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240310 121500 240751
rect 121460 240304 121512 240310
rect 121460 240246 121512 240252
rect 121458 240136 121514 240145
rect 121458 240071 121514 240080
rect 121472 239018 121500 240071
rect 120816 239012 120868 239018
rect 120816 238954 120868 238960
rect 121460 239012 121512 239018
rect 121460 238954 121512 238960
rect 120632 235816 120684 235822
rect 120632 235758 120684 235764
rect 120172 202836 120224 202842
rect 120172 202778 120224 202784
rect 118608 191140 118660 191146
rect 118608 191082 118660 191088
rect 114468 188420 114520 188426
rect 114468 188362 114520 188368
rect 110420 187128 110472 187134
rect 110420 187070 110472 187076
rect 122116 185842 122144 254351
rect 122194 253736 122250 253745
rect 122194 253671 122250 253680
rect 122208 206446 122236 253671
rect 122760 232529 122788 277306
rect 122746 232520 122802 232529
rect 122746 232455 122802 232464
rect 122196 206440 122248 206446
rect 122196 206382 122248 206388
rect 123496 195401 123524 292742
rect 123772 289746 123800 303962
rect 124128 292732 124180 292738
rect 124128 292674 124180 292680
rect 124140 292398 124168 292674
rect 124220 292460 124272 292466
rect 124220 292402 124272 292408
rect 124128 292392 124180 292398
rect 124128 292334 124180 292340
rect 124036 289876 124088 289882
rect 124036 289818 124088 289824
rect 124048 289746 124076 289818
rect 123760 289740 123812 289746
rect 123760 289682 123812 289688
rect 124036 289740 124088 289746
rect 124036 289682 124088 289688
rect 123576 289128 123628 289134
rect 123576 289070 123628 289076
rect 123588 238950 123616 289070
rect 123760 273284 123812 273290
rect 123760 273226 123812 273232
rect 123772 262070 123800 273226
rect 124140 264246 124168 292334
rect 124232 287026 124260 292402
rect 124220 287020 124272 287026
rect 124220 286962 124272 286968
rect 124324 286958 124352 331162
rect 124864 297016 124916 297022
rect 124864 296958 124916 296964
rect 124402 293176 124458 293185
rect 124402 293111 124458 293120
rect 124312 286952 124364 286958
rect 124312 286894 124364 286900
rect 124128 264240 124180 264246
rect 124128 264182 124180 264188
rect 123760 262064 123812 262070
rect 123760 262006 123812 262012
rect 123668 261520 123720 261526
rect 123668 261462 123720 261468
rect 123576 238944 123628 238950
rect 123576 238886 123628 238892
rect 123680 235929 123708 261462
rect 123760 244316 123812 244322
rect 123760 244258 123812 244264
rect 123666 235920 123722 235929
rect 123666 235855 123722 235864
rect 123772 226302 123800 244258
rect 124416 238882 124444 293111
rect 124404 238876 124456 238882
rect 124404 238818 124456 238824
rect 123760 226296 123812 226302
rect 123760 226238 123812 226244
rect 123482 195392 123538 195401
rect 123482 195327 123538 195336
rect 124876 188562 124904 296958
rect 124968 294914 124996 368698
rect 125048 365832 125100 365838
rect 125048 365774 125100 365780
rect 124956 294908 125008 294914
rect 124956 294850 125008 294856
rect 125060 294846 125088 365774
rect 125508 332580 125560 332586
rect 125508 332522 125560 332528
rect 125520 331809 125548 332522
rect 125506 331800 125562 331809
rect 125506 331735 125562 331744
rect 125612 300286 125640 381482
rect 125704 335306 125732 385630
rect 126060 382356 126112 382362
rect 126060 382298 126112 382304
rect 126072 381546 126100 382298
rect 126060 381540 126112 381546
rect 126060 381482 126112 381488
rect 125692 335300 125744 335306
rect 125692 335242 125744 335248
rect 125784 310480 125836 310486
rect 125784 310422 125836 310428
rect 125796 309233 125824 310422
rect 125782 309224 125838 309233
rect 125782 309159 125838 309168
rect 125600 300280 125652 300286
rect 125600 300222 125652 300228
rect 125598 300112 125654 300121
rect 125598 300047 125654 300056
rect 125048 294840 125100 294846
rect 125048 294782 125100 294788
rect 124956 282940 125008 282946
rect 124956 282882 125008 282888
rect 124968 271182 124996 282882
rect 124956 271176 125008 271182
rect 124956 271118 125008 271124
rect 124956 269680 125008 269686
rect 124956 269622 125008 269628
rect 124968 196654 124996 269622
rect 125612 264926 125640 300047
rect 126256 284238 126284 386582
rect 126348 363089 126376 394742
rect 126980 386436 127032 386442
rect 126980 386378 127032 386384
rect 126888 386368 126940 386374
rect 126888 386310 126940 386316
rect 126900 385762 126928 386310
rect 126888 385756 126940 385762
rect 126888 385698 126940 385704
rect 126334 363080 126390 363089
rect 126334 363015 126390 363024
rect 126886 363080 126942 363089
rect 126886 363015 126942 363024
rect 126794 343632 126850 343641
rect 126794 343567 126850 343576
rect 126808 342990 126836 343567
rect 126796 342984 126848 342990
rect 126794 342952 126796 342961
rect 126848 342952 126850 342961
rect 126794 342887 126850 342896
rect 126336 337816 126388 337822
rect 126336 337758 126388 337764
rect 126348 336870 126376 337758
rect 126336 336864 126388 336870
rect 126336 336806 126388 336812
rect 126244 284232 126296 284238
rect 126244 284174 126296 284180
rect 125600 264920 125652 264926
rect 125600 264862 125652 264868
rect 126244 256760 126296 256766
rect 126244 256702 126296 256708
rect 125048 246220 125100 246226
rect 125048 246162 125100 246168
rect 124956 196648 125008 196654
rect 124956 196590 125008 196596
rect 124864 188556 124916 188562
rect 124864 188498 124916 188504
rect 122104 185836 122156 185842
rect 122104 185778 122156 185784
rect 125060 185638 125088 246162
rect 126256 194070 126284 256702
rect 126348 237289 126376 336806
rect 126900 309126 126928 363015
rect 126888 309120 126940 309126
rect 126888 309062 126940 309068
rect 126426 291952 126482 291961
rect 126426 291887 126482 291896
rect 126334 237280 126390 237289
rect 126334 237215 126390 237224
rect 126348 226273 126376 237215
rect 126334 226264 126390 226273
rect 126334 226199 126390 226208
rect 126440 211886 126468 291887
rect 126992 237318 127020 386378
rect 127176 342922 127204 396714
rect 127268 395486 127296 494770
rect 127636 444514 127664 537678
rect 128372 534886 128400 579702
rect 134156 578264 134208 578270
rect 134156 578206 134208 578212
rect 129832 576904 129884 576910
rect 129832 576846 129884 576852
rect 129004 568608 129056 568614
rect 129004 568550 129056 568556
rect 128544 536172 128596 536178
rect 128544 536114 128596 536120
rect 128360 534880 128412 534886
rect 128360 534822 128412 534828
rect 128360 529236 128412 529242
rect 128360 529178 128412 529184
rect 128372 459610 128400 529178
rect 128452 493400 128504 493406
rect 128452 493342 128504 493348
rect 128360 459604 128412 459610
rect 128360 459546 128412 459552
rect 127624 444508 127676 444514
rect 127624 444450 127676 444456
rect 127636 443057 127664 444450
rect 127622 443048 127678 443057
rect 127622 442983 127678 442992
rect 127348 399492 127400 399498
rect 127348 399434 127400 399440
rect 127256 395480 127308 395486
rect 127256 395422 127308 395428
rect 127164 342916 127216 342922
rect 127164 342858 127216 342864
rect 127360 335238 127388 399434
rect 128464 395350 128492 493342
rect 128556 439006 128584 536114
rect 129016 478922 129044 568550
rect 129740 541680 129792 541686
rect 129740 541622 129792 541628
rect 129752 541074 129780 541622
rect 129740 541068 129792 541074
rect 129740 541010 129792 541016
rect 129004 478916 129056 478922
rect 129004 478858 129056 478864
rect 128636 463752 128688 463758
rect 128636 463694 128688 463700
rect 128544 439000 128596 439006
rect 128544 438942 128596 438948
rect 128544 405068 128596 405074
rect 128544 405010 128596 405016
rect 128452 395344 128504 395350
rect 128452 395286 128504 395292
rect 127624 382288 127676 382294
rect 127624 382230 127676 382236
rect 127636 368490 127664 382230
rect 127624 368484 127676 368490
rect 127624 368426 127676 368432
rect 127348 335232 127400 335238
rect 127348 335174 127400 335180
rect 127360 334014 127388 335174
rect 127348 334008 127400 334014
rect 127348 333950 127400 333956
rect 127636 332042 127664 368426
rect 128360 334008 128412 334014
rect 128360 333950 128412 333956
rect 127624 332036 127676 332042
rect 127624 331978 127676 331984
rect 128268 322924 128320 322930
rect 128268 322866 128320 322872
rect 127624 292936 127676 292942
rect 127624 292878 127676 292884
rect 126980 237312 127032 237318
rect 126980 237254 127032 237260
rect 127636 213314 127664 292878
rect 128280 262274 128308 322866
rect 128372 289134 128400 333950
rect 128556 333946 128584 405010
rect 128648 354686 128676 463694
rect 129752 444446 129780 541010
rect 129844 499574 129872 576846
rect 131120 575612 131172 575618
rect 131120 575554 131172 575560
rect 130384 573368 130436 573374
rect 130384 573310 130436 573316
rect 129844 499546 129964 499574
rect 129936 487218 129964 499546
rect 129924 487212 129976 487218
rect 129924 487154 129976 487160
rect 129832 481772 129884 481778
rect 129832 481714 129884 481720
rect 129844 481642 129872 481714
rect 129832 481636 129884 481642
rect 129832 481578 129884 481584
rect 129832 478916 129884 478922
rect 129832 478858 129884 478864
rect 129844 476814 129872 478858
rect 129832 476808 129884 476814
rect 129832 476750 129884 476756
rect 129740 444440 129792 444446
rect 129740 444382 129792 444388
rect 129004 393984 129056 393990
rect 129004 393926 129056 393932
rect 128636 354680 128688 354686
rect 128636 354622 128688 354628
rect 128648 354074 128676 354622
rect 128636 354068 128688 354074
rect 128636 354010 128688 354016
rect 129016 336802 129044 393926
rect 129096 360256 129148 360262
rect 129096 360198 129148 360204
rect 129108 340814 129136 360198
rect 129096 340808 129148 340814
rect 129096 340750 129148 340756
rect 129752 336870 129780 444382
rect 129844 370598 129872 476750
rect 129936 382362 129964 487154
rect 130396 481778 130424 573310
rect 131132 485081 131160 575554
rect 133880 571396 133932 571402
rect 133880 571338 133932 571344
rect 133144 564460 133196 564466
rect 133144 564402 133196 564408
rect 132500 549364 132552 549370
rect 132500 549306 132552 549312
rect 131212 536104 131264 536110
rect 131212 536046 131264 536052
rect 131118 485072 131174 485081
rect 131118 485007 131174 485016
rect 130384 481772 130436 481778
rect 130384 481714 130436 481720
rect 131224 451274 131252 536046
rect 131304 497480 131356 497486
rect 131304 497422 131356 497428
rect 131132 451246 131252 451274
rect 131132 448594 131160 451246
rect 131120 448588 131172 448594
rect 131120 448530 131172 448536
rect 130016 387116 130068 387122
rect 130016 387058 130068 387064
rect 129924 382356 129976 382362
rect 129924 382298 129976 382304
rect 129832 370592 129884 370598
rect 129832 370534 129884 370540
rect 129740 336864 129792 336870
rect 129740 336806 129792 336812
rect 129004 336796 129056 336802
rect 129004 336738 129056 336744
rect 128544 333940 128596 333946
rect 128544 333882 128596 333888
rect 128634 318744 128690 318753
rect 128634 318679 128690 318688
rect 128648 317558 128676 318679
rect 128636 317552 128688 317558
rect 128636 317494 128688 317500
rect 129096 313336 129148 313342
rect 129096 313278 129148 313284
rect 129004 296880 129056 296886
rect 129004 296822 129056 296828
rect 128360 289128 128412 289134
rect 128360 289070 128412 289076
rect 128268 262268 128320 262274
rect 128268 262210 128320 262216
rect 127624 213308 127676 213314
rect 127624 213250 127676 213256
rect 126428 211880 126480 211886
rect 126428 211822 126480 211828
rect 126244 194064 126296 194070
rect 126244 194006 126296 194012
rect 129016 191185 129044 296822
rect 129108 249694 129136 313278
rect 129740 298784 129792 298790
rect 129740 298726 129792 298732
rect 129280 290488 129332 290494
rect 129280 290430 129332 290436
rect 129188 280220 129240 280226
rect 129188 280162 129240 280168
rect 129096 249688 129148 249694
rect 129096 249630 129148 249636
rect 129002 191176 129058 191185
rect 129002 191111 129058 191120
rect 129200 191049 129228 280162
rect 129292 235890 129320 290430
rect 129752 288425 129780 298726
rect 129844 292398 129872 370534
rect 130028 361554 130056 387058
rect 130016 361548 130068 361554
rect 130016 361490 130068 361496
rect 130028 360262 130056 361490
rect 130016 360256 130068 360262
rect 130016 360198 130068 360204
rect 131132 336598 131160 448530
rect 131316 437238 131344 497422
rect 132512 456142 132540 549306
rect 132592 537532 132644 537538
rect 132592 537474 132644 537480
rect 132500 456136 132552 456142
rect 132500 456078 132552 456084
rect 131304 437232 131356 437238
rect 131304 437174 131356 437180
rect 131304 401056 131356 401062
rect 131304 400998 131356 401004
rect 131212 396840 131264 396846
rect 131212 396782 131264 396788
rect 131224 338094 131252 396782
rect 131212 338088 131264 338094
rect 131212 338030 131264 338036
rect 131224 337414 131252 338030
rect 131212 337408 131264 337414
rect 131212 337350 131264 337356
rect 131120 336592 131172 336598
rect 131120 336534 131172 336540
rect 131212 334620 131264 334626
rect 131212 334562 131264 334568
rect 131120 330540 131172 330546
rect 131120 330482 131172 330488
rect 130568 303000 130620 303006
rect 130568 302942 130620 302948
rect 130476 292868 130528 292874
rect 130476 292810 130528 292816
rect 129832 292392 129884 292398
rect 129832 292334 129884 292340
rect 129738 288416 129794 288425
rect 129738 288351 129794 288360
rect 130384 254652 130436 254658
rect 130384 254594 130436 254600
rect 129280 235884 129332 235890
rect 129280 235826 129332 235832
rect 129186 191040 129242 191049
rect 129186 190975 129242 190984
rect 125048 185632 125100 185638
rect 125048 185574 125100 185580
rect 125508 183592 125560 183598
rect 125508 183534 125560 183540
rect 109040 182844 109092 182850
rect 109040 182786 109092 182792
rect 110696 182368 110748 182374
rect 110696 182310 110748 182316
rect 110328 178288 110380 178294
rect 110328 178230 110380 178236
rect 102046 177712 102102 177721
rect 102046 177647 102102 177656
rect 105726 177712 105782 177721
rect 105726 177647 105782 177656
rect 107566 177712 107622 177721
rect 107566 177647 107622 177656
rect 108120 176996 108172 177002
rect 108120 176938 108172 176944
rect 103336 176928 103388 176934
rect 103336 176870 103388 176876
rect 103348 176769 103376 176870
rect 104624 176792 104676 176798
rect 98734 176760 98790 176769
rect 98734 176695 98790 176704
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 104622 176760 104624 176769
rect 108132 176769 108160 176938
rect 110340 176769 110368 178230
rect 110708 177721 110736 182310
rect 112444 182300 112496 182306
rect 112444 182242 112496 182248
rect 112456 177721 112484 182242
rect 119528 182232 119580 182238
rect 119528 182174 119580 182180
rect 118424 180872 118476 180878
rect 118424 180814 118476 180820
rect 115848 179512 115900 179518
rect 115848 179454 115900 179460
rect 113732 178220 113784 178226
rect 113732 178162 113784 178168
rect 110694 177712 110750 177721
rect 110694 177647 110750 177656
rect 112442 177712 112498 177721
rect 112442 177647 112498 177656
rect 113744 176769 113772 178162
rect 115860 177041 115888 179454
rect 118436 177721 118464 180814
rect 119540 177721 119568 182174
rect 124036 180940 124088 180946
rect 124036 180882 124088 180888
rect 124048 177721 124076 180882
rect 125520 177721 125548 183534
rect 129464 181008 129516 181014
rect 129464 180950 129516 180956
rect 126612 179580 126664 179586
rect 126612 179522 126664 179528
rect 118422 177712 118478 177721
rect 118422 177647 118478 177656
rect 119526 177712 119582 177721
rect 119526 177647 119582 177656
rect 124034 177712 124090 177721
rect 124034 177647 124090 177656
rect 125506 177712 125562 177721
rect 125506 177647 125562 177656
rect 126624 177041 126652 179522
rect 127072 178152 127124 178158
rect 127072 178094 127124 178100
rect 115846 177032 115902 177041
rect 115846 176967 115902 176976
rect 126610 177032 126666 177041
rect 126610 176967 126666 176976
rect 127084 176769 127112 178094
rect 129476 177721 129504 180950
rect 130396 178673 130424 254594
rect 130488 217394 130516 292810
rect 130580 251297 130608 302942
rect 130566 251288 130622 251297
rect 130566 251223 130622 251232
rect 130580 238746 130608 251223
rect 130568 238740 130620 238746
rect 130568 238682 130620 238688
rect 131132 235754 131160 330482
rect 131224 244254 131252 334562
rect 131316 317422 131344 400998
rect 132512 347750 132540 456078
rect 132604 441590 132632 537474
rect 133156 473346 133184 564402
rect 133892 479534 133920 571338
rect 133972 545216 134024 545222
rect 133972 545158 134024 545164
rect 133880 479528 133932 479534
rect 133880 479470 133932 479476
rect 133144 473340 133196 473346
rect 133144 473282 133196 473288
rect 133788 473340 133840 473346
rect 133788 473282 133840 473288
rect 133800 472666 133828 473282
rect 133788 472660 133840 472666
rect 133788 472602 133840 472608
rect 133788 466540 133840 466546
rect 133788 466482 133840 466488
rect 133800 466410 133828 466482
rect 133788 466404 133840 466410
rect 133788 466346 133840 466352
rect 132592 441584 132644 441590
rect 132592 441526 132644 441532
rect 132604 440366 132632 441526
rect 132592 440360 132644 440366
rect 132592 440302 132644 440308
rect 132592 405000 132644 405006
rect 132592 404942 132644 404948
rect 132500 347744 132552 347750
rect 132500 347686 132552 347692
rect 132500 339516 132552 339522
rect 132500 339458 132552 339464
rect 131304 317416 131356 317422
rect 131304 317358 131356 317364
rect 131488 317416 131540 317422
rect 131488 317358 131540 317364
rect 131500 316878 131528 317358
rect 131488 316872 131540 316878
rect 131488 316814 131540 316820
rect 131304 309120 131356 309126
rect 131304 309062 131356 309068
rect 131316 284306 131344 309062
rect 131304 284300 131356 284306
rect 131304 284242 131356 284248
rect 132512 277302 132540 339458
rect 132604 333878 132632 404942
rect 132684 391264 132736 391270
rect 132684 391206 132736 391212
rect 133696 391264 133748 391270
rect 133696 391206 133748 391212
rect 132696 339318 132724 391206
rect 133708 390590 133736 391206
rect 133696 390584 133748 390590
rect 133696 390526 133748 390532
rect 133800 360126 133828 466346
rect 133892 375358 133920 479470
rect 133984 452606 134012 545158
rect 134064 494760 134116 494766
rect 134064 494702 134116 494708
rect 133972 452600 134024 452606
rect 133972 452542 134024 452548
rect 133972 440360 134024 440366
rect 133972 440302 134024 440308
rect 133880 375352 133932 375358
rect 133880 375294 133932 375300
rect 133788 360120 133840 360126
rect 133788 360062 133840 360068
rect 133800 359514 133828 360062
rect 133788 359508 133840 359514
rect 133788 359450 133840 359456
rect 133788 347744 133840 347750
rect 133788 347686 133840 347692
rect 133800 347070 133828 347686
rect 133788 347064 133840 347070
rect 133788 347006 133840 347012
rect 132960 340196 133012 340202
rect 132960 340138 133012 340144
rect 132972 339522 133000 340138
rect 132960 339516 133012 339522
rect 132960 339458 133012 339464
rect 132684 339312 132736 339318
rect 132684 339254 132736 339260
rect 133880 337408 133932 337414
rect 133880 337350 133932 337356
rect 132592 333872 132644 333878
rect 132592 333814 132644 333820
rect 133236 300960 133288 300966
rect 133236 300902 133288 300908
rect 133144 298852 133196 298858
rect 133144 298794 133196 298800
rect 132592 282940 132644 282946
rect 132592 282882 132644 282888
rect 132500 277296 132552 277302
rect 132500 277238 132552 277244
rect 131764 259480 131816 259486
rect 131764 259422 131816 259428
rect 131212 244248 131264 244254
rect 131212 244190 131264 244196
rect 131120 235748 131172 235754
rect 131120 235690 131172 235696
rect 130476 217388 130528 217394
rect 130476 217330 130528 217336
rect 131776 185774 131804 259422
rect 132604 233102 132632 282882
rect 132592 233096 132644 233102
rect 132592 233038 132644 233044
rect 133156 199578 133184 298794
rect 133248 273970 133276 300902
rect 133604 284232 133656 284238
rect 133604 284174 133656 284180
rect 133616 282946 133644 284174
rect 133604 282940 133656 282946
rect 133604 282882 133656 282888
rect 133236 273964 133288 273970
rect 133236 273906 133288 273912
rect 133892 273222 133920 337350
rect 133984 336666 134012 440302
rect 134076 392698 134104 494702
rect 134168 489190 134196 578206
rect 136640 559564 136692 559570
rect 136640 559506 136692 559512
rect 135444 559020 135496 559026
rect 135444 558962 135496 558968
rect 135260 546508 135312 546514
rect 135260 546450 135312 546456
rect 134156 489184 134208 489190
rect 134156 489126 134208 489132
rect 135272 456074 135300 546450
rect 135352 496120 135404 496126
rect 135352 496062 135404 496068
rect 135260 456068 135312 456074
rect 135260 456010 135312 456016
rect 135168 452600 135220 452606
rect 135168 452542 135220 452548
rect 135180 451926 135208 452542
rect 135168 451920 135220 451926
rect 135168 451862 135220 451868
rect 135260 445868 135312 445874
rect 135260 445810 135312 445816
rect 134708 396024 134760 396030
rect 134708 395966 134760 395972
rect 134720 395350 134748 395966
rect 134708 395344 134760 395350
rect 134708 395286 134760 395292
rect 134720 394913 134748 395286
rect 134706 394904 134762 394913
rect 134706 394839 134762 394848
rect 134156 393440 134208 393446
rect 134156 393382 134208 393388
rect 134064 392692 134116 392698
rect 134064 392634 134116 392640
rect 134076 392154 134104 392634
rect 134064 392148 134116 392154
rect 134064 392090 134116 392096
rect 133972 336660 134024 336666
rect 133972 336602 134024 336608
rect 134168 322930 134196 393382
rect 135168 375352 135220 375358
rect 135168 375294 135220 375300
rect 135180 374649 135208 375294
rect 135166 374640 135222 374649
rect 135166 374575 135222 374584
rect 135272 339250 135300 445810
rect 135364 389910 135392 496062
rect 135456 468518 135484 558962
rect 136652 558958 136680 559506
rect 136640 558952 136692 558958
rect 136640 558894 136692 558900
rect 135444 468512 135496 468518
rect 135444 468454 135496 468460
rect 136652 466410 136680 558894
rect 136732 542428 136784 542434
rect 136732 542370 136784 542376
rect 136640 466404 136692 466410
rect 136640 466346 136692 466352
rect 136744 452538 136772 542370
rect 136836 500274 136864 581703
rect 142160 569968 142212 569974
rect 142160 569910 142212 569916
rect 138020 563712 138072 563718
rect 138020 563654 138072 563660
rect 136824 500268 136876 500274
rect 136824 500210 136876 500216
rect 137100 500268 137152 500274
rect 137100 500210 137152 500216
rect 137112 499633 137140 500210
rect 137098 499624 137154 499633
rect 137098 499559 137154 499568
rect 137284 493332 137336 493338
rect 137284 493274 137336 493280
rect 136732 452532 136784 452538
rect 136732 452474 136784 452480
rect 136732 440292 136784 440298
rect 136732 440234 136784 440240
rect 135444 394052 135496 394058
rect 135444 393994 135496 394000
rect 135456 393446 135484 393994
rect 135444 393440 135496 393446
rect 135444 393382 135496 393388
rect 135352 389904 135404 389910
rect 135352 389846 135404 389852
rect 135260 339244 135312 339250
rect 135260 339186 135312 339192
rect 135456 335170 135484 393382
rect 136640 390652 136692 390658
rect 136640 390594 136692 390600
rect 136548 389904 136600 389910
rect 136546 389872 136548 389881
rect 136600 389872 136602 389881
rect 136546 389807 136602 389816
rect 135904 385076 135956 385082
rect 135904 385018 135956 385024
rect 135444 335164 135496 335170
rect 135444 335106 135496 335112
rect 134156 322924 134208 322930
rect 134156 322866 134208 322872
rect 134524 320952 134576 320958
rect 134524 320894 134576 320900
rect 133880 273216 133932 273222
rect 133880 273158 133932 273164
rect 133236 269136 133288 269142
rect 133236 269078 133288 269084
rect 133144 199572 133196 199578
rect 133144 199514 133196 199520
rect 131764 185768 131816 185774
rect 131764 185710 131816 185716
rect 132408 182436 132460 182442
rect 132408 182378 132460 182384
rect 130382 178664 130438 178673
rect 130382 178599 130438 178608
rect 132420 177721 132448 182378
rect 133248 181393 133276 269078
rect 133892 256766 133920 256797
rect 133880 256760 133932 256766
rect 133878 256728 133880 256737
rect 133932 256728 133934 256737
rect 133878 256663 133934 256672
rect 133328 249824 133380 249830
rect 133328 249766 133380 249772
rect 133340 183054 133368 249766
rect 133892 237250 133920 256663
rect 133880 237244 133932 237250
rect 133880 237186 133932 237192
rect 134536 185910 134564 320894
rect 134616 304292 134668 304298
rect 134616 304234 134668 304240
rect 134628 242894 134656 304234
rect 134800 295452 134852 295458
rect 134800 295394 134852 295400
rect 134812 268394 134840 295394
rect 134800 268388 134852 268394
rect 134800 268330 134852 268336
rect 134708 267776 134760 267782
rect 134708 267718 134760 267724
rect 134616 242888 134668 242894
rect 134616 242830 134668 242836
rect 134720 234598 134748 267718
rect 135916 246566 135944 385018
rect 135996 307148 136048 307154
rect 135996 307090 136048 307096
rect 135904 246560 135956 246566
rect 135904 246502 135956 246508
rect 135168 243024 135220 243030
rect 135168 242966 135220 242972
rect 135180 242894 135208 242966
rect 135168 242888 135220 242894
rect 135168 242830 135220 242836
rect 134708 234592 134760 234598
rect 134708 234534 134760 234540
rect 136008 189922 136036 307090
rect 136088 299736 136140 299742
rect 136088 299678 136140 299684
rect 136100 210594 136128 299678
rect 136652 259418 136680 390594
rect 136744 314634 136772 440234
rect 136824 392148 136876 392154
rect 136824 392090 136876 392096
rect 136836 315314 136864 392090
rect 137296 390658 137324 493274
rect 138032 470558 138060 563654
rect 140780 560312 140832 560318
rect 140780 560254 140832 560260
rect 138112 550656 138164 550662
rect 138112 550598 138164 550604
rect 138020 470552 138072 470558
rect 138020 470494 138072 470500
rect 138032 469266 138060 470494
rect 138020 469260 138072 469266
rect 138020 469202 138072 469208
rect 138124 460222 138152 550598
rect 139492 545148 139544 545154
rect 139492 545090 139544 545096
rect 139400 491972 139452 491978
rect 139400 491914 139452 491920
rect 138204 469260 138256 469266
rect 138204 469202 138256 469208
rect 138112 460216 138164 460222
rect 138112 460158 138164 460164
rect 138112 458244 138164 458250
rect 138112 458186 138164 458192
rect 137376 452532 137428 452538
rect 137376 452474 137428 452480
rect 137388 451314 137416 452474
rect 137376 451308 137428 451314
rect 137376 451250 137428 451256
rect 137284 390652 137336 390658
rect 137284 390594 137336 390600
rect 137296 389366 137324 390594
rect 137284 389360 137336 389366
rect 137284 389302 137336 389308
rect 137388 373726 137416 451250
rect 138020 393508 138072 393514
rect 138020 393450 138072 393456
rect 137376 373720 137428 373726
rect 137376 373662 137428 373668
rect 137284 354000 137336 354006
rect 137282 353968 137284 353977
rect 137336 353968 137338 353977
rect 137282 353903 137338 353912
rect 136824 315308 136876 315314
rect 136824 315250 136876 315256
rect 136732 314628 136784 314634
rect 136732 314570 136784 314576
rect 136744 313954 136772 314570
rect 136732 313948 136784 313954
rect 136732 313890 136784 313896
rect 136732 305788 136784 305794
rect 136732 305730 136784 305736
rect 136640 259412 136692 259418
rect 136640 259354 136692 259360
rect 136744 256698 136772 305730
rect 137284 301640 137336 301646
rect 137284 301582 137336 301588
rect 137100 259412 137152 259418
rect 137100 259354 137152 259360
rect 137112 258738 137140 259354
rect 137100 258732 137152 258738
rect 137100 258674 137152 258680
rect 136732 256692 136784 256698
rect 136732 256634 136784 256640
rect 136744 256086 136772 256634
rect 136732 256080 136784 256086
rect 136732 256022 136784 256028
rect 136640 246560 136692 246566
rect 136640 246502 136692 246508
rect 136652 245682 136680 246502
rect 136640 245676 136692 245682
rect 136640 245618 136692 245624
rect 136652 231742 136680 245618
rect 136640 231736 136692 231742
rect 136640 231678 136692 231684
rect 136088 210588 136140 210594
rect 136088 210530 136140 210536
rect 137296 202298 137324 301582
rect 138032 261526 138060 393450
rect 138124 345030 138152 458186
rect 138216 365702 138244 469202
rect 139412 392766 139440 491914
rect 139504 454714 139532 545090
rect 140792 469878 140820 560254
rect 141516 554056 141568 554062
rect 141516 553998 141568 554004
rect 141528 553450 141556 553998
rect 141516 553444 141568 553450
rect 141516 553386 141568 553392
rect 142068 553444 142120 553450
rect 142068 553386 142120 553392
rect 141056 485852 141108 485858
rect 141056 485794 141108 485800
rect 140964 469940 141016 469946
rect 140964 469882 141016 469888
rect 140780 469872 140832 469878
rect 140780 469814 140832 469820
rect 140778 462360 140834 462369
rect 140778 462295 140780 462304
rect 140832 462295 140834 462304
rect 140780 462266 140832 462272
rect 139492 454708 139544 454714
rect 139492 454650 139544 454656
rect 139492 448520 139544 448526
rect 139492 448462 139544 448468
rect 140688 448520 140740 448526
rect 140688 448462 140740 448468
rect 139504 447846 139532 448462
rect 139492 447840 139544 447846
rect 139492 447782 139544 447788
rect 139400 392760 139452 392766
rect 139400 392702 139452 392708
rect 139400 383716 139452 383722
rect 139400 383658 139452 383664
rect 138296 373720 138348 373726
rect 138296 373662 138348 373668
rect 138308 372638 138336 373662
rect 138296 372632 138348 372638
rect 138296 372574 138348 372580
rect 138204 365696 138256 365702
rect 138204 365638 138256 365644
rect 138112 345024 138164 345030
rect 138112 344966 138164 344972
rect 138124 344350 138152 344966
rect 138112 344344 138164 344350
rect 138112 344286 138164 344292
rect 138308 340882 138336 372574
rect 138296 340876 138348 340882
rect 138296 340818 138348 340824
rect 138112 336796 138164 336802
rect 138112 336738 138164 336744
rect 138124 263498 138152 336738
rect 138664 308576 138716 308582
rect 138664 308518 138716 308524
rect 138112 263492 138164 263498
rect 138112 263434 138164 263440
rect 138124 263090 138152 263434
rect 138112 263084 138164 263090
rect 138112 263026 138164 263032
rect 138020 261520 138072 261526
rect 138020 261462 138072 261468
rect 137468 258120 137520 258126
rect 137468 258062 137520 258068
rect 137376 247172 137428 247178
rect 137376 247114 137428 247120
rect 137284 202292 137336 202298
rect 137284 202234 137336 202240
rect 135996 189916 136048 189922
rect 135996 189858 136048 189864
rect 137388 187202 137416 247114
rect 137480 244934 137508 258062
rect 137468 244928 137520 244934
rect 137468 244870 137520 244876
rect 138676 196722 138704 308518
rect 139412 300218 139440 383658
rect 140700 374338 140728 448462
rect 140872 444508 140924 444514
rect 140872 444450 140924 444456
rect 140780 390652 140832 390658
rect 140780 390594 140832 390600
rect 140044 374332 140096 374338
rect 140044 374274 140096 374280
rect 140688 374332 140740 374338
rect 140688 374274 140740 374280
rect 140056 337958 140084 374274
rect 140700 374066 140728 374274
rect 140688 374060 140740 374066
rect 140688 374002 140740 374008
rect 140044 337952 140096 337958
rect 140044 337894 140096 337900
rect 140226 322144 140282 322153
rect 140226 322079 140282 322088
rect 140044 303068 140096 303074
rect 140044 303010 140096 303016
rect 139400 300212 139452 300218
rect 139400 300154 139452 300160
rect 138756 263628 138808 263634
rect 138756 263570 138808 263576
rect 138664 196716 138716 196722
rect 138664 196658 138716 196664
rect 138768 189854 138796 263570
rect 140056 205154 140084 303010
rect 140136 295724 140188 295730
rect 140136 295666 140188 295672
rect 140148 218754 140176 295666
rect 140240 249830 140268 322079
rect 140228 249824 140280 249830
rect 140228 249766 140280 249772
rect 140686 242856 140742 242865
rect 140686 242791 140742 242800
rect 140700 241534 140728 242791
rect 140688 241528 140740 241534
rect 140688 241470 140740 241476
rect 140700 234433 140728 241470
rect 140686 234424 140742 234433
rect 140686 234359 140742 234368
rect 140136 218748 140188 218754
rect 140136 218690 140188 218696
rect 140792 218006 140820 390594
rect 140884 327078 140912 444450
rect 140976 362914 141004 469882
rect 141068 382226 141096 485794
rect 142080 462369 142108 553386
rect 142172 477494 142200 569910
rect 155224 564460 155276 564466
rect 155224 564402 155276 564408
rect 142252 549296 142304 549302
rect 142252 549238 142304 549244
rect 142160 477488 142212 477494
rect 142160 477430 142212 477436
rect 142160 472660 142212 472666
rect 142160 472602 142212 472608
rect 142066 462360 142122 462369
rect 142066 462295 142122 462304
rect 141056 382220 141108 382226
rect 141056 382162 141108 382168
rect 141068 381614 141096 382162
rect 141056 381608 141108 381614
rect 141056 381550 141108 381556
rect 142172 367062 142200 472602
rect 142264 458862 142292 549238
rect 142344 541000 142396 541006
rect 142344 540942 142396 540948
rect 142252 458856 142304 458862
rect 142252 458798 142304 458804
rect 142252 456068 142304 456074
rect 142252 456010 142304 456016
rect 142160 367056 142212 367062
rect 142160 366998 142212 367004
rect 140964 362908 141016 362914
rect 140964 362850 141016 362856
rect 140976 362234 141004 362850
rect 140964 362228 141016 362234
rect 140964 362170 141016 362176
rect 142160 354000 142212 354006
rect 142160 353942 142212 353948
rect 141424 327820 141476 327826
rect 141424 327762 141476 327768
rect 140872 327072 140924 327078
rect 140872 327014 140924 327020
rect 140884 326466 140912 327014
rect 140872 326460 140924 326466
rect 140872 326402 140924 326408
rect 140780 218000 140832 218006
rect 140780 217942 140832 217948
rect 140044 205148 140096 205154
rect 140044 205090 140096 205096
rect 141436 192778 141464 327762
rect 141516 295656 141568 295662
rect 141516 295598 141568 295604
rect 141528 200870 141556 295598
rect 141608 263084 141660 263090
rect 141608 263026 141660 263032
rect 141620 256018 141648 263026
rect 141608 256012 141660 256018
rect 141608 255954 141660 255960
rect 142172 235958 142200 353942
rect 142264 346390 142292 456010
rect 142356 448526 142384 540942
rect 155236 538218 155264 564402
rect 159376 554062 159404 643078
rect 201512 559570 201540 703326
rect 218992 698970 219020 703520
rect 235184 700330 235212 703520
rect 267660 703322 267688 703520
rect 267648 703316 267700 703322
rect 267648 703258 267700 703264
rect 283852 700330 283880 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 238024 700324 238076 700330
rect 238024 700266 238076 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 218980 698964 219032 698970
rect 218980 698906 219032 698912
rect 238036 594114 238064 700266
rect 276664 630692 276716 630698
rect 276664 630634 276716 630640
rect 238024 594108 238076 594114
rect 238024 594050 238076 594056
rect 201500 559564 201552 559570
rect 201500 559506 201552 559512
rect 159364 554056 159416 554062
rect 159364 553998 159416 554004
rect 155224 538212 155276 538218
rect 155224 538154 155276 538160
rect 151820 489184 151872 489190
rect 151820 489126 151872 489132
rect 143724 481772 143776 481778
rect 143724 481714 143776 481720
rect 143632 456816 143684 456822
rect 143632 456758 143684 456764
rect 142344 448520 142396 448526
rect 142344 448462 142396 448468
rect 143540 445800 143592 445806
rect 143540 445742 143592 445748
rect 142344 395480 142396 395486
rect 142344 395422 142396 395428
rect 142252 346384 142304 346390
rect 142252 346326 142304 346332
rect 142250 338056 142306 338065
rect 142250 337991 142252 338000
rect 142304 337991 142306 338000
rect 142252 337962 142304 337968
rect 142356 288318 142384 395422
rect 142804 371884 142856 371890
rect 142804 371826 142856 371832
rect 142816 356726 142844 371826
rect 142436 356720 142488 356726
rect 142436 356662 142488 356668
rect 142804 356720 142856 356726
rect 142804 356662 142856 356668
rect 142448 290494 142476 356662
rect 143448 346384 143500 346390
rect 143448 346326 143500 346332
rect 143460 345681 143488 346326
rect 143446 345672 143502 345681
rect 143446 345607 143502 345616
rect 143448 338020 143500 338026
rect 143448 337962 143500 337968
rect 143460 336802 143488 337962
rect 143448 336796 143500 336802
rect 143448 336738 143500 336744
rect 143552 318782 143580 445742
rect 143644 345710 143672 456758
rect 143736 376038 143764 481714
rect 146300 481704 146352 481710
rect 146300 481646 146352 481652
rect 145012 471300 145064 471306
rect 145012 471242 145064 471248
rect 145024 470626 145052 471242
rect 145012 470620 145064 470626
rect 145012 470562 145064 470568
rect 144920 466472 144972 466478
rect 144920 466414 144972 466420
rect 143816 389836 143868 389842
rect 143816 389778 143868 389784
rect 143724 376032 143776 376038
rect 143724 375974 143776 375980
rect 143724 359508 143776 359514
rect 143724 359450 143776 359456
rect 143632 345704 143684 345710
rect 143632 345646 143684 345652
rect 143540 318776 143592 318782
rect 143540 318718 143592 318724
rect 142804 305720 142856 305726
rect 142804 305662 142856 305668
rect 142436 290488 142488 290494
rect 142436 290430 142488 290436
rect 142344 288312 142396 288318
rect 142344 288254 142396 288260
rect 142160 235952 142212 235958
rect 142160 235894 142212 235900
rect 141516 200864 141568 200870
rect 141516 200806 141568 200812
rect 142816 193934 142844 305662
rect 143448 288312 143500 288318
rect 143448 288254 143500 288260
rect 143460 287706 143488 288254
rect 143448 287700 143500 287706
rect 143448 287642 143500 287648
rect 143736 286890 143764 359450
rect 143828 301578 143856 389778
rect 143906 389056 143962 389065
rect 143906 388991 143962 389000
rect 143920 388074 143948 388991
rect 143908 388068 143960 388074
rect 143908 388010 143960 388016
rect 144932 357406 144960 466414
rect 145024 365022 145052 470562
rect 146312 376718 146340 481646
rect 146392 472048 146444 472054
rect 146392 471990 146444 471996
rect 146300 376712 146352 376718
rect 146300 376654 146352 376660
rect 146300 367056 146352 367062
rect 146300 366998 146352 367004
rect 145012 365016 145064 365022
rect 145012 364958 145064 364964
rect 144920 357400 144972 357406
rect 144920 357342 144972 357348
rect 144920 352504 144972 352510
rect 144920 352446 144972 352452
rect 144274 346352 144330 346361
rect 144274 346287 144330 346296
rect 144288 345710 144316 346287
rect 144276 345704 144328 345710
rect 144276 345646 144328 345652
rect 144828 318776 144880 318782
rect 144828 318718 144880 318724
rect 144840 318102 144868 318718
rect 144828 318096 144880 318102
rect 144828 318038 144880 318044
rect 144184 314084 144236 314090
rect 144184 314026 144236 314032
rect 143816 301572 143868 301578
rect 143816 301514 143868 301520
rect 143724 286884 143776 286890
rect 143724 286826 143776 286832
rect 143736 286346 143764 286826
rect 143724 286340 143776 286346
rect 143724 286282 143776 286288
rect 142896 277432 142948 277438
rect 142896 277374 142948 277380
rect 142908 237318 142936 277374
rect 142988 253972 143040 253978
rect 142988 253914 143040 253920
rect 142896 237312 142948 237318
rect 142896 237254 142948 237260
rect 143000 220794 143028 253914
rect 142988 220788 143040 220794
rect 142988 220730 143040 220736
rect 144196 198150 144224 314026
rect 144276 296948 144328 296954
rect 144276 296890 144328 296896
rect 144288 202162 144316 296890
rect 144368 274780 144420 274786
rect 144368 274722 144420 274728
rect 144380 231742 144408 274722
rect 144460 266484 144512 266490
rect 144460 266426 144512 266432
rect 144472 240786 144500 266426
rect 144460 240780 144512 240786
rect 144460 240722 144512 240728
rect 144932 238542 144960 352446
rect 145024 285598 145052 364958
rect 145564 360324 145616 360330
rect 145564 360266 145616 360272
rect 145576 352510 145604 360266
rect 146208 357400 146260 357406
rect 146208 357342 146260 357348
rect 146220 356697 146248 357342
rect 146206 356688 146262 356697
rect 146206 356623 146262 356632
rect 145564 352504 145616 352510
rect 145564 352446 145616 352452
rect 145564 297424 145616 297430
rect 145564 297366 145616 297372
rect 145012 285592 145064 285598
rect 145012 285534 145064 285540
rect 145024 284986 145052 285534
rect 145012 284980 145064 284986
rect 145012 284922 145064 284928
rect 144920 238536 144972 238542
rect 144920 238478 144972 238484
rect 144368 231736 144420 231742
rect 144368 231678 144420 231684
rect 144276 202156 144328 202162
rect 144276 202098 144328 202104
rect 144184 198144 144236 198150
rect 144184 198086 144236 198092
rect 145576 195294 145604 297366
rect 145656 265056 145708 265062
rect 145656 264998 145708 265004
rect 145668 243574 145696 264998
rect 145656 243568 145708 243574
rect 145656 243510 145708 243516
rect 146312 238649 146340 366998
rect 146404 364342 146432 471990
rect 147864 469872 147916 469878
rect 147864 469814 147916 469820
rect 147772 460964 147824 460970
rect 147772 460906 147824 460912
rect 147680 451920 147732 451926
rect 147680 451862 147732 451868
rect 146944 392760 146996 392766
rect 146944 392702 146996 392708
rect 146956 364546 146984 392702
rect 147588 384328 147640 384334
rect 147588 384270 147640 384276
rect 147600 381546 147628 384270
rect 147588 381540 147640 381546
rect 147588 381482 147640 381488
rect 146944 364540 146996 364546
rect 146944 364482 146996 364488
rect 146392 364336 146444 364342
rect 146956 364334 146984 364482
rect 146956 364306 147076 364334
rect 146392 364278 146444 364284
rect 146404 363633 146432 364278
rect 146390 363624 146446 363633
rect 146390 363559 146446 363568
rect 146484 361412 146536 361418
rect 146484 361354 146536 361360
rect 146496 360369 146524 361354
rect 146482 360360 146538 360369
rect 146482 360295 146484 360304
rect 146536 360295 146538 360304
rect 146484 360266 146536 360272
rect 146392 358148 146444 358154
rect 146392 358090 146444 358096
rect 146404 357474 146432 358090
rect 146392 357468 146444 357474
rect 146392 357410 146444 357416
rect 146404 300150 146432 357410
rect 146944 308440 146996 308446
rect 146944 308382 146996 308388
rect 146392 300144 146444 300150
rect 146392 300086 146444 300092
rect 146298 238640 146354 238649
rect 146298 238575 146354 238584
rect 146312 238474 146340 238575
rect 146300 238468 146352 238474
rect 146300 238410 146352 238416
rect 145656 228404 145708 228410
rect 145656 228346 145708 228352
rect 145668 216034 145696 228346
rect 145656 216028 145708 216034
rect 145656 215970 145708 215976
rect 145564 195288 145616 195294
rect 145564 195230 145616 195236
rect 142804 193928 142856 193934
rect 142804 193870 142856 193876
rect 141424 192772 141476 192778
rect 141424 192714 141476 192720
rect 138756 189848 138808 189854
rect 138756 189790 138808 189796
rect 137376 187196 137428 187202
rect 137376 187138 137428 187144
rect 146956 187066 146984 308382
rect 147048 302938 147076 364306
rect 147692 342242 147720 451862
rect 147784 351898 147812 460906
rect 147876 361486 147904 469814
rect 149152 468512 149204 468518
rect 149152 468454 149204 468460
rect 149060 376712 149112 376718
rect 149060 376654 149112 376660
rect 148416 365764 148468 365770
rect 148416 365706 148468 365712
rect 147864 361480 147916 361486
rect 147864 361422 147916 361428
rect 148324 358080 148376 358086
rect 148324 358022 148376 358028
rect 147772 351892 147824 351898
rect 147772 351834 147824 351840
rect 147784 351121 147812 351834
rect 147770 351112 147826 351121
rect 147770 351047 147826 351056
rect 147680 342236 147732 342242
rect 147680 342178 147732 342184
rect 147692 341562 147720 342178
rect 147680 341556 147732 341562
rect 147680 341498 147732 341504
rect 147036 302932 147088 302938
rect 147036 302874 147088 302880
rect 147126 298208 147182 298217
rect 147126 298143 147182 298152
rect 147036 296812 147088 296818
rect 147036 296754 147088 296760
rect 147048 203794 147076 296754
rect 147140 231606 147168 298143
rect 147128 231600 147180 231606
rect 147128 231542 147180 231548
rect 148336 204270 148364 358022
rect 148428 320890 148456 365706
rect 148416 320884 148468 320890
rect 148416 320826 148468 320832
rect 148416 311160 148468 311166
rect 148416 311102 148468 311108
rect 147680 204264 147732 204270
rect 147680 204206 147732 204212
rect 148324 204264 148376 204270
rect 148324 204206 148376 204212
rect 147036 203788 147088 203794
rect 147036 203730 147088 203736
rect 147692 203590 147720 204206
rect 147680 203584 147732 203590
rect 147680 203526 147732 203532
rect 148428 197985 148456 311102
rect 148508 300280 148560 300286
rect 148508 300222 148560 300228
rect 148520 219434 148548 300222
rect 148598 295352 148654 295361
rect 148598 295287 148654 295296
rect 148612 237114 148640 295287
rect 149072 238678 149100 376654
rect 149164 360194 149192 468454
rect 150624 465112 150676 465118
rect 150624 465054 150676 465060
rect 150532 454708 150584 454714
rect 150532 454650 150584 454656
rect 149244 398880 149296 398886
rect 149244 398822 149296 398828
rect 149152 360188 149204 360194
rect 149152 360130 149204 360136
rect 149256 294710 149284 398822
rect 150440 395412 150492 395418
rect 150440 395354 150492 395360
rect 149704 360188 149756 360194
rect 149704 360130 149756 360136
rect 149716 359417 149744 360130
rect 149702 359408 149758 359417
rect 149702 359343 149758 359352
rect 149704 304360 149756 304366
rect 149704 304302 149756 304308
rect 149244 294704 149296 294710
rect 149244 294646 149296 294652
rect 149060 238672 149112 238678
rect 149060 238614 149112 238620
rect 148600 237108 148652 237114
rect 148600 237050 148652 237056
rect 148508 219428 148560 219434
rect 148508 219370 148560 219376
rect 149716 206514 149744 304302
rect 149796 295996 149848 296002
rect 149796 295938 149848 295944
rect 149808 237386 149836 295938
rect 150452 269074 150480 395354
rect 150544 343602 150572 454650
rect 150636 371890 150664 465054
rect 150624 371884 150676 371890
rect 150624 371826 150676 371832
rect 151832 368490 151860 489126
rect 151912 460216 151964 460222
rect 151912 460158 151964 460164
rect 151820 368484 151872 368490
rect 151820 368426 151872 368432
rect 151084 356720 151136 356726
rect 151084 356662 151136 356668
rect 150532 343596 150584 343602
rect 150532 343538 150584 343544
rect 150544 342961 150572 343538
rect 150530 342952 150586 342961
rect 150530 342887 150586 342896
rect 150532 340264 150584 340270
rect 150532 340206 150584 340212
rect 150544 337482 150572 340206
rect 150532 337476 150584 337482
rect 150532 337418 150584 337424
rect 151096 329186 151124 356662
rect 151924 354674 151952 460158
rect 152004 458856 152056 458862
rect 152004 458798 152056 458804
rect 151832 354646 151952 354674
rect 151832 349110 151860 354646
rect 151820 349104 151872 349110
rect 151820 349046 151872 349052
rect 152016 349042 152044 458798
rect 173164 405816 173216 405822
rect 173164 405758 173216 405764
rect 153844 403028 153896 403034
rect 153844 402970 153896 402976
rect 152096 392624 152148 392630
rect 152096 392566 152148 392572
rect 152004 349036 152056 349042
rect 152004 348978 152056 348984
rect 151728 337476 151780 337482
rect 151728 337418 151780 337424
rect 151084 329180 151136 329186
rect 151084 329122 151136 329128
rect 151084 316872 151136 316878
rect 151084 316814 151136 316820
rect 150440 269068 150492 269074
rect 150440 269010 150492 269016
rect 150452 267782 150480 269010
rect 150440 267776 150492 267782
rect 150440 267718 150492 267724
rect 150440 260840 150492 260846
rect 150440 260782 150492 260788
rect 150452 260166 150480 260782
rect 150440 260160 150492 260166
rect 150440 260102 150492 260108
rect 149796 237380 149848 237386
rect 149796 237322 149848 237328
rect 149704 206508 149756 206514
rect 149704 206450 149756 206456
rect 148414 197976 148470 197985
rect 148414 197911 148470 197920
rect 151096 196790 151124 316814
rect 151174 296848 151230 296857
rect 151174 296783 151230 296792
rect 151188 227633 151216 296783
rect 151360 264988 151412 264994
rect 151360 264930 151412 264936
rect 151268 245744 151320 245750
rect 151268 245686 151320 245692
rect 151174 227624 151230 227633
rect 151174 227559 151230 227568
rect 151084 196784 151136 196790
rect 151084 196726 151136 196732
rect 151280 192846 151308 245686
rect 151372 237250 151400 264930
rect 151740 260166 151768 337418
rect 152108 292534 152136 392566
rect 153108 349104 153160 349110
rect 153108 349046 153160 349052
rect 153016 349036 153068 349042
rect 153016 348978 153068 348984
rect 153028 348401 153056 348978
rect 153120 348430 153148 349046
rect 153108 348424 153160 348430
rect 153014 348392 153070 348401
rect 153108 348366 153160 348372
rect 153014 348327 153070 348336
rect 152648 326460 152700 326466
rect 152648 326402 152700 326408
rect 152464 309800 152516 309806
rect 152464 309742 152516 309748
rect 152096 292528 152148 292534
rect 152096 292470 152148 292476
rect 151728 260160 151780 260166
rect 151728 260102 151780 260108
rect 151360 237244 151412 237250
rect 151360 237186 151412 237192
rect 151268 192840 151320 192846
rect 151268 192782 151320 192788
rect 146944 187060 146996 187066
rect 146944 187002 146996 187008
rect 134524 185904 134576 185910
rect 134524 185846 134576 185852
rect 152476 184278 152504 309742
rect 152556 290012 152608 290018
rect 152556 289954 152608 289960
rect 152568 216102 152596 289954
rect 152660 278050 152688 326402
rect 152740 298376 152792 298382
rect 152740 298318 152792 298324
rect 152648 278044 152700 278050
rect 152648 277986 152700 277992
rect 152648 262268 152700 262274
rect 152648 262210 152700 262216
rect 152556 216096 152608 216102
rect 152556 216038 152608 216044
rect 152660 193866 152688 262210
rect 152752 238882 152780 298318
rect 152740 238876 152792 238882
rect 152740 238818 152792 238824
rect 153856 212022 153884 402970
rect 166264 400988 166316 400994
rect 166264 400930 166316 400936
rect 159364 398948 159416 398954
rect 159364 398890 159416 398896
rect 157984 398200 158036 398206
rect 157984 398142 158036 398148
rect 155224 385756 155276 385762
rect 155224 385698 155276 385704
rect 154580 376100 154632 376106
rect 154580 376042 154632 376048
rect 154592 375465 154620 376042
rect 154578 375456 154634 375465
rect 154578 375391 154634 375400
rect 153936 314016 153988 314022
rect 153936 313958 153988 313964
rect 153844 212016 153896 212022
rect 153844 211958 153896 211964
rect 152648 193860 152700 193866
rect 152648 193802 152700 193808
rect 153948 190126 153976 313958
rect 154028 267776 154080 267782
rect 154028 267718 154080 267724
rect 154040 224738 154068 267718
rect 154592 258058 154620 375391
rect 154580 258052 154632 258058
rect 154580 257994 154632 258000
rect 154028 224732 154080 224738
rect 154028 224674 154080 224680
rect 153936 190120 153988 190126
rect 153936 190062 153988 190068
rect 155236 188630 155264 385698
rect 155960 374672 156012 374678
rect 155960 374614 156012 374620
rect 155972 374202 156000 374614
rect 155960 374196 156012 374202
rect 155960 374138 156012 374144
rect 155316 317552 155368 317558
rect 155316 317494 155368 317500
rect 155328 235929 155356 317494
rect 155408 292528 155460 292534
rect 155408 292470 155460 292476
rect 155420 238785 155448 292470
rect 155500 252680 155552 252686
rect 155500 252622 155552 252628
rect 155512 242214 155540 252622
rect 155972 252550 156000 374138
rect 156604 311228 156656 311234
rect 156604 311170 156656 311176
rect 155960 252544 156012 252550
rect 155960 252486 156012 252492
rect 155500 242208 155552 242214
rect 155500 242150 155552 242156
rect 155500 240304 155552 240310
rect 155500 240246 155552 240252
rect 155406 238776 155462 238785
rect 155406 238711 155462 238720
rect 155314 235920 155370 235929
rect 155314 235855 155370 235864
rect 155512 199646 155540 240246
rect 155592 239012 155644 239018
rect 155592 238954 155644 238960
rect 155604 229022 155632 238954
rect 155592 229016 155644 229022
rect 155592 228958 155644 228964
rect 155500 199640 155552 199646
rect 155500 199582 155552 199588
rect 155224 188624 155276 188630
rect 155224 188566 155276 188572
rect 152464 184272 152516 184278
rect 152464 184214 152516 184220
rect 133328 183048 133380 183054
rect 133328 182990 133380 182996
rect 133234 181384 133290 181393
rect 133234 181319 133290 181328
rect 156616 180130 156644 311170
rect 156696 291236 156748 291242
rect 156696 291178 156748 291184
rect 156708 218822 156736 291178
rect 156788 249824 156840 249830
rect 156788 249766 156840 249772
rect 156800 233102 156828 249766
rect 156788 233096 156840 233102
rect 156788 233038 156840 233044
rect 156696 218816 156748 218822
rect 156696 218758 156748 218764
rect 157996 201074 158024 398142
rect 158168 358828 158220 358834
rect 158168 358770 158220 358776
rect 158076 295588 158128 295594
rect 158076 295530 158128 295536
rect 158088 220726 158116 295530
rect 158180 285054 158208 358770
rect 158168 285048 158220 285054
rect 158168 284990 158220 284996
rect 158168 266416 158220 266422
rect 158168 266358 158220 266364
rect 158180 235958 158208 266358
rect 158168 235952 158220 235958
rect 158168 235894 158220 235900
rect 158076 220720 158128 220726
rect 158076 220662 158128 220668
rect 157984 201068 158036 201074
rect 157984 201010 158036 201016
rect 159376 181626 159404 398890
rect 162124 398132 162176 398138
rect 162124 398074 162176 398080
rect 159456 388068 159508 388074
rect 159456 388010 159508 388016
rect 159468 209166 159496 388010
rect 160744 367192 160796 367198
rect 160744 367134 160796 367140
rect 159548 331968 159600 331974
rect 159548 331910 159600 331916
rect 159560 224806 159588 331910
rect 160756 330546 160784 367134
rect 160836 361752 160888 361758
rect 160836 361694 160888 361700
rect 160744 330540 160796 330546
rect 160744 330482 160796 330488
rect 160744 323672 160796 323678
rect 160744 323614 160796 323620
rect 159640 295520 159692 295526
rect 159640 295462 159692 295468
rect 159652 234394 159680 295462
rect 159640 234388 159692 234394
rect 159640 234330 159692 234336
rect 159548 224800 159600 224806
rect 159548 224742 159600 224748
rect 159456 209160 159508 209166
rect 159456 209102 159508 209108
rect 160756 183122 160784 323614
rect 160848 277370 160876 361694
rect 160836 277364 160888 277370
rect 160836 277306 160888 277312
rect 160928 276072 160980 276078
rect 160928 276014 160980 276020
rect 160836 260160 160888 260166
rect 160836 260102 160888 260108
rect 160848 184210 160876 260102
rect 160940 236774 160968 276014
rect 161020 258732 161072 258738
rect 161020 258674 161072 258680
rect 160928 236768 160980 236774
rect 160928 236710 160980 236716
rect 161032 230489 161060 258674
rect 161018 230480 161074 230489
rect 161018 230415 161074 230424
rect 160836 184204 160888 184210
rect 160836 184146 160888 184152
rect 160744 183116 160796 183122
rect 160744 183058 160796 183064
rect 159364 181620 159416 181626
rect 159364 181562 159416 181568
rect 156604 180124 156656 180130
rect 156604 180066 156656 180072
rect 134708 179648 134760 179654
rect 134708 179590 134760 179596
rect 129462 177712 129518 177721
rect 129462 177647 129518 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 133144 177064 133196 177070
rect 134720 177041 134748 179590
rect 148232 178356 148284 178362
rect 148232 178298 148284 178304
rect 133144 177006 133196 177012
rect 134706 177032 134762 177041
rect 133156 176769 133184 177006
rect 134706 176967 134762 176976
rect 136088 176860 136140 176866
rect 136088 176802 136140 176808
rect 136100 176769 136128 176802
rect 148244 176769 148272 178298
rect 159916 178084 159968 178090
rect 159916 178026 159968 178032
rect 159928 176769 159956 178026
rect 162136 177313 162164 398074
rect 162216 369980 162268 369986
rect 162216 369922 162268 369928
rect 162228 326534 162256 369922
rect 163596 364812 163648 364818
rect 163596 364754 163648 364760
rect 162216 326528 162268 326534
rect 162216 326470 162268 326476
rect 163504 313948 163556 313954
rect 163504 313890 163556 313896
rect 162216 306468 162268 306474
rect 162216 306410 162268 306416
rect 162228 209234 162256 306410
rect 162308 301572 162360 301578
rect 162308 301514 162360 301520
rect 162320 228886 162348 301514
rect 162400 300892 162452 300898
rect 162400 300834 162452 300840
rect 162412 240854 162440 300834
rect 162400 240848 162452 240854
rect 162400 240790 162452 240796
rect 162308 228880 162360 228886
rect 162308 228822 162360 228828
rect 162216 209228 162268 209234
rect 162216 209170 162268 209176
rect 162122 177304 162178 177313
rect 162122 177239 162178 177248
rect 104676 176760 104678 176769
rect 104622 176695 104678 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 110326 176760 110382 176769
rect 110326 176695 110382 176704
rect 113730 176760 113786 176769
rect 113730 176695 113786 176704
rect 127070 176760 127126 176769
rect 133142 176760 133198 176769
rect 127070 176695 127126 176704
rect 128176 176724 128228 176730
rect 133142 176695 133198 176704
rect 136086 176760 136142 176769
rect 136086 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 159914 176760 159970 176769
rect 159914 176695 159970 176704
rect 128176 176666 128228 176672
rect 128188 176497 128216 176666
rect 128174 176488 128230 176497
rect 128174 176423 128230 176432
rect 163516 176322 163544 313890
rect 163608 312594 163636 364754
rect 164884 362976 164936 362982
rect 164884 362918 164936 362924
rect 164896 323610 164924 362918
rect 165528 328500 165580 328506
rect 165528 328442 165580 328448
rect 164884 323604 164936 323610
rect 164884 323546 164936 323552
rect 164884 312656 164936 312662
rect 164884 312598 164936 312604
rect 163596 312588 163648 312594
rect 163596 312530 163648 312536
rect 163596 302320 163648 302326
rect 163596 302262 163648 302268
rect 163608 235482 163636 302262
rect 163688 287700 163740 287706
rect 163688 287642 163740 287648
rect 163596 235476 163648 235482
rect 163596 235418 163648 235424
rect 163700 222086 163728 287642
rect 164896 222873 164924 312598
rect 165436 308440 165488 308446
rect 165436 308382 165488 308388
rect 165448 307873 165476 308382
rect 165434 307864 165490 307873
rect 165434 307799 165490 307808
rect 164882 222864 164938 222873
rect 164882 222799 164938 222808
rect 163688 222080 163740 222086
rect 163688 222022 163740 222028
rect 164884 182436 164936 182442
rect 164884 182378 164936 182384
rect 163504 176316 163556 176322
rect 163504 176258 163556 176264
rect 120816 176248 120868 176254
rect 120816 176190 120868 176196
rect 102048 176112 102100 176118
rect 102048 176054 102100 176060
rect 102060 175409 102088 176054
rect 116952 175976 117004 175982
rect 116952 175918 117004 175924
rect 116964 175409 116992 175918
rect 120828 175409 120856 176190
rect 121920 176180 121972 176186
rect 121920 176122 121972 176128
rect 121932 175409 121960 176122
rect 130752 176044 130804 176050
rect 130752 175986 130804 175992
rect 130764 175409 130792 175986
rect 102046 175400 102102 175409
rect 102046 175335 102102 175344
rect 116950 175400 117006 175409
rect 116950 175335 117006 175344
rect 120814 175400 120870 175409
rect 120814 175335 120870 175344
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 130750 175400 130806 175409
rect 130750 175335 130806 175344
rect 164896 173874 164924 182378
rect 165448 180266 165476 307799
rect 165540 192506 165568 328442
rect 166276 200802 166304 400930
rect 167644 390720 167696 390726
rect 167644 390662 167696 390668
rect 166356 369912 166408 369918
rect 166356 369854 166408 369860
rect 166368 325038 166396 369854
rect 166356 325032 166408 325038
rect 166356 324974 166408 324980
rect 166540 315308 166592 315314
rect 166540 315250 166592 315256
rect 166356 305652 166408 305658
rect 166356 305594 166408 305600
rect 166264 200796 166316 200802
rect 166264 200738 166316 200744
rect 165528 192500 165580 192506
rect 165528 192442 165580 192448
rect 166368 181558 166396 305594
rect 166448 281580 166500 281586
rect 166448 281522 166500 281528
rect 166356 181552 166408 181558
rect 166356 181494 166408 181500
rect 165436 180260 165488 180266
rect 165436 180202 165488 180208
rect 165436 179648 165488 179654
rect 165436 179590 165488 179596
rect 165448 175234 165476 179590
rect 166264 179512 166316 179518
rect 166264 179454 166316 179460
rect 165528 177064 165580 177070
rect 165528 177006 165580 177012
rect 165436 175228 165488 175234
rect 165436 175170 165488 175176
rect 165540 175166 165568 177006
rect 165528 175160 165580 175166
rect 165528 175102 165580 175108
rect 164884 173868 164936 173874
rect 164884 173810 164936 173816
rect 166276 165578 166304 179454
rect 166460 175982 166488 281522
rect 166552 233034 166580 315250
rect 166540 233028 166592 233034
rect 166540 232970 166592 232976
rect 167656 210458 167684 390662
rect 171784 365968 171836 365974
rect 171784 365910 171836 365916
rect 169116 358896 169168 358902
rect 169116 358838 169168 358844
rect 167828 320884 167880 320890
rect 167828 320826 167880 320832
rect 167840 305046 167868 320826
rect 167828 305040 167880 305046
rect 167828 304982 167880 304988
rect 167736 254584 167788 254590
rect 167736 254526 167788 254532
rect 167644 210452 167696 210458
rect 167644 210394 167696 210400
rect 166540 181008 166592 181014
rect 166540 180950 166592 180956
rect 166356 175976 166408 175982
rect 166356 175918 166408 175924
rect 166448 175976 166500 175982
rect 166448 175918 166500 175924
rect 166368 167006 166396 175918
rect 166552 172514 166580 180950
rect 167552 176928 167604 176934
rect 167552 176870 167604 176876
rect 166632 176248 166684 176254
rect 166632 176190 166684 176196
rect 166540 172508 166592 172514
rect 166540 172450 166592 172456
rect 166644 168366 166672 176190
rect 167564 171134 167592 176870
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 167656 171358 167684 171527
rect 167644 171352 167696 171358
rect 167644 171294 167696 171300
rect 167564 171106 167684 171134
rect 166632 168360 166684 168366
rect 166632 168302 166684 168308
rect 166356 167000 166408 167006
rect 166356 166942 166408 166948
rect 166264 165572 166316 165578
rect 166264 165514 166316 165520
rect 167656 159390 167684 171106
rect 167644 159384 167696 159390
rect 167644 159326 167696 159332
rect 166264 153264 166316 153270
rect 166264 153206 166316 153212
rect 67362 128072 67418 128081
rect 67362 128007 67418 128016
rect 67270 122632 67326 122641
rect 67270 122567 67326 122576
rect 67284 89729 67312 122567
rect 67376 93809 67404 128007
rect 67454 125216 67510 125225
rect 67454 125151 67510 125160
rect 67362 93800 67418 93809
rect 67362 93735 67418 93744
rect 67468 91089 67496 125151
rect 67638 120864 67694 120873
rect 67638 120799 67694 120808
rect 67454 91080 67510 91089
rect 67652 91050 67680 120799
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67454 91015 67510 91024
rect 67640 91044 67692 91050
rect 67640 90986 67692 90992
rect 67270 89720 67326 89729
rect 67270 89655 67326 89664
rect 67744 85542 67772 100671
rect 164884 99408 164936 99414
rect 164884 99350 164936 99356
rect 85578 94752 85634 94761
rect 85578 94687 85634 94696
rect 112350 94752 112406 94761
rect 112350 94687 112406 94696
rect 122838 94752 122894 94761
rect 122838 94687 122894 94696
rect 124494 94752 124550 94761
rect 124494 94687 124550 94696
rect 85592 93906 85620 94687
rect 112364 94042 112392 94687
rect 112352 94036 112404 94042
rect 112352 93978 112404 93984
rect 122852 93974 122880 94687
rect 124508 94110 124536 94687
rect 129556 94512 129608 94518
rect 129556 94454 129608 94460
rect 124496 94104 124548 94110
rect 124496 94046 124548 94052
rect 122840 93968 122892 93974
rect 122840 93910 122892 93916
rect 85580 93900 85632 93906
rect 85580 93842 85632 93848
rect 123206 93528 123262 93537
rect 123206 93463 123262 93472
rect 123220 93294 123248 93463
rect 123208 93288 123260 93294
rect 100574 93256 100630 93265
rect 100574 93191 100630 93200
rect 110142 93256 110198 93265
rect 123208 93230 123260 93236
rect 110142 93191 110198 93200
rect 100588 93158 100616 93191
rect 100576 93152 100628 93158
rect 100576 93094 100628 93100
rect 88064 92472 88116 92478
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 84842 92440 84898 92449
rect 84842 92375 84898 92384
rect 86774 92440 86830 92449
rect 86774 92375 86830 92384
rect 88062 92440 88064 92449
rect 88116 92440 88118 92449
rect 88062 92375 88118 92384
rect 100114 92440 100170 92449
rect 100114 92375 100170 92384
rect 101954 92440 102010 92449
rect 101954 92375 102010 92384
rect 103426 92440 103482 92449
rect 103426 92375 103482 92384
rect 104438 92440 104494 92449
rect 104438 92375 104494 92384
rect 105726 92440 105782 92449
rect 105726 92375 105782 92384
rect 107566 92440 107622 92449
rect 107566 92375 107622 92384
rect 107934 92440 107990 92449
rect 107934 92375 107990 92384
rect 108302 92440 108358 92449
rect 108302 92375 108358 92384
rect 110050 92440 110106 92449
rect 110050 92375 110106 92384
rect 74828 91118 74856 92375
rect 84856 91186 84884 92375
rect 86788 92342 86816 92375
rect 86776 92336 86828 92342
rect 86776 92278 86828 92284
rect 88982 91760 89038 91769
rect 88982 91695 89038 91704
rect 84844 91180 84896 91186
rect 84844 91122 84896 91128
rect 74816 91112 74868 91118
rect 74816 91054 74868 91060
rect 88996 89690 89024 91695
rect 97446 91488 97502 91497
rect 97446 91423 97502 91432
rect 99194 91488 99250 91497
rect 99194 91423 99250 91432
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 90638 91216 90694 91225
rect 90638 91151 90694 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 88984 89684 89036 89690
rect 88984 89626 89036 89632
rect 90652 86970 90680 91151
rect 90640 86964 90692 86970
rect 90640 86906 90692 86912
rect 67732 85536 67784 85542
rect 67732 85478 67784 85484
rect 92400 84046 92428 91151
rect 92388 84040 92440 84046
rect 92388 83982 92440 83988
rect 93780 79898 93808 91151
rect 95068 82754 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97078 91216 97134 91225
rect 97078 91151 97134 91160
rect 95056 82748 95108 82754
rect 95056 82690 95108 82696
rect 95160 81258 95188 91151
rect 95148 81252 95200 81258
rect 95148 81194 95200 81200
rect 96540 79966 96568 91151
rect 97092 86766 97120 91151
rect 97460 88194 97488 91423
rect 99102 91216 99158 91225
rect 99102 91151 99158 91160
rect 97448 88188 97500 88194
rect 97448 88130 97500 88136
rect 97080 86760 97132 86766
rect 97080 86702 97132 86708
rect 99116 81433 99144 91151
rect 99102 81424 99158 81433
rect 99102 81359 99158 81368
rect 99208 80073 99236 91423
rect 99286 91352 99342 91361
rect 99286 91287 99342 91296
rect 99194 80064 99250 80073
rect 99194 79999 99250 80008
rect 96528 79960 96580 79966
rect 96528 79902 96580 79908
rect 93768 79892 93820 79898
rect 93768 79834 93820 79840
rect 99300 77178 99328 91287
rect 100128 85406 100156 92375
rect 101862 92304 101918 92313
rect 101862 92239 101918 92248
rect 100116 85400 100168 85406
rect 100116 85342 100168 85348
rect 101876 78577 101904 92239
rect 101968 79830 101996 92375
rect 103334 92304 103390 92313
rect 103334 92239 103390 92248
rect 102046 92168 102102 92177
rect 102046 92103 102102 92112
rect 102060 89554 102088 92103
rect 102048 89548 102100 89554
rect 102048 89490 102100 89496
rect 103348 84114 103376 92239
rect 103336 84108 103388 84114
rect 103336 84050 103388 84056
rect 103440 82822 103468 92375
rect 104452 88126 104480 92375
rect 104622 92304 104678 92313
rect 104622 92239 104678 92248
rect 104440 88120 104492 88126
rect 104440 88062 104492 88068
rect 104636 85474 104664 92239
rect 105740 88233 105768 92375
rect 106186 92304 106242 92313
rect 106186 92239 106242 92248
rect 107474 92304 107530 92313
rect 107474 92239 107530 92248
rect 105726 88224 105782 88233
rect 105726 88159 105782 88168
rect 104624 85468 104676 85474
rect 104624 85410 104676 85416
rect 103428 82816 103480 82822
rect 103428 82758 103480 82764
rect 106200 82686 106228 92239
rect 106188 82680 106240 82686
rect 106188 82622 106240 82628
rect 107488 81394 107516 92239
rect 107476 81388 107528 81394
rect 107476 81330 107528 81336
rect 101956 79824 102008 79830
rect 101956 79766 102008 79772
rect 101862 78568 101918 78577
rect 101862 78503 101918 78512
rect 107580 78441 107608 92375
rect 107948 86834 107976 92375
rect 108316 86873 108344 92375
rect 110064 90982 110092 92375
rect 110052 90976 110104 90982
rect 110052 90918 110104 90924
rect 108302 86864 108358 86873
rect 107936 86828 107988 86834
rect 108302 86799 108358 86808
rect 107936 86770 107988 86776
rect 110156 85338 110184 93191
rect 110694 92440 110750 92449
rect 110694 92375 110750 92384
rect 113822 92440 113878 92449
rect 113822 92375 113878 92384
rect 119342 92440 119398 92449
rect 119342 92375 119344 92384
rect 110708 92206 110736 92375
rect 110696 92200 110748 92206
rect 110696 92142 110748 92148
rect 111614 91760 111670 91769
rect 111614 91695 111670 91704
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 111156 91180 111208 91186
rect 110144 85332 110196 85338
rect 110144 85274 110196 85280
rect 110340 78674 110368 91151
rect 111156 91122 111208 91128
rect 111064 91112 111116 91118
rect 111064 91054 111116 91060
rect 110328 78668 110380 78674
rect 110328 78610 110380 78616
rect 107566 78432 107622 78441
rect 107566 78367 107622 78376
rect 99288 77172 99340 77178
rect 99288 77114 99340 77120
rect 86960 76628 87012 76634
rect 86960 76570 87012 76576
rect 69020 75268 69072 75274
rect 69020 75210 69072 75216
rect 67640 55956 67692 55962
rect 67640 55898 67692 55904
rect 67180 45552 67232 45558
rect 67180 45494 67232 45500
rect 64788 12436 64840 12442
rect 64788 12378 64840 12384
rect 65524 8968 65576 8974
rect 65524 8910 65576 8916
rect 65536 480 65564 8910
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 66732 480 66760 3538
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 55898
rect 69032 3534 69060 75210
rect 80060 73908 80112 73914
rect 80060 73850 80112 73856
rect 73160 64184 73212 64190
rect 73160 64126 73212 64132
rect 70400 54664 70452 54670
rect 70400 54606 70452 54612
rect 69112 51740 69164 51746
rect 69112 51682 69164 51688
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 51682
rect 70412 16574 70440 54606
rect 71780 50516 71832 50522
rect 71780 50458 71832 50464
rect 71792 16574 71820 50458
rect 73172 16574 73200 64126
rect 74540 58812 74592 58818
rect 74540 58754 74592 58760
rect 74552 16574 74580 58754
rect 78680 54732 78732 54738
rect 78680 54674 78732 54680
rect 77298 51776 77354 51785
rect 77298 51711 77354 51720
rect 75920 18760 75972 18766
rect 75920 18702 75972 18708
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 18702
rect 77312 3602 77340 51711
rect 77392 25560 77444 25566
rect 77392 25502 77444 25508
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77404 480 77432 25502
rect 78692 16574 78720 54674
rect 80072 16574 80100 73850
rect 84200 71052 84252 71058
rect 84200 70994 84252 71000
rect 82820 29708 82872 29714
rect 82820 29650 82872 29656
rect 81440 24268 81492 24274
rect 81440 24210 81492 24216
rect 81452 16574 81480 24210
rect 82832 16574 82860 29650
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3538
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 70994
rect 85580 50448 85632 50454
rect 85580 50390 85632 50396
rect 85592 6914 85620 50390
rect 85672 43444 85724 43450
rect 85672 43386 85724 43392
rect 85684 16574 85712 43386
rect 86972 16574 87000 76570
rect 111076 75818 111104 91054
rect 111168 77246 111196 91122
rect 111628 89486 111656 91695
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 111616 89480 111668 89486
rect 111616 89422 111668 89428
rect 113100 84153 113128 91151
rect 113836 90914 113864 92375
rect 119396 92375 119398 92384
rect 119894 92440 119950 92449
rect 119894 92375 119950 92384
rect 129462 92440 129518 92449
rect 129462 92375 129518 92384
rect 119344 92346 119396 92352
rect 117134 92168 117190 92177
rect 117134 92103 117190 92112
rect 115754 91352 115810 91361
rect 115754 91287 115810 91296
rect 114374 91216 114430 91225
rect 114374 91151 114430 91160
rect 115294 91216 115350 91225
rect 115294 91151 115350 91160
rect 113824 90908 113876 90914
rect 113824 90850 113876 90856
rect 113086 84144 113142 84153
rect 113086 84079 113142 84088
rect 114388 80034 114416 91151
rect 115308 87990 115336 91151
rect 115296 87984 115348 87990
rect 115296 87926 115348 87932
rect 115768 86698 115796 91287
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 115756 86692 115808 86698
rect 115756 86634 115808 86640
rect 115860 82793 115888 91151
rect 117148 85270 117176 92103
rect 118054 91624 118110 91633
rect 118054 91559 118110 91568
rect 118068 89418 118096 91559
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 118056 89412 118108 89418
rect 118056 89354 118108 89360
rect 117136 85264 117188 85270
rect 117136 85206 117188 85212
rect 115846 82784 115902 82793
rect 115846 82719 115902 82728
rect 118620 81190 118648 91151
rect 119908 90846 119936 92375
rect 129476 92274 129504 92375
rect 129568 92342 129596 94454
rect 151726 93664 151782 93673
rect 151726 93599 151782 93608
rect 151740 93362 151768 93599
rect 151728 93356 151780 93362
rect 151728 93298 151780 93304
rect 134708 93220 134760 93226
rect 134708 93162 134760 93168
rect 133142 92440 133198 92449
rect 133142 92375 133198 92384
rect 133156 92342 133184 92375
rect 129556 92336 129608 92342
rect 129556 92278 129608 92284
rect 133144 92336 133196 92342
rect 133144 92278 133196 92284
rect 129464 92268 129516 92274
rect 129464 92210 129516 92216
rect 134720 92206 134748 93162
rect 136086 92440 136142 92449
rect 136086 92375 136142 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152094 92440 152150 92449
rect 152094 92375 152150 92384
rect 134708 92200 134760 92206
rect 134708 92142 134760 92148
rect 136100 92138 136128 92375
rect 136088 92132 136140 92138
rect 136088 92074 136140 92080
rect 134890 91760 134946 91769
rect 134890 91695 134946 91704
rect 120906 91624 120962 91633
rect 120906 91559 120962 91568
rect 119896 90840 119948 90846
rect 119896 90782 119948 90788
rect 120920 89350 120948 91559
rect 122102 91352 122158 91361
rect 122102 91287 122158 91296
rect 126702 91352 126758 91361
rect 126702 91287 126758 91296
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 120908 89344 120960 89350
rect 120908 89286 120960 89292
rect 121380 81326 121408 91151
rect 122116 88330 122144 91287
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 126058 91216 126114 91225
rect 126058 91151 126114 91160
rect 122104 88324 122156 88330
rect 122104 88266 122156 88272
rect 122760 82618 122788 91151
rect 124140 88262 124168 91151
rect 124128 88256 124180 88262
rect 124128 88198 124180 88204
rect 125520 83978 125548 91151
rect 126072 86902 126100 91151
rect 126060 86896 126112 86902
rect 126060 86838 126112 86844
rect 126716 85202 126744 91287
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 131026 91216 131082 91225
rect 131026 91151 131082 91160
rect 126704 85196 126756 85202
rect 126704 85138 126756 85144
rect 125508 83972 125560 83978
rect 125508 83914 125560 83920
rect 122748 82612 122800 82618
rect 122748 82554 122800 82560
rect 126900 82550 126928 91151
rect 126888 82544 126940 82550
rect 126888 82486 126940 82492
rect 121368 81320 121420 81326
rect 121368 81262 121420 81268
rect 118608 81184 118660 81190
rect 118608 81126 118660 81132
rect 114376 80028 114428 80034
rect 114376 79970 114428 79976
rect 128280 78606 128308 91151
rect 131040 83910 131068 91151
rect 134904 89622 134932 91695
rect 151556 90778 151584 92375
rect 152108 92206 152136 92375
rect 152096 92200 152148 92206
rect 152096 92142 152148 92148
rect 151634 91216 151690 91225
rect 151634 91151 151690 91160
rect 151544 90772 151596 90778
rect 151544 90714 151596 90720
rect 134892 89616 134944 89622
rect 134892 89558 134944 89564
rect 151648 88058 151676 91151
rect 164896 89690 164924 99350
rect 166276 93362 166304 153206
rect 167644 125656 167696 125662
rect 167644 125598 167696 125604
rect 166356 110492 166408 110498
rect 166356 110434 166408 110440
rect 166264 93356 166316 93362
rect 166264 93298 166316 93304
rect 164884 89684 164936 89690
rect 164884 89626 164936 89632
rect 151636 88052 151688 88058
rect 151636 87994 151688 88000
rect 166368 85406 166396 110434
rect 166448 109064 166500 109070
rect 166448 109006 166500 109012
rect 166460 88194 166488 109006
rect 166540 97300 166592 97306
rect 166540 97242 166592 97248
rect 166552 92274 166580 97242
rect 166540 92268 166592 92274
rect 166540 92210 166592 92216
rect 166448 88188 166500 88194
rect 166448 88130 166500 88136
rect 166356 85400 166408 85406
rect 166356 85342 166408 85348
rect 131028 83904 131080 83910
rect 131028 83846 131080 83852
rect 167656 82550 167684 125598
rect 167748 101425 167776 254526
rect 167840 180198 167868 304982
rect 169024 299600 169076 299606
rect 169024 299542 169076 299548
rect 167920 298240 167972 298246
rect 167920 298182 167972 298188
rect 167932 250510 167960 298182
rect 167920 250504 167972 250510
rect 167920 250446 167972 250452
rect 169036 189990 169064 299542
rect 169128 288386 169156 358838
rect 170404 351212 170456 351218
rect 170404 351154 170456 351160
rect 169668 339516 169720 339522
rect 169668 339458 169720 339464
rect 169116 288380 169168 288386
rect 169116 288322 169168 288328
rect 169116 273352 169168 273358
rect 169116 273294 169168 273300
rect 169024 189984 169076 189990
rect 169024 189926 169076 189932
rect 169128 183190 169156 273294
rect 169208 256080 169260 256086
rect 169208 256022 169260 256028
rect 169220 237289 169248 256022
rect 169206 237280 169262 237289
rect 169206 237215 169262 237224
rect 169680 232558 169708 339458
rect 169668 232552 169720 232558
rect 169668 232494 169720 232500
rect 169116 183184 169168 183190
rect 169116 183126 169168 183132
rect 170416 182889 170444 351154
rect 170496 322244 170548 322250
rect 170496 322186 170548 322192
rect 170508 217326 170536 322186
rect 171796 319462 171824 365910
rect 172426 333296 172482 333305
rect 172426 333231 172482 333240
rect 172440 332625 172468 333231
rect 172426 332616 172482 332625
rect 172426 332551 172482 332560
rect 172336 320204 172388 320210
rect 172336 320146 172388 320152
rect 171784 319456 171836 319462
rect 171784 319398 171836 319404
rect 171784 318096 171836 318102
rect 171784 318038 171836 318044
rect 170588 300212 170640 300218
rect 170588 300154 170640 300160
rect 170600 223446 170628 300154
rect 170588 223440 170640 223446
rect 170588 223382 170640 223388
rect 170496 217320 170548 217326
rect 170496 217262 170548 217268
rect 170402 182880 170458 182889
rect 170402 182815 170458 182824
rect 170496 182368 170548 182374
rect 170496 182310 170548 182316
rect 167920 180940 167972 180946
rect 167920 180882 167972 180888
rect 167828 180192 167880 180198
rect 167828 180134 167880 180140
rect 167828 176112 167880 176118
rect 167828 176054 167880 176060
rect 167840 158710 167868 176054
rect 167932 169726 167960 180882
rect 169208 180872 169260 180878
rect 169208 180814 169260 180820
rect 169024 178084 169076 178090
rect 169024 178026 169076 178032
rect 167920 169720 167972 169726
rect 167920 169662 167972 169668
rect 167828 158704 167880 158710
rect 167828 158646 167880 158652
rect 169036 149054 169064 178026
rect 169116 176996 169168 177002
rect 169116 176938 169168 176944
rect 169128 161430 169156 176938
rect 169220 166938 169248 180814
rect 170404 178356 170456 178362
rect 170404 178298 170456 178304
rect 169208 166932 169260 166938
rect 169208 166874 169260 166880
rect 169116 161424 169168 161430
rect 169116 161366 169168 161372
rect 170416 150414 170444 178298
rect 170508 162858 170536 182310
rect 170680 179580 170732 179586
rect 170680 179522 170732 179528
rect 170588 171352 170640 171358
rect 170588 171294 170640 171300
rect 170496 162852 170548 162858
rect 170496 162794 170548 162800
rect 170600 155242 170628 171294
rect 170692 171086 170720 179522
rect 170680 171080 170732 171086
rect 170680 171022 170732 171028
rect 170588 155236 170640 155242
rect 170588 155178 170640 155184
rect 170404 150408 170456 150414
rect 170404 150350 170456 150356
rect 169024 149048 169076 149054
rect 169024 148990 169076 148996
rect 169024 144220 169076 144226
rect 169024 144162 169076 144168
rect 167920 140072 167972 140078
rect 167920 140014 167972 140020
rect 167828 121508 167880 121514
rect 167828 121450 167880 121456
rect 167734 101416 167790 101425
rect 167734 101351 167790 101360
rect 167736 100020 167788 100026
rect 167736 99962 167788 99968
rect 167748 92138 167776 99962
rect 167736 92132 167788 92138
rect 167736 92074 167788 92080
rect 167840 90846 167868 121450
rect 167932 113174 167960 140014
rect 167932 113146 168052 113174
rect 167920 111784 167972 111790
rect 167918 111752 167920 111761
rect 167972 111752 167974 111761
rect 167918 111687 167974 111696
rect 168024 110129 168052 113146
rect 168010 110120 168066 110129
rect 168010 110055 168066 110064
rect 169036 108769 169064 144162
rect 170404 140820 170456 140826
rect 170404 140762 170456 140768
rect 169116 117360 169168 117366
rect 169116 117302 169168 117308
rect 169022 108760 169078 108769
rect 169022 108695 169078 108704
rect 167920 107704 167972 107710
rect 167920 107646 167972 107652
rect 167828 90840 167880 90846
rect 167828 90782 167880 90788
rect 167644 82544 167696 82550
rect 167644 82486 167696 82492
rect 167932 81258 167960 107646
rect 169024 106344 169076 106350
rect 169024 106286 169076 106292
rect 167920 81252 167972 81258
rect 167920 81194 167972 81200
rect 169036 79898 169064 106286
rect 169128 85338 169156 117302
rect 169300 113212 169352 113218
rect 169300 113154 169352 113160
rect 169208 107772 169260 107778
rect 169208 107714 169260 107720
rect 169116 85332 169168 85338
rect 169116 85274 169168 85280
rect 169220 82754 169248 107714
rect 169312 88126 169340 113154
rect 170416 93294 170444 140762
rect 170496 138032 170548 138038
rect 170496 137974 170548 137980
rect 170404 93288 170456 93294
rect 170404 93230 170456 93236
rect 170508 89418 170536 137974
rect 170588 122868 170640 122874
rect 170588 122810 170640 122816
rect 170496 89412 170548 89418
rect 170496 89354 170548 89360
rect 170600 89350 170628 122810
rect 170680 118856 170732 118862
rect 170680 118798 170732 118804
rect 170588 89344 170640 89350
rect 170588 89286 170640 89292
rect 170404 89004 170456 89010
rect 170404 88946 170456 88952
rect 169300 88120 169352 88126
rect 169300 88062 169352 88068
rect 169208 82748 169260 82754
rect 169208 82690 169260 82696
rect 169024 79892 169076 79898
rect 169024 79834 169076 79840
rect 128268 78600 128320 78606
rect 128268 78542 128320 78548
rect 111156 77240 111208 77246
rect 111156 77182 111208 77188
rect 111064 75812 111116 75818
rect 111064 75754 111116 75760
rect 110420 73976 110472 73982
rect 110420 73918 110472 73924
rect 93860 68400 93912 68406
rect 93860 68342 93912 68348
rect 89720 39364 89772 39370
rect 89720 39306 89772 39312
rect 89732 16574 89760 39306
rect 92480 26920 92532 26926
rect 92480 26862 92532 26868
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 89732 16546 89944 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89168 16040 89220 16046
rect 89168 15982 89220 15988
rect 89180 480 89208 15982
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 9036 91612 9042
rect 91560 8978 91612 8984
rect 91572 480 91600 8978
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 26862
rect 93872 3602 93900 68342
rect 98000 62892 98052 62898
rect 98000 62834 98052 62840
rect 96620 40724 96672 40730
rect 96620 40666 96672 40672
rect 93952 37936 94004 37942
rect 93952 37878 94004 37884
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93964 480 93992 37878
rect 95240 29640 95292 29646
rect 95240 29582 95292 29588
rect 95252 16574 95280 29582
rect 96632 16574 96660 40666
rect 98012 16574 98040 62834
rect 104900 61532 104952 61538
rect 104900 61474 104952 61480
rect 102140 57384 102192 57390
rect 102140 57326 102192 57332
rect 99380 32496 99432 32502
rect 99380 32438 99432 32444
rect 99392 16574 99420 32438
rect 100760 31136 100812 31142
rect 100760 31078 100812 31084
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 94780 3596 94832 3602
rect 94780 3538 94832 3544
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3538
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 31078
rect 102152 16574 102180 57326
rect 103520 32428 103572 32434
rect 103520 32370 103572 32376
rect 103532 16574 103560 32370
rect 104912 16574 104940 61474
rect 106280 43512 106332 43518
rect 106280 43454 106332 43460
rect 106292 16574 106320 43454
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 102244 480 102272 16546
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 6248 108172 6254
rect 108120 6190 108172 6196
rect 108132 480 108160 6190
rect 109316 3664 109368 3670
rect 109316 3606 109368 3612
rect 109328 480 109356 3606
rect 110432 3398 110460 73918
rect 114560 72616 114612 72622
rect 114560 72558 114612 72564
rect 113180 40792 113232 40798
rect 113180 40734 113232 40740
rect 110512 39432 110564 39438
rect 110512 39374 110564 39380
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 39374
rect 111800 22908 111852 22914
rect 111800 22850 111852 22856
rect 111812 16574 111840 22850
rect 113192 16574 113220 40734
rect 114572 16574 114600 72558
rect 121460 65612 121512 65618
rect 121460 65554 121512 65560
rect 118700 60104 118752 60110
rect 118700 60046 118752 60052
rect 117320 55888 117372 55894
rect 117320 55830 117372 55836
rect 115940 44940 115992 44946
rect 115940 44882 115992 44888
rect 115952 16574 115980 44882
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 55830
rect 118712 3398 118740 60046
rect 120078 37904 120134 37913
rect 120078 37839 120134 37848
rect 118792 26988 118844 26994
rect 118792 26930 118844 26936
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 26930
rect 120092 16574 120120 37839
rect 121472 16574 121500 65554
rect 124220 49156 124272 49162
rect 124220 49098 124272 49104
rect 122840 47728 122892 47734
rect 122840 47670 122892 47676
rect 122852 16574 122880 47670
rect 124232 16574 124260 49098
rect 133144 39500 133196 39506
rect 133144 39442 133196 39448
rect 128360 27056 128412 27062
rect 128360 26998 128412 27004
rect 128372 16574 128400 26998
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 132960 6316 133012 6322
rect 132960 6258 133012 6264
rect 132972 480 133000 6258
rect 133156 3398 133184 39442
rect 164424 14544 164476 14550
rect 164424 14486 164476 14492
rect 133144 3392 133196 3398
rect 133144 3334 133196 3340
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136468 480 136496 3334
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14486
rect 170416 3534 170444 88946
rect 170692 87990 170720 118798
rect 171796 117978 171824 318038
rect 172348 310486 172376 320146
rect 172336 310480 172388 310486
rect 172336 310422 172388 310428
rect 171876 291848 171928 291854
rect 171876 291790 171928 291796
rect 171888 233986 171916 291790
rect 171876 233980 171928 233986
rect 171876 233922 171928 233928
rect 172440 198014 172468 332551
rect 173176 204921 173204 405758
rect 226984 400240 227036 400246
rect 226984 400182 227036 400188
rect 204904 398880 204956 398886
rect 204904 398822 204956 398828
rect 178684 387932 178736 387938
rect 178684 387874 178736 387880
rect 174544 378208 174596 378214
rect 174544 378150 174596 378156
rect 174556 327894 174584 378150
rect 177396 372768 177448 372774
rect 177396 372710 177448 372716
rect 176016 364744 176068 364750
rect 176016 364686 176068 364692
rect 175924 336796 175976 336802
rect 175924 336738 175976 336744
rect 175188 331900 175240 331906
rect 175188 331842 175240 331848
rect 175200 331294 175228 331842
rect 175188 331288 175240 331294
rect 175188 331230 175240 331236
rect 174544 327888 174596 327894
rect 174544 327830 174596 327836
rect 173348 310480 173400 310486
rect 173348 310422 173400 310428
rect 173256 289944 173308 289950
rect 173256 289886 173308 289892
rect 173162 204912 173218 204921
rect 173162 204847 173218 204856
rect 172428 198008 172480 198014
rect 172428 197950 172480 197956
rect 173268 184346 173296 289886
rect 173360 211818 173388 310422
rect 174636 296744 174688 296750
rect 174636 296686 174688 296692
rect 174544 270564 174596 270570
rect 174544 270506 174596 270512
rect 173348 211812 173400 211818
rect 173348 211754 173400 211760
rect 173256 184340 173308 184346
rect 173256 184282 173308 184288
rect 173164 183660 173216 183666
rect 173164 183602 173216 183608
rect 171968 182300 172020 182306
rect 171968 182242 172020 182248
rect 171876 179444 171928 179450
rect 171876 179386 171928 179392
rect 171888 155922 171916 179386
rect 171980 164218 172008 182242
rect 171968 164212 172020 164218
rect 171968 164154 172020 164160
rect 173176 161362 173204 183602
rect 174556 177546 174584 270506
rect 174648 235890 174676 296686
rect 175096 274780 175148 274786
rect 175096 274722 175148 274728
rect 175108 263634 175136 274722
rect 175096 263628 175148 263634
rect 175096 263570 175148 263576
rect 174636 235884 174688 235890
rect 174636 235826 174688 235832
rect 175096 235340 175148 235346
rect 175096 235282 175148 235288
rect 175108 235142 175136 235282
rect 175096 235136 175148 235142
rect 175096 235078 175148 235084
rect 175108 192642 175136 235078
rect 175200 221474 175228 331230
rect 175188 221468 175240 221474
rect 175188 221410 175240 221416
rect 175096 192636 175148 192642
rect 175096 192578 175148 192584
rect 174544 177540 174596 177546
rect 174544 177482 174596 177488
rect 174636 176792 174688 176798
rect 174636 176734 174688 176740
rect 173256 176180 173308 176186
rect 173256 176122 173308 176128
rect 173268 168298 173296 176122
rect 174648 169046 174676 176734
rect 174636 169040 174688 169046
rect 174636 168982 174688 168988
rect 173256 168292 173308 168298
rect 173256 168234 173308 168240
rect 173164 161356 173216 161362
rect 173164 161298 173216 161304
rect 171876 155916 171928 155922
rect 171876 155858 171928 155864
rect 174544 153332 174596 153338
rect 174544 153274 174596 153280
rect 171876 144968 171928 144974
rect 171876 144910 171928 144916
rect 171784 117972 171836 117978
rect 171784 117914 171836 117920
rect 171784 98660 171836 98666
rect 171784 98602 171836 98608
rect 171796 92478 171824 98602
rect 171784 92472 171836 92478
rect 171784 92414 171836 92420
rect 170680 87984 170732 87990
rect 170680 87926 170732 87932
rect 171888 83910 171916 144910
rect 171968 131164 172020 131170
rect 171968 131106 172020 131112
rect 171980 85474 172008 131106
rect 173256 129804 173308 129810
rect 173256 129746 173308 129752
rect 173164 127016 173216 127022
rect 173164 126958 173216 126964
rect 172060 118788 172112 118794
rect 172060 118730 172112 118736
rect 172072 94042 172100 118730
rect 172060 94036 172112 94042
rect 172060 93978 172112 93984
rect 173176 86766 173204 126958
rect 173164 86760 173216 86766
rect 173164 86702 173216 86708
rect 171968 85468 172020 85474
rect 171968 85410 172020 85416
rect 171876 83904 171928 83910
rect 171876 83846 171928 83852
rect 173268 79830 173296 129746
rect 173440 117428 173492 117434
rect 173440 117370 173492 117376
rect 173348 110560 173400 110566
rect 173348 110502 173400 110508
rect 173256 79824 173308 79830
rect 173256 79766 173308 79772
rect 173164 79348 173216 79354
rect 173164 79290 173216 79296
rect 173176 3670 173204 79290
rect 173360 77178 173388 110502
rect 173452 89486 173480 117370
rect 174556 90778 174584 153274
rect 174636 140888 174688 140894
rect 174636 140830 174688 140836
rect 174648 94110 174676 140830
rect 174728 120148 174780 120154
rect 174728 120090 174780 120096
rect 174636 94104 174688 94110
rect 174636 94046 174688 94052
rect 174544 90772 174596 90778
rect 174544 90714 174596 90720
rect 173440 89480 173492 89486
rect 173440 89422 173492 89428
rect 174740 85270 174768 120090
rect 174820 111852 174872 111858
rect 174820 111794 174872 111800
rect 174832 89554 174860 111794
rect 174820 89548 174872 89554
rect 174820 89490 174872 89496
rect 174728 85264 174780 85270
rect 174728 85206 174780 85212
rect 173348 77172 173400 77178
rect 173348 77114 173400 77120
rect 175936 30326 175964 336738
rect 176028 326398 176056 364686
rect 177304 351212 177356 351218
rect 177304 351154 177356 351160
rect 176016 326392 176068 326398
rect 176016 326334 176068 326340
rect 176568 300144 176620 300150
rect 176568 300086 176620 300092
rect 176580 299674 176608 300086
rect 176568 299668 176620 299674
rect 176568 299610 176620 299616
rect 176016 269340 176068 269346
rect 176016 269282 176068 269288
rect 176028 235142 176056 269282
rect 176108 243024 176160 243030
rect 176108 242966 176160 242972
rect 176120 238513 176148 242966
rect 176106 238504 176162 238513
rect 176106 238439 176162 238448
rect 176016 235136 176068 235142
rect 176016 235078 176068 235084
rect 176580 214606 176608 299610
rect 176568 214600 176620 214606
rect 176568 214542 176620 214548
rect 176016 146328 176068 146334
rect 176016 146270 176068 146276
rect 176028 92342 176056 146270
rect 176108 125724 176160 125730
rect 176108 125666 176160 125672
rect 176016 92336 176068 92342
rect 176016 92278 176068 92284
rect 176120 83978 176148 125666
rect 176108 83972 176160 83978
rect 176108 83914 176160 83920
rect 175924 30320 175976 30326
rect 175924 30262 175976 30268
rect 173164 3664 173216 3670
rect 173164 3606 173216 3612
rect 170404 3528 170456 3534
rect 170404 3470 170456 3476
rect 177316 3058 177344 351154
rect 177408 336025 177436 372710
rect 177488 370048 177540 370054
rect 177488 369990 177540 369996
rect 177394 336016 177450 336025
rect 177394 335951 177450 335960
rect 177396 329112 177448 329118
rect 177396 329054 177448 329060
rect 177408 4146 177436 329054
rect 177500 319530 177528 369990
rect 177488 319524 177540 319530
rect 177488 319466 177540 319472
rect 177488 316804 177540 316810
rect 177488 316746 177540 316752
rect 177500 220318 177528 316746
rect 177948 273284 178000 273290
rect 177948 273226 178000 273232
rect 177488 220312 177540 220318
rect 177488 220254 177540 220260
rect 177960 199510 177988 273226
rect 177948 199504 178000 199510
rect 177948 199446 178000 199452
rect 177488 133952 177540 133958
rect 177488 133894 177540 133900
rect 177500 78674 177528 133894
rect 177580 114572 177632 114578
rect 177580 114514 177632 114520
rect 177592 82686 177620 114514
rect 178696 86290 178724 387874
rect 184204 387864 184256 387870
rect 184204 387806 184256 387812
rect 181444 381608 181496 381614
rect 181444 381550 181496 381556
rect 180248 367328 180300 367334
rect 180248 367270 180300 367276
rect 178868 363112 178920 363118
rect 178868 363054 178920 363060
rect 178776 341556 178828 341562
rect 178776 341498 178828 341504
rect 178788 280838 178816 341498
rect 178880 327758 178908 363054
rect 180156 362228 180208 362234
rect 180156 362170 180208 362176
rect 180064 347064 180116 347070
rect 180064 347006 180116 347012
rect 178868 327752 178920 327758
rect 178868 327694 178920 327700
rect 178868 309256 178920 309262
rect 178868 309198 178920 309204
rect 178776 280832 178828 280838
rect 178776 280774 178828 280780
rect 178776 263628 178828 263634
rect 178776 263570 178828 263576
rect 178788 182850 178816 263570
rect 178880 233170 178908 309198
rect 179418 267064 179474 267073
rect 179418 266999 179474 267008
rect 179432 266422 179460 266999
rect 179420 266416 179472 266422
rect 179420 266358 179472 266364
rect 178960 247104 179012 247110
rect 178960 247046 179012 247052
rect 178868 233164 178920 233170
rect 178868 233106 178920 233112
rect 178880 195430 178908 233106
rect 178972 227662 179000 247046
rect 178960 227656 179012 227662
rect 178960 227598 179012 227604
rect 178868 195424 178920 195430
rect 178868 195366 178920 195372
rect 178776 182844 178828 182850
rect 178776 182786 178828 182792
rect 178776 178288 178828 178294
rect 178776 178230 178828 178236
rect 178788 162790 178816 178230
rect 178776 162784 178828 162790
rect 178776 162726 178828 162732
rect 178776 135312 178828 135318
rect 178776 135254 178828 135260
rect 178788 90914 178816 135254
rect 178868 120216 178920 120222
rect 178868 120158 178920 120164
rect 178776 90908 178828 90914
rect 178776 90850 178828 90856
rect 178880 86698 178908 120158
rect 178960 109132 179012 109138
rect 178960 109074 179012 109080
rect 178868 86692 178920 86698
rect 178868 86634 178920 86640
rect 178684 86284 178736 86290
rect 178684 86226 178736 86232
rect 178682 84824 178738 84833
rect 178682 84759 178738 84768
rect 177580 82680 177632 82686
rect 177580 82622 177632 82628
rect 177488 78668 177540 78674
rect 177488 78610 177540 78616
rect 177396 4140 177448 4146
rect 177396 4082 177448 4088
rect 178696 3466 178724 84759
rect 178972 79966 179000 109074
rect 178960 79960 179012 79966
rect 178960 79902 179012 79908
rect 180076 4826 180104 347006
rect 180168 66978 180196 362170
rect 180260 319598 180288 367270
rect 180248 319592 180300 319598
rect 180248 319534 180300 319540
rect 180248 294024 180300 294030
rect 180248 293966 180300 293972
rect 180260 178838 180288 293966
rect 180340 281580 180392 281586
rect 180340 281522 180392 281528
rect 180352 269346 180380 281522
rect 180340 269340 180392 269346
rect 180340 269282 180392 269288
rect 180708 266416 180760 266422
rect 180708 266358 180760 266364
rect 180720 206310 180748 266358
rect 180708 206304 180760 206310
rect 180708 206246 180760 206252
rect 180248 178832 180300 178838
rect 180248 178774 180300 178780
rect 180248 131232 180300 131238
rect 180248 131174 180300 131180
rect 180260 88233 180288 131174
rect 180246 88224 180302 88233
rect 180246 88159 180302 88168
rect 180156 66972 180208 66978
rect 180156 66914 180208 66920
rect 181456 11762 181484 381550
rect 182824 354748 182876 354754
rect 182824 354690 182876 354696
rect 181536 312588 181588 312594
rect 181536 312530 181588 312536
rect 181548 227526 181576 312530
rect 181628 289944 181680 289950
rect 181628 289886 181680 289892
rect 181640 288425 181668 289886
rect 181626 288416 181682 288425
rect 181626 288351 181682 288360
rect 181536 227520 181588 227526
rect 181536 227462 181588 227468
rect 181548 189786 181576 227462
rect 181640 220114 181668 288351
rect 181812 256012 181864 256018
rect 181812 255954 181864 255960
rect 181824 255338 181852 255954
rect 181812 255332 181864 255338
rect 181812 255274 181864 255280
rect 182088 255332 182140 255338
rect 182088 255274 182140 255280
rect 182100 231130 182128 255274
rect 182088 231124 182140 231130
rect 182088 231066 182140 231072
rect 181628 220108 181680 220114
rect 181628 220050 181680 220056
rect 181536 189780 181588 189786
rect 181536 189722 181588 189728
rect 181536 142180 181588 142186
rect 181536 142122 181588 142128
rect 181548 85202 181576 142122
rect 181628 106412 181680 106418
rect 181628 106354 181680 106360
rect 181536 85196 181588 85202
rect 181536 85138 181588 85144
rect 181640 84046 181668 106354
rect 181628 84040 181680 84046
rect 181628 83982 181680 83988
rect 182836 38622 182864 354690
rect 183008 346452 183060 346458
rect 183008 346394 183060 346400
rect 182916 298172 182968 298178
rect 182916 298114 182968 298120
rect 182928 213382 182956 298114
rect 183020 296002 183048 346394
rect 183008 295996 183060 296002
rect 183008 295938 183060 295944
rect 183468 278044 183520 278050
rect 183468 277986 183520 277992
rect 183480 277438 183508 277986
rect 183468 277432 183520 277438
rect 183468 277374 183520 277380
rect 183376 264240 183428 264246
rect 183376 264182 183428 264188
rect 183388 263634 183416 264182
rect 183376 263628 183428 263634
rect 183376 263570 183428 263576
rect 183388 237046 183416 263570
rect 183376 237040 183428 237046
rect 183376 236982 183428 236988
rect 183480 222902 183508 277374
rect 183468 222896 183520 222902
rect 183468 222838 183520 222844
rect 182916 213376 182968 213382
rect 182916 213318 182968 213324
rect 182916 121576 182968 121582
rect 182916 121518 182968 121524
rect 182928 81190 182956 121518
rect 182916 81184 182968 81190
rect 182916 81126 182968 81132
rect 182824 38616 182876 38622
rect 182824 38558 182876 38564
rect 184216 33114 184244 387806
rect 192484 380180 192536 380186
rect 192484 380122 192536 380128
rect 185584 373312 185636 373318
rect 185584 373254 185636 373260
rect 184848 314696 184900 314702
rect 184848 314638 184900 314644
rect 184756 301504 184808 301510
rect 184756 301446 184808 301452
rect 184768 300218 184796 301446
rect 184756 300212 184808 300218
rect 184756 300154 184808 300160
rect 184296 251252 184348 251258
rect 184296 251194 184348 251200
rect 184308 238066 184336 251194
rect 184296 238060 184348 238066
rect 184296 238002 184348 238008
rect 184768 215966 184796 300154
rect 184756 215960 184808 215966
rect 184756 215902 184808 215908
rect 184860 182918 184888 314638
rect 184848 182912 184900 182918
rect 184848 182854 184900 182860
rect 184296 122936 184348 122942
rect 184296 122878 184348 122884
rect 184308 82618 184336 122878
rect 184296 82612 184348 82618
rect 184296 82554 184348 82560
rect 185596 39506 185624 373254
rect 189724 365900 189776 365906
rect 189724 365842 189776 365848
rect 188436 364676 188488 364682
rect 188436 364618 188488 364624
rect 187056 363248 187108 363254
rect 187056 363190 187108 363196
rect 186964 344344 187016 344350
rect 186964 344286 187016 344292
rect 185676 327140 185728 327146
rect 185676 327082 185728 327088
rect 185688 309194 185716 327082
rect 186320 311160 186372 311166
rect 186320 311102 186372 311108
rect 186332 310554 186360 311102
rect 186320 310548 186372 310554
rect 186320 310490 186372 310496
rect 185676 309188 185728 309194
rect 185676 309130 185728 309136
rect 185688 225758 185716 309130
rect 186228 302932 186280 302938
rect 186228 302874 186280 302880
rect 186240 302297 186268 302874
rect 186226 302288 186282 302297
rect 186226 302223 186282 302232
rect 186136 280832 186188 280838
rect 186136 280774 186188 280780
rect 186148 280226 186176 280774
rect 186136 280220 186188 280226
rect 186136 280162 186188 280168
rect 185676 225752 185728 225758
rect 185676 225694 185728 225700
rect 186148 214878 186176 280162
rect 186136 214872 186188 214878
rect 186136 214814 186188 214820
rect 185676 124228 185728 124234
rect 185676 124170 185728 124176
rect 185688 93974 185716 124170
rect 186240 96626 186268 302223
rect 186320 261520 186372 261526
rect 186320 261462 186372 261468
rect 186332 260914 186360 261462
rect 186320 260908 186372 260914
rect 186320 260850 186372 260856
rect 186228 96620 186280 96626
rect 186228 96562 186280 96568
rect 185676 93968 185728 93974
rect 185676 93910 185728 93916
rect 186976 71126 187004 344286
rect 187068 281518 187096 363190
rect 188344 348424 188396 348430
rect 188344 348366 188396 348372
rect 187608 311160 187660 311166
rect 187608 311102 187660 311108
rect 187056 281512 187108 281518
rect 187056 281454 187108 281460
rect 187056 274712 187108 274718
rect 187056 274654 187108 274660
rect 187068 235414 187096 274654
rect 187516 260908 187568 260914
rect 187516 260850 187568 260856
rect 187056 235408 187108 235414
rect 187056 235350 187108 235356
rect 187528 213246 187556 260850
rect 187620 227118 187648 311102
rect 187700 289128 187752 289134
rect 187700 289070 187752 289076
rect 187712 288454 187740 289070
rect 187700 288448 187752 288454
rect 187700 288390 187752 288396
rect 187700 230308 187752 230314
rect 187700 230250 187752 230256
rect 187712 229770 187740 230250
rect 187700 229764 187752 229770
rect 187700 229706 187752 229712
rect 187608 227112 187660 227118
rect 187608 227054 187660 227060
rect 187516 213240 187568 213246
rect 187516 213182 187568 213188
rect 187148 143608 187200 143614
rect 187148 143550 187200 143556
rect 187056 80708 187108 80714
rect 187056 80650 187108 80656
rect 186964 71120 187016 71126
rect 186964 71062 187016 71068
rect 185584 39500 185636 39506
rect 185584 39442 185636 39448
rect 184204 33108 184256 33114
rect 184204 33050 184256 33056
rect 181444 11756 181496 11762
rect 181444 11698 181496 11704
rect 180064 4820 180116 4826
rect 180064 4762 180116 4768
rect 187068 3602 187096 80650
rect 187160 78606 187188 143550
rect 187148 78600 187200 78606
rect 187148 78542 187200 78548
rect 188356 27606 188384 348366
rect 188448 334626 188476 364618
rect 188436 334620 188488 334626
rect 188436 334562 188488 334568
rect 189736 333946 189764 365842
rect 191104 356244 191156 356250
rect 191104 356186 191156 356192
rect 191116 339386 191144 356186
rect 191104 339380 191156 339386
rect 191104 339322 191156 339328
rect 189724 333940 189776 333946
rect 189724 333882 189776 333888
rect 189080 333260 189132 333266
rect 189080 333202 189132 333208
rect 190368 333260 190420 333266
rect 190368 333202 190420 333208
rect 189092 332654 189120 333202
rect 189080 332648 189132 332654
rect 189080 332590 189132 332596
rect 188988 310616 189040 310622
rect 188988 310558 189040 310564
rect 188896 288448 188948 288454
rect 188896 288390 188948 288396
rect 188804 258732 188856 258738
rect 188804 258674 188856 258680
rect 188816 229770 188844 258674
rect 188804 229764 188856 229770
rect 188804 229706 188856 229712
rect 188908 204950 188936 288390
rect 188896 204944 188948 204950
rect 188896 204886 188948 204892
rect 188436 103556 188488 103562
rect 188436 103498 188488 103504
rect 188448 93770 188476 103498
rect 189000 95169 189028 310558
rect 189724 298308 189776 298314
rect 189724 298250 189776 298256
rect 189736 196858 189764 298250
rect 190276 282940 190328 282946
rect 190276 282882 190328 282888
rect 189816 244928 189868 244934
rect 189816 244870 189868 244876
rect 189828 232626 189856 244870
rect 189816 232620 189868 232626
rect 189816 232562 189868 232568
rect 190288 228410 190316 282882
rect 190380 237969 190408 333202
rect 191104 316736 191156 316742
rect 191104 316678 191156 316684
rect 190366 237960 190422 237969
rect 190366 237895 190422 237904
rect 190276 228404 190328 228410
rect 190276 228346 190328 228352
rect 189724 196852 189776 196858
rect 189724 196794 189776 196800
rect 189724 151836 189776 151842
rect 189724 151778 189776 151784
rect 188986 95160 189042 95169
rect 188986 95095 189042 95104
rect 188436 93764 188488 93770
rect 188436 93706 188488 93712
rect 189736 92206 189764 151778
rect 189724 92200 189776 92206
rect 189724 92142 189776 92148
rect 188344 27600 188396 27606
rect 188344 27542 188396 27548
rect 191116 4078 191144 316678
rect 191196 285728 191248 285734
rect 191196 285670 191248 285676
rect 191208 240242 191236 285670
rect 191748 252612 191800 252618
rect 191748 252554 191800 252560
rect 191656 242956 191708 242962
rect 191656 242898 191708 242904
rect 191196 240236 191248 240242
rect 191196 240178 191248 240184
rect 191208 185706 191236 240178
rect 191668 239426 191696 242898
rect 191656 239420 191708 239426
rect 191656 239362 191708 239368
rect 191760 200938 191788 252554
rect 191748 200932 191800 200938
rect 191748 200874 191800 200880
rect 191196 185700 191248 185706
rect 191196 185642 191248 185648
rect 192496 83502 192524 380122
rect 197268 376780 197320 376786
rect 197268 376722 197320 376728
rect 193956 372836 194008 372842
rect 193956 372778 194008 372784
rect 193496 361820 193548 361826
rect 193496 361762 193548 361768
rect 193508 358086 193536 361762
rect 193864 358964 193916 358970
rect 193864 358906 193916 358912
rect 193496 358080 193548 358086
rect 193496 358022 193548 358028
rect 193128 317484 193180 317490
rect 193128 317426 193180 317432
rect 193036 302252 193088 302258
rect 193036 302194 193088 302200
rect 192576 278792 192628 278798
rect 192576 278734 192628 278740
rect 192588 190058 192616 278734
rect 192852 251660 192904 251666
rect 192852 251602 192904 251608
rect 192864 251297 192892 251602
rect 192850 251288 192906 251297
rect 192850 251223 192906 251232
rect 193048 231198 193076 302194
rect 193140 233889 193168 317426
rect 193876 285666 193904 358906
rect 193968 356726 193996 372778
rect 197280 368490 197308 376722
rect 204916 374066 204944 398822
rect 222844 389292 222896 389298
rect 222844 389234 222896 389240
rect 204904 374060 204956 374066
rect 204904 374002 204956 374008
rect 209780 374060 209832 374066
rect 209780 374002 209832 374008
rect 200764 371408 200816 371414
rect 200764 371350 200816 371356
rect 197268 368484 197320 368490
rect 197268 368426 197320 368432
rect 198004 368484 198056 368490
rect 198004 368426 198056 368432
rect 195244 363316 195296 363322
rect 195244 363258 195296 363264
rect 193956 356720 194008 356726
rect 193956 356662 194008 356668
rect 194508 297288 194560 297294
rect 194508 297230 194560 297236
rect 193864 285660 193916 285666
rect 193864 285602 193916 285608
rect 194324 268252 194376 268258
rect 194324 268194 194376 268200
rect 194232 243840 194284 243846
rect 194232 243782 194284 243788
rect 193864 242208 193916 242214
rect 193864 242150 193916 242156
rect 193126 233880 193182 233889
rect 193126 233815 193182 233824
rect 193036 231192 193088 231198
rect 193036 231134 193088 231140
rect 193876 226166 193904 242150
rect 194244 235550 194272 243782
rect 194336 243710 194364 268194
rect 194416 259480 194468 259486
rect 194416 259422 194468 259428
rect 194428 258738 194456 259422
rect 194416 258732 194468 258738
rect 194416 258674 194468 258680
rect 194416 250504 194468 250510
rect 194416 250446 194468 250452
rect 194428 249966 194456 250446
rect 194416 249960 194468 249966
rect 194416 249902 194468 249908
rect 194324 243704 194376 243710
rect 194324 243646 194376 243652
rect 194232 235544 194284 235550
rect 194232 235486 194284 235492
rect 193864 226160 193916 226166
rect 193864 226102 193916 226108
rect 194428 207670 194456 249902
rect 194520 240106 194548 297230
rect 195256 289814 195284 363258
rect 195336 363180 195388 363186
rect 195336 363122 195388 363128
rect 195348 294545 195376 363122
rect 196624 363044 196676 363050
rect 196624 362986 196676 362992
rect 195428 335640 195480 335646
rect 195428 335582 195480 335588
rect 195440 312594 195468 335582
rect 195428 312588 195480 312594
rect 195428 312530 195480 312536
rect 195704 295384 195756 295390
rect 195704 295326 195756 295332
rect 195334 294536 195390 294545
rect 195334 294471 195390 294480
rect 195336 292664 195388 292670
rect 195336 292606 195388 292612
rect 195244 289808 195296 289814
rect 195244 289750 195296 289756
rect 195244 273964 195296 273970
rect 195244 273906 195296 273912
rect 194508 240100 194560 240106
rect 194508 240042 194560 240048
rect 195060 239488 195112 239494
rect 195060 239430 195112 239436
rect 195072 236609 195100 239430
rect 195058 236600 195114 236609
rect 195058 236535 195114 236544
rect 195150 235240 195206 235249
rect 195150 235175 195206 235184
rect 195164 234530 195192 235175
rect 195152 234524 195204 234530
rect 195152 234466 195204 234472
rect 195256 221610 195284 273906
rect 195348 249014 195376 292606
rect 195336 249008 195388 249014
rect 195336 248950 195388 248956
rect 195348 245070 195376 248950
rect 195336 245064 195388 245070
rect 195336 245006 195388 245012
rect 195336 243568 195388 243574
rect 195336 243510 195388 243516
rect 195348 238542 195376 243510
rect 195716 240281 195744 295326
rect 196636 294642 196664 362986
rect 196716 362228 196768 362234
rect 196716 362170 196768 362176
rect 196728 307086 196756 362170
rect 196808 361684 196860 361690
rect 196808 361626 196860 361632
rect 196820 324970 196848 361626
rect 196900 360256 196952 360262
rect 196900 360198 196952 360204
rect 196912 337414 196940 360198
rect 197358 356280 197414 356289
rect 197358 356215 197360 356224
rect 197412 356215 197414 356224
rect 197360 356186 197412 356192
rect 198016 353705 198044 368426
rect 199384 366036 199436 366042
rect 199384 365978 199436 365984
rect 198648 364404 198700 364410
rect 198648 364346 198700 364352
rect 198188 360936 198240 360942
rect 198188 360878 198240 360884
rect 198096 357468 198148 357474
rect 198096 357410 198148 357416
rect 198002 353696 198058 353705
rect 198002 353631 198058 353640
rect 198108 349625 198136 357410
rect 198200 354006 198228 360878
rect 198660 356289 198688 364346
rect 198740 356992 198792 356998
rect 198740 356934 198792 356940
rect 198646 356280 198702 356289
rect 198646 356215 198702 356224
rect 198188 354000 198240 354006
rect 198188 353942 198240 353948
rect 198186 351520 198242 351529
rect 198186 351455 198242 351464
rect 198094 349616 198150 349625
rect 198094 349551 198150 349560
rect 197358 347440 197414 347449
rect 197358 347375 197414 347384
rect 197372 346458 197400 347375
rect 197360 346452 197412 346458
rect 197360 346394 197412 346400
rect 198094 344720 198150 344729
rect 198094 344655 198150 344664
rect 198002 342680 198058 342689
rect 198002 342615 198058 342624
rect 197358 340640 197414 340649
rect 197358 340575 197414 340584
rect 197372 339522 197400 340575
rect 197360 339516 197412 339522
rect 197360 339458 197412 339464
rect 197358 337920 197414 337929
rect 197358 337855 197414 337864
rect 197372 337482 197400 337855
rect 197360 337476 197412 337482
rect 197360 337418 197412 337424
rect 196900 337408 196952 337414
rect 196900 337350 196952 337356
rect 197726 335880 197782 335889
rect 197726 335815 197782 335824
rect 197740 335646 197768 335815
rect 197728 335640 197780 335646
rect 197728 335582 197780 335588
rect 197358 331800 197414 331809
rect 197358 331735 197414 331744
rect 197372 331294 197400 331735
rect 197360 331288 197412 331294
rect 197360 331230 197412 331236
rect 197358 329080 197414 329089
rect 197358 329015 197414 329024
rect 197372 328506 197400 329015
rect 197360 328500 197412 328506
rect 197360 328442 197412 328448
rect 197358 327176 197414 327185
rect 197358 327111 197360 327120
rect 197412 327111 197414 327120
rect 197360 327082 197412 327088
rect 196808 324964 196860 324970
rect 196808 324906 196860 324912
rect 197360 322924 197412 322930
rect 197360 322866 197412 322872
rect 197372 322425 197400 322866
rect 197358 322416 197414 322425
rect 197358 322351 197414 322360
rect 197358 320240 197414 320249
rect 197358 320175 197360 320184
rect 197412 320175 197414 320184
rect 197360 320146 197412 320152
rect 197358 318200 197414 318209
rect 197358 318135 197414 318144
rect 197372 317490 197400 318135
rect 197360 317484 197412 317490
rect 197360 317426 197412 317432
rect 197358 315480 197414 315489
rect 197358 315415 197414 315424
rect 197372 314702 197400 315415
rect 197360 314696 197412 314702
rect 197360 314638 197412 314644
rect 197358 313440 197414 313449
rect 197358 313375 197414 313384
rect 197372 313342 197400 313375
rect 197360 313336 197412 313342
rect 197360 313278 197412 313284
rect 197358 311400 197414 311409
rect 197358 311335 197414 311344
rect 197372 310622 197400 311335
rect 197360 310616 197412 310622
rect 197360 310558 197412 310564
rect 197358 309360 197414 309369
rect 197358 309295 197414 309304
rect 197372 309262 197400 309295
rect 197360 309256 197412 309262
rect 197360 309198 197412 309204
rect 196716 307080 196768 307086
rect 196716 307022 196768 307028
rect 197266 306640 197322 306649
rect 197266 306575 197322 306584
rect 197280 300150 197308 306575
rect 197452 306332 197504 306338
rect 197452 306274 197504 306280
rect 197358 302560 197414 302569
rect 197358 302495 197414 302504
rect 197372 302258 197400 302495
rect 197360 302252 197412 302258
rect 197360 302194 197412 302200
rect 197360 300212 197412 300218
rect 197360 300154 197412 300160
rect 197268 300144 197320 300150
rect 197268 300086 197320 300092
rect 197372 299985 197400 300154
rect 197358 299976 197414 299985
rect 197358 299911 197414 299920
rect 197358 297800 197414 297809
rect 197358 297735 197414 297744
rect 197372 297294 197400 297735
rect 197360 297288 197412 297294
rect 197360 297230 197412 297236
rect 197464 296714 197492 306274
rect 197726 304600 197782 304609
rect 197726 304535 197782 304544
rect 197740 303686 197768 304535
rect 197728 303680 197780 303686
rect 197728 303622 197780 303628
rect 198016 302938 198044 342615
rect 198108 311166 198136 344655
rect 198200 320890 198228 351455
rect 198752 351218 198780 356934
rect 198740 351212 198792 351218
rect 198740 351154 198792 351160
rect 198922 333840 198978 333849
rect 198922 333775 198978 333784
rect 198278 325000 198334 325009
rect 198278 324935 198334 324944
rect 198188 320884 198240 320890
rect 198188 320826 198240 320832
rect 198096 311160 198148 311166
rect 198096 311102 198148 311108
rect 198292 308446 198320 324935
rect 198646 324864 198702 324873
rect 198936 324850 198964 333775
rect 198702 324822 198964 324850
rect 198646 324799 198702 324808
rect 198830 313440 198886 313449
rect 198830 313375 198886 313384
rect 198280 308440 198332 308446
rect 198280 308382 198332 308388
rect 198648 303680 198700 303686
rect 198648 303622 198700 303628
rect 198004 302932 198056 302938
rect 198004 302874 198056 302880
rect 197372 296686 197492 296714
rect 196624 294636 196676 294642
rect 196624 294578 196676 294584
rect 196714 293720 196770 293729
rect 196714 293655 196770 293664
rect 196624 292596 196676 292602
rect 196624 292538 196676 292544
rect 195980 284980 196032 284986
rect 195980 284922 196032 284928
rect 195888 245676 195940 245682
rect 195888 245618 195940 245624
rect 195796 240848 195848 240854
rect 195796 240790 195848 240796
rect 195702 240272 195758 240281
rect 195702 240207 195758 240216
rect 195808 238754 195836 240790
rect 195900 239737 195928 245618
rect 195992 243846 196020 284922
rect 195980 243840 196032 243846
rect 195980 243782 196032 243788
rect 195980 243704 196032 243710
rect 195980 243646 196032 243652
rect 195886 239728 195942 239737
rect 195886 239663 195942 239672
rect 195992 239018 196020 243646
rect 196532 240780 196584 240786
rect 196532 240722 196584 240728
rect 195980 239012 196032 239018
rect 195980 238954 196032 238960
rect 195808 238726 195928 238754
rect 195336 238536 195388 238542
rect 195336 238478 195388 238484
rect 195900 237182 195928 238726
rect 195888 237176 195940 237182
rect 195888 237118 195940 237124
rect 195980 237108 196032 237114
rect 195980 237050 196032 237056
rect 195336 236768 195388 236774
rect 195992 236745 196020 237050
rect 195336 236710 195388 236716
rect 195978 236736 196034 236745
rect 195348 230314 195376 236710
rect 195978 236671 196034 236680
rect 195886 236056 195942 236065
rect 195886 235991 195942 236000
rect 195336 230308 195388 230314
rect 195336 230250 195388 230256
rect 195244 221604 195296 221610
rect 195244 221546 195296 221552
rect 194416 207664 194468 207670
rect 194416 207606 194468 207612
rect 195244 205148 195296 205154
rect 195244 205090 195296 205096
rect 192576 190052 192628 190058
rect 192576 189994 192628 190000
rect 193864 124296 193916 124302
rect 193864 124238 193916 124244
rect 192576 116000 192628 116006
rect 192576 115942 192628 115948
rect 192588 86834 192616 115942
rect 192668 102196 192720 102202
rect 192668 102138 192720 102144
rect 192680 93838 192708 102138
rect 192668 93832 192720 93838
rect 192668 93774 192720 93780
rect 193876 88262 193904 124238
rect 193864 88256 193916 88262
rect 193864 88198 193916 88204
rect 192576 86828 192628 86834
rect 192576 86770 192628 86776
rect 192484 83496 192536 83502
rect 192484 83438 192536 83444
rect 195256 42770 195284 205090
rect 195336 190120 195388 190126
rect 195336 190062 195388 190068
rect 195348 82142 195376 190062
rect 195900 178702 195928 235991
rect 196544 234530 196572 240722
rect 196636 238134 196664 292538
rect 196728 251666 196756 293655
rect 196808 286340 196860 286346
rect 196808 286282 196860 286288
rect 196716 251660 196768 251666
rect 196716 251602 196768 251608
rect 196716 245064 196768 245070
rect 196716 245006 196768 245012
rect 196624 238128 196676 238134
rect 196624 238070 196676 238076
rect 196624 235476 196676 235482
rect 196624 235418 196676 235424
rect 196532 234524 196584 234530
rect 196532 234466 196584 234472
rect 195980 222216 196032 222222
rect 195980 222158 196032 222164
rect 195992 222018 196020 222158
rect 195980 222012 196032 222018
rect 195980 221954 196032 221960
rect 196636 207874 196664 235418
rect 196624 207868 196676 207874
rect 196624 207810 196676 207816
rect 196624 206508 196676 206514
rect 196624 206450 196676 206456
rect 195888 178696 195940 178702
rect 195888 178638 195940 178644
rect 195336 82136 195388 82142
rect 195336 82078 195388 82084
rect 196636 78062 196664 206450
rect 196728 181490 196756 245006
rect 196820 242185 196848 286282
rect 197372 267734 197400 296686
rect 197450 295760 197506 295769
rect 197450 295695 197506 295704
rect 197464 295390 197492 295695
rect 197452 295384 197504 295390
rect 197452 295326 197504 295332
rect 197450 291000 197506 291009
rect 197450 290935 197506 290944
rect 197464 289950 197492 290935
rect 197452 289944 197504 289950
rect 197452 289886 197504 289892
rect 198004 289876 198056 289882
rect 198004 289818 198056 289824
rect 197450 288960 197506 288969
rect 197450 288895 197506 288904
rect 197464 288454 197492 288895
rect 197452 288448 197504 288454
rect 197452 288390 197504 288396
rect 197450 286920 197506 286929
rect 197450 286855 197506 286864
rect 197464 285734 197492 286855
rect 197452 285728 197504 285734
rect 197452 285670 197504 285676
rect 197450 284200 197506 284209
rect 197450 284135 197506 284144
rect 197464 282946 197492 284135
rect 197452 282940 197504 282946
rect 197452 282882 197504 282888
rect 197450 282160 197506 282169
rect 197450 282095 197506 282104
rect 197464 281586 197492 282095
rect 197452 281580 197504 281586
rect 197452 281522 197504 281528
rect 197450 280256 197506 280265
rect 197450 280191 197452 280200
rect 197504 280191 197506 280200
rect 197452 280162 197504 280168
rect 197450 277536 197506 277545
rect 197450 277471 197506 277480
rect 197464 277438 197492 277471
rect 197452 277432 197504 277438
rect 197452 277374 197504 277380
rect 197450 275360 197506 275369
rect 197450 275295 197506 275304
rect 197464 274786 197492 275295
rect 197452 274780 197504 274786
rect 197452 274722 197504 274728
rect 197450 273320 197506 273329
rect 197450 273255 197452 273264
rect 197504 273255 197506 273264
rect 197452 273226 197504 273232
rect 197450 271280 197506 271289
rect 197450 271215 197506 271224
rect 197464 271182 197492 271215
rect 197452 271176 197504 271182
rect 197452 271118 197504 271124
rect 197450 268560 197506 268569
rect 197450 268495 197506 268504
rect 197464 268258 197492 268495
rect 197452 268252 197504 268258
rect 197452 268194 197504 268200
rect 197372 267706 197492 267734
rect 197358 266520 197414 266529
rect 197358 266455 197414 266464
rect 197372 266422 197400 266455
rect 197360 266416 197412 266422
rect 197360 266358 197412 266364
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197372 263634 197400 264415
rect 197360 263628 197412 263634
rect 197360 263570 197412 263576
rect 197358 261760 197414 261769
rect 197358 261695 197414 261704
rect 197372 260914 197400 261695
rect 197360 260908 197412 260914
rect 197360 260850 197412 260856
rect 197358 259720 197414 259729
rect 197358 259655 197414 259664
rect 197372 259486 197400 259655
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197358 257680 197414 257689
rect 197358 257615 197414 257624
rect 197372 256766 197400 257615
rect 197360 256760 197412 256766
rect 197360 256702 197412 256708
rect 197358 255640 197414 255649
rect 197358 255575 197414 255584
rect 197372 255338 197400 255575
rect 197360 255332 197412 255338
rect 197360 255274 197412 255280
rect 197358 252920 197414 252929
rect 197358 252855 197414 252864
rect 197372 252618 197400 252855
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197464 252521 197492 267706
rect 197450 252512 197506 252521
rect 197450 252447 197506 252456
rect 197358 250880 197414 250889
rect 197358 250815 197414 250824
rect 197372 249966 197400 250815
rect 197360 249960 197412 249966
rect 197360 249902 197412 249908
rect 197360 249008 197412 249014
rect 197358 248976 197360 248985
rect 197412 248976 197414 248985
rect 197358 248911 197414 248920
rect 196806 242176 196862 242185
rect 196806 242111 196862 242120
rect 196808 240100 196860 240106
rect 196808 240042 196860 240048
rect 196820 222222 196848 240042
rect 198016 237386 198044 289818
rect 198554 271280 198610 271289
rect 198554 271215 198610 271224
rect 198094 246120 198150 246129
rect 198094 246055 198150 246064
rect 198108 245682 198136 246055
rect 198096 245676 198148 245682
rect 198096 245618 198148 245624
rect 198278 244080 198334 244089
rect 198278 244015 198334 244024
rect 198292 243846 198320 244015
rect 198280 243840 198332 243846
rect 198280 243782 198332 243788
rect 198004 237380 198056 237386
rect 198004 237322 198056 237328
rect 196808 222216 196860 222222
rect 196808 222158 196860 222164
rect 198568 202434 198596 271215
rect 198556 202428 198608 202434
rect 198556 202370 198608 202376
rect 198004 189916 198056 189922
rect 198004 189858 198056 189864
rect 196808 182232 196860 182238
rect 196808 182174 196860 182180
rect 196716 181484 196768 181490
rect 196716 181426 196768 181432
rect 196716 178424 196768 178430
rect 196716 178366 196768 178372
rect 196728 155854 196756 178366
rect 196820 166870 196848 182174
rect 196900 178220 196952 178226
rect 196900 178162 196952 178168
rect 196808 166864 196860 166870
rect 196808 166806 196860 166812
rect 196912 164150 196940 178162
rect 196900 164144 196952 164150
rect 196900 164086 196952 164092
rect 196716 155848 196768 155854
rect 196716 155790 196768 155796
rect 196716 150476 196768 150482
rect 196716 150418 196768 150424
rect 196728 111790 196756 150418
rect 196808 114640 196860 114646
rect 196808 114582 196860 114588
rect 196716 111784 196768 111790
rect 196716 111726 196768 111732
rect 196820 81394 196848 114582
rect 196900 113280 196952 113286
rect 196900 113222 196952 113228
rect 196912 84114 196940 113222
rect 196900 84108 196952 84114
rect 196900 84050 196952 84056
rect 196808 81388 196860 81394
rect 196808 81330 196860 81336
rect 196624 78056 196676 78062
rect 196624 77998 196676 78004
rect 195244 42764 195296 42770
rect 195244 42706 195296 42712
rect 198016 10402 198044 189858
rect 198096 181620 198148 181626
rect 198096 181562 198148 181568
rect 198108 79422 198136 181562
rect 198660 177342 198688 303622
rect 198844 235346 198872 313375
rect 198832 235340 198884 235346
rect 198832 235282 198884 235288
rect 198936 217462 198964 324822
rect 199396 306338 199424 365978
rect 199568 362296 199620 362302
rect 199568 362238 199620 362244
rect 199474 361856 199530 361865
rect 199474 361791 199530 361800
rect 199488 333266 199516 361791
rect 199580 339114 199608 362238
rect 200776 361418 200804 371350
rect 209044 367396 209096 367402
rect 209044 367338 209096 367344
rect 209056 365770 209084 367338
rect 209044 365764 209096 365770
rect 209044 365706 209096 365712
rect 206466 364440 206522 364449
rect 206466 364375 206522 364384
rect 206480 363322 206508 364375
rect 206468 363316 206520 363322
rect 206468 363258 206520 363264
rect 204536 361820 204588 361826
rect 204536 361762 204588 361768
rect 202604 361752 202656 361758
rect 202604 361694 202656 361700
rect 200764 361412 200816 361418
rect 200764 361354 200816 361360
rect 202616 359924 202644 361694
rect 204548 359924 204576 361762
rect 206480 359924 206508 363258
rect 209056 359924 209084 365706
rect 209792 364334 209820 374002
rect 212540 371884 212592 371890
rect 212540 371826 212592 371832
rect 213828 371884 213880 371890
rect 213828 371826 213880 371832
rect 209792 364306 210648 364334
rect 210620 359938 210648 364306
rect 212552 359938 212580 371826
rect 213840 371346 213868 371826
rect 213828 371340 213880 371346
rect 213828 371282 213880 371288
rect 222856 367266 222884 389234
rect 224224 374264 224276 374270
rect 224224 374206 224276 374212
rect 223488 368552 223540 368558
rect 223488 368494 223540 368500
rect 222844 367260 222896 367266
rect 222844 367202 222896 367208
rect 216588 365764 216640 365770
rect 216588 365706 216640 365712
rect 214840 364608 214892 364614
rect 214840 364550 214892 364556
rect 210620 359910 211002 359938
rect 212552 359910 212934 359938
rect 214852 359924 214880 364550
rect 216600 360942 216628 365706
rect 219346 361856 219402 361865
rect 222856 361826 222884 367202
rect 223500 362302 223528 368494
rect 224236 364750 224264 374206
rect 224224 364744 224276 364750
rect 224224 364686 224276 364692
rect 223488 362296 223540 362302
rect 223488 362238 223540 362244
rect 223500 362114 223528 362238
rect 223500 362086 223620 362114
rect 219346 361791 219402 361800
rect 221280 361820 221332 361826
rect 216588 360936 216640 360942
rect 216588 360878 216640 360884
rect 217140 360936 217192 360942
rect 217140 360878 217192 360884
rect 217152 359938 217180 360878
rect 217152 359910 217442 359938
rect 219360 359924 219388 361791
rect 221280 361762 221332 361768
rect 222844 361820 222896 361826
rect 222844 361762 222896 361768
rect 221292 359924 221320 361762
rect 223592 359938 223620 362086
rect 224236 361826 224264 364686
rect 226996 362506 227024 400182
rect 268384 397520 268436 397526
rect 268384 397462 268436 397468
rect 231860 394732 231912 394738
rect 231860 394674 231912 394680
rect 227720 366036 227772 366042
rect 227720 365978 227772 365984
rect 226984 362500 227036 362506
rect 226984 362442 227036 362448
rect 224224 361820 224276 361826
rect 224224 361762 224276 361768
rect 225788 361820 225840 361826
rect 225788 361762 225840 361768
rect 223592 359910 223882 359938
rect 225800 359924 225828 361762
rect 227732 359924 227760 365978
rect 229652 362500 229704 362506
rect 229652 362442 229704 362448
rect 229664 359924 229692 362442
rect 231872 359938 231900 394674
rect 253204 389224 253256 389230
rect 253204 389166 253256 389172
rect 233884 378344 233936 378350
rect 233884 378286 233936 378292
rect 233896 363254 233924 378286
rect 253216 378282 253244 389166
rect 267004 388272 267056 388278
rect 267004 388214 267056 388220
rect 264244 386504 264296 386510
rect 264244 386446 264296 386452
rect 264256 379574 264284 386446
rect 263600 379568 263652 379574
rect 263600 379510 263652 379516
rect 264244 379568 264296 379574
rect 264244 379510 264296 379516
rect 244280 378276 244332 378282
rect 244280 378218 244332 378224
rect 253204 378276 253256 378282
rect 253204 378218 253256 378224
rect 244292 377466 244320 378218
rect 244280 377460 244332 377466
rect 244280 377402 244332 377408
rect 249708 376848 249760 376854
rect 244922 376816 244978 376825
rect 249708 376790 249760 376796
rect 244922 376751 244978 376760
rect 244936 369918 244964 376751
rect 242164 369912 242216 369918
rect 242164 369854 242216 369860
rect 244648 369912 244700 369918
rect 244648 369854 244700 369860
rect 244924 369912 244976 369918
rect 244924 369854 244976 369860
rect 238208 367192 238260 367198
rect 238208 367134 238260 367140
rect 233884 363248 233936 363254
rect 233884 363190 233936 363196
rect 233896 359938 233924 363190
rect 236092 363112 236144 363118
rect 236092 363054 236144 363060
rect 231872 359910 232254 359938
rect 233896 359910 234186 359938
rect 236104 359924 236132 363054
rect 238220 359938 238248 367134
rect 242176 363254 242204 369854
rect 242164 363248 242216 363254
rect 242164 363190 242216 363196
rect 242532 363248 242584 363254
rect 242532 363190 242584 363196
rect 240600 361888 240652 361894
rect 240600 361830 240652 361836
rect 238220 359910 238694 359938
rect 240612 359924 240640 361830
rect 242544 359924 242572 363190
rect 244660 359938 244688 369854
rect 247040 362976 247092 362982
rect 247040 362918 247092 362924
rect 244660 359910 245134 359938
rect 247052 359924 247080 362918
rect 249720 362234 249748 376790
rect 253216 373994 253244 378218
rect 253124 373966 253244 373994
rect 249708 362228 249760 362234
rect 249708 362170 249760 362176
rect 250904 362228 250956 362234
rect 250904 362170 250956 362176
rect 249708 361752 249760 361758
rect 248970 361720 249026 361729
rect 248970 361655 249026 361664
rect 249706 361720 249708 361729
rect 249760 361720 249762 361729
rect 249706 361655 249762 361664
rect 248984 359924 249012 361655
rect 250916 359924 250944 362170
rect 252468 361616 252520 361622
rect 252468 361558 252520 361564
rect 252480 361486 252508 361558
rect 252468 361480 252520 361486
rect 252468 361422 252520 361428
rect 253124 359938 253152 373966
rect 255320 369164 255372 369170
rect 255320 369106 255372 369112
rect 255332 368694 255360 369106
rect 255320 368688 255372 368694
rect 255320 368630 255372 368636
rect 255332 364334 255360 368630
rect 261852 366104 261904 366110
rect 261852 366046 261904 366052
rect 259368 366036 259420 366042
rect 259368 365978 259420 365984
rect 259380 364818 259408 365978
rect 258264 364812 258316 364818
rect 258264 364754 258316 364760
rect 259368 364812 259420 364818
rect 259368 364754 259420 364760
rect 257344 364472 257396 364478
rect 257344 364414 257396 364420
rect 255332 364306 255452 364334
rect 253124 359910 253506 359938
rect 255424 359924 255452 364306
rect 257356 360262 257384 364414
rect 258276 361962 258304 364754
rect 258264 361956 258316 361962
rect 258264 361898 258316 361904
rect 259920 361956 259972 361962
rect 259920 361898 259972 361904
rect 257344 360256 257396 360262
rect 257344 360198 257396 360204
rect 257356 359924 257384 360198
rect 259932 359924 259960 361898
rect 261864 359924 261892 366046
rect 263612 359938 263640 379510
rect 267016 377466 267044 388214
rect 265256 377460 265308 377466
rect 265256 377402 265308 377408
rect 267004 377460 267056 377466
rect 267004 377402 267056 377408
rect 265268 375426 265296 377402
rect 265256 375420 265308 375426
rect 265256 375362 265308 375368
rect 265268 359938 265296 375362
rect 268396 362982 268424 397462
rect 276676 396030 276704 630634
rect 299492 541686 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703254 332548 703520
rect 332508 703248 332560 703254
rect 332508 703190 332560 703196
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 364996 703050 365024 703520
rect 397472 703118 397500 703520
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 358728 703044 358780 703050
rect 358728 702986 358780 702992
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 334624 696992 334676 696998
rect 334624 696934 334676 696940
rect 320824 683188 320876 683194
rect 320824 683130 320876 683136
rect 299480 541680 299532 541686
rect 299480 541622 299532 541628
rect 286324 484424 286376 484430
rect 286324 484366 286376 484372
rect 286336 396137 286364 484366
rect 300122 396264 300178 396273
rect 300122 396199 300178 396208
rect 286322 396128 286378 396137
rect 286322 396063 286378 396072
rect 276020 396024 276072 396030
rect 276020 395966 276072 395972
rect 276664 396024 276716 396030
rect 276664 395966 276716 395972
rect 276032 395350 276060 395966
rect 276020 395344 276072 395350
rect 276020 395286 276072 395292
rect 276032 378842 276060 395286
rect 278044 393372 278096 393378
rect 278044 393314 278096 393320
rect 278056 383654 278084 393314
rect 286336 383654 286364 396063
rect 292488 395344 292540 395350
rect 292488 395286 292540 395292
rect 278056 383626 278176 383654
rect 286336 383626 286640 383654
rect 275940 378814 276060 378842
rect 269856 368824 269908 368830
rect 269856 368766 269908 368772
rect 268384 362976 268436 362982
rect 268384 362918 268436 362924
rect 268396 359938 268424 362918
rect 263612 359910 263810 359938
rect 265268 359910 265742 359938
rect 268318 359910 268424 359938
rect 269868 359938 269896 368766
rect 275940 361962 275968 378814
rect 276664 371476 276716 371482
rect 276664 371418 276716 371424
rect 274732 361956 274784 361962
rect 274732 361898 274784 361904
rect 275928 361956 275980 361962
rect 275928 361898 275980 361904
rect 272156 360256 272208 360262
rect 272156 360198 272208 360204
rect 272168 359938 272196 360198
rect 269868 359910 270250 359938
rect 271984 359924 272196 359938
rect 274744 359924 274772 361898
rect 276676 361690 276704 371418
rect 278148 361826 278176 383626
rect 282920 372836 282972 372842
rect 282920 372778 282972 372784
rect 282932 369889 282960 372778
rect 282918 369880 282974 369889
rect 282918 369815 282974 369824
rect 278136 361820 278188 361826
rect 278136 361762 278188 361768
rect 278596 361820 278648 361826
rect 278596 361762 278648 361768
rect 276664 361684 276716 361690
rect 276664 361626 276716 361632
rect 276676 359924 276704 361626
rect 278608 359924 278636 361762
rect 281172 361684 281224 361690
rect 281172 361626 281224 361632
rect 281184 359924 281212 361626
rect 282932 359938 282960 369815
rect 285036 363180 285088 363186
rect 285036 363122 285088 363128
rect 285048 360398 285076 363122
rect 285036 360392 285088 360398
rect 286612 360369 286640 383626
rect 292500 362001 292528 395286
rect 297364 382968 297416 382974
rect 297364 382910 297416 382916
rect 297376 367198 297404 382910
rect 297364 367192 297416 367198
rect 297364 367134 297416 367140
rect 295340 365968 295392 365974
rect 295340 365910 295392 365916
rect 295352 365838 295380 365910
rect 293408 365832 293460 365838
rect 293408 365774 293460 365780
rect 295340 365832 295392 365838
rect 295340 365774 295392 365780
rect 295984 365832 296036 365838
rect 295984 365774 296036 365780
rect 293420 363225 293448 365774
rect 293406 363216 293462 363225
rect 293406 363151 293462 363160
rect 292486 361992 292542 362001
rect 292486 361927 292542 361936
rect 289544 361888 289596 361894
rect 289544 361830 289596 361836
rect 289556 361554 289584 361830
rect 289544 361548 289596 361554
rect 289544 361490 289596 361496
rect 285036 360334 285088 360340
rect 286598 360360 286654 360369
rect 271984 359910 272182 359924
rect 282932 359910 283130 359938
rect 285048 359924 285076 360334
rect 286598 360295 286654 360304
rect 286612 359938 286640 360295
rect 286612 359910 286994 359938
rect 289556 359924 289584 361490
rect 292500 360233 292528 361927
rect 291474 360224 291530 360233
rect 291474 360159 291530 360168
rect 292486 360224 292542 360233
rect 292486 360159 292542 360168
rect 291488 359924 291516 360159
rect 293420 359924 293448 363151
rect 295996 359924 296024 365774
rect 297376 364334 297404 367134
rect 297376 364306 297496 364334
rect 297468 359938 297496 364306
rect 300136 361865 300164 396199
rect 316684 393440 316736 393446
rect 316684 393382 316736 393388
rect 313280 390584 313332 390590
rect 313280 390526 313332 390532
rect 301504 386436 301556 386442
rect 301504 386378 301556 386384
rect 301516 363186 301544 386378
rect 308404 377460 308456 377466
rect 308404 377402 308456 377408
rect 305092 370048 305144 370054
rect 305092 369990 305144 369996
rect 305000 365968 305052 365974
rect 305000 365910 305052 365916
rect 303528 364676 303580 364682
rect 303528 364618 303580 364624
rect 301504 363180 301556 363186
rect 301504 363122 301556 363128
rect 300768 361888 300820 361894
rect 300122 361856 300178 361865
rect 300768 361830 300820 361836
rect 300122 361791 300178 361800
rect 300136 359938 300164 361791
rect 300780 360942 300808 361830
rect 300768 360936 300820 360942
rect 300768 360878 300820 360884
rect 297468 359910 297942 359938
rect 299874 359910 300164 359938
rect 301516 359938 301544 363122
rect 303540 361622 303568 364618
rect 305012 362914 305040 365910
rect 305104 364682 305132 369990
rect 305092 364676 305144 364682
rect 305092 364618 305144 364624
rect 305644 364676 305696 364682
rect 305644 364618 305696 364624
rect 305656 364334 305684 364618
rect 305656 364306 305960 364334
rect 305000 362908 305052 362914
rect 305000 362850 305052 362856
rect 303528 361616 303580 361622
rect 303528 361558 303580 361564
rect 304356 361616 304408 361622
rect 304356 361558 304408 361564
rect 304368 360233 304396 361558
rect 304354 360224 304410 360233
rect 304354 360159 304410 360168
rect 301516 359910 301806 359938
rect 304368 359924 304396 360159
rect 305932 359938 305960 364306
rect 308416 360330 308444 377402
rect 312544 368756 312596 368762
rect 312544 368698 312596 368704
rect 310796 362024 310848 362030
rect 310796 361966 310848 361972
rect 308220 360324 308272 360330
rect 308220 360266 308272 360272
rect 308404 360324 308456 360330
rect 308404 360266 308456 360272
rect 305932 359910 306314 359938
rect 308232 359924 308260 360266
rect 310808 359924 310836 361966
rect 312556 360466 312584 368698
rect 313292 362234 313320 390526
rect 316696 383654 316724 393382
rect 316696 383626 316816 383654
rect 313280 362228 313332 362234
rect 313280 362170 313332 362176
rect 313292 362030 313320 362170
rect 313280 362024 313332 362030
rect 313280 361966 313332 361972
rect 314660 360868 314712 360874
rect 314660 360810 314712 360816
rect 312544 360460 312596 360466
rect 312544 360402 312596 360408
rect 312556 359938 312584 360402
rect 314672 359938 314700 360810
rect 312556 359910 312754 359938
rect 314672 359924 314884 359938
rect 314686 359910 314884 359924
rect 271984 359553 272012 359910
rect 314856 359553 314884 359910
rect 271970 359544 272026 359553
rect 271970 359479 272026 359488
rect 314842 359544 314898 359553
rect 316788 359530 316816 383626
rect 319536 376032 319588 376038
rect 319536 375974 319588 375980
rect 316868 361752 316920 361758
rect 316868 361694 316920 361700
rect 319258 361720 319314 361729
rect 316880 359689 316908 361694
rect 319258 361655 319314 361664
rect 316866 359680 316922 359689
rect 316866 359615 316922 359624
rect 316788 359514 317552 359530
rect 316788 359508 317564 359514
rect 316788 359502 317512 359508
rect 314842 359479 314898 359488
rect 317512 359450 317564 359456
rect 319272 359258 319300 361655
rect 319444 360392 319496 360398
rect 319444 360334 319496 360340
rect 319350 359680 319406 359689
rect 319350 359615 319406 359624
rect 319364 359417 319392 359615
rect 319350 359408 319406 359417
rect 319350 359343 319406 359352
rect 199672 359230 200054 359258
rect 319194 359230 319392 359258
rect 199672 356998 199700 359230
rect 199660 356992 199712 356998
rect 199660 356934 199712 356940
rect 319364 356697 319392 359230
rect 319350 356688 319406 356697
rect 319350 356623 319406 356632
rect 199568 339108 199620 339114
rect 199568 339050 199620 339056
rect 199476 333260 199528 333266
rect 199476 333202 199528 333208
rect 199384 306332 199436 306338
rect 199384 306274 199436 306280
rect 319350 244352 319406 244361
rect 319350 244287 319406 244296
rect 199672 240230 200054 240258
rect 199672 240174 199700 240230
rect 199660 240168 199712 240174
rect 199660 240110 199712 240116
rect 199856 239154 199884 240230
rect 318523 240094 318564 240122
rect 201926 239850 201954 240040
rect 201512 239822 201954 239850
rect 200946 239728 201002 239737
rect 200946 239663 201002 239672
rect 200960 239222 200988 239663
rect 200948 239216 201000 239222
rect 200948 239158 201000 239164
rect 199844 239148 199896 239154
rect 199844 239090 199896 239096
rect 200120 239080 200172 239086
rect 200120 239022 200172 239028
rect 200132 238474 200160 239022
rect 200120 238468 200172 238474
rect 200120 238410 200172 238416
rect 200672 238060 200724 238066
rect 200672 238002 200724 238008
rect 200684 234462 200712 238002
rect 200672 234456 200724 234462
rect 200672 234398 200724 234404
rect 201512 226098 201540 239822
rect 202236 239148 202288 239154
rect 202236 239090 202288 239096
rect 202144 239012 202196 239018
rect 202144 238954 202196 238960
rect 201592 238808 201644 238814
rect 201592 238750 201644 238756
rect 201604 238513 201632 238750
rect 201590 238504 201646 238513
rect 201590 238439 201646 238448
rect 201500 226092 201552 226098
rect 201500 226034 201552 226040
rect 198924 217456 198976 217462
rect 198924 217398 198976 217404
rect 199476 200796 199528 200802
rect 199476 200738 199528 200744
rect 199384 195288 199436 195294
rect 199384 195230 199436 195236
rect 198648 177336 198700 177342
rect 198648 177278 198700 177284
rect 198188 136672 198240 136678
rect 198188 136614 198240 136620
rect 198200 92313 198228 136614
rect 198280 116068 198332 116074
rect 198280 116010 198332 116016
rect 198186 92304 198242 92313
rect 198186 92239 198242 92248
rect 198292 90982 198320 116010
rect 198280 90976 198332 90982
rect 198280 90918 198332 90924
rect 198096 79416 198148 79422
rect 198096 79358 198148 79364
rect 199396 76702 199424 195230
rect 199488 91798 199516 200738
rect 200764 198008 200816 198014
rect 200764 197950 200816 197956
rect 200776 93673 200804 197950
rect 200948 111920 201000 111926
rect 200948 111862 201000 111868
rect 200856 100768 200908 100774
rect 200856 100710 200908 100716
rect 200762 93664 200818 93673
rect 200762 93599 200818 93608
rect 199476 91792 199528 91798
rect 199476 91734 199528 91740
rect 200868 77246 200896 100710
rect 200960 93158 200988 111862
rect 200948 93152 201000 93158
rect 200948 93094 201000 93100
rect 202156 92478 202184 238954
rect 202248 191282 202276 239090
rect 203522 237960 203578 237969
rect 203522 237895 203578 237904
rect 202788 233912 202840 233918
rect 202788 233854 202840 233860
rect 202696 226364 202748 226370
rect 202696 226306 202748 226312
rect 202708 226098 202736 226306
rect 202696 226092 202748 226098
rect 202696 226034 202748 226040
rect 202236 191276 202288 191282
rect 202236 191218 202288 191224
rect 202236 184272 202288 184278
rect 202236 184214 202288 184220
rect 202144 92472 202196 92478
rect 202144 92414 202196 92420
rect 200856 77240 200908 77246
rect 200856 77182 200908 77188
rect 199384 76696 199436 76702
rect 199384 76638 199436 76644
rect 202248 52290 202276 184214
rect 202800 182986 202828 233854
rect 202788 182980 202840 182986
rect 202788 182922 202840 182928
rect 202788 176860 202840 176866
rect 202788 176802 202840 176808
rect 202800 176662 202828 176802
rect 202788 176656 202840 176662
rect 202788 176598 202840 176604
rect 202328 138100 202380 138106
rect 202328 138042 202380 138048
rect 202340 92410 202368 138042
rect 202420 104916 202472 104922
rect 202420 104858 202472 104864
rect 202328 92404 202380 92410
rect 202328 92346 202380 92352
rect 202432 86970 202460 104858
rect 203536 95198 203564 237895
rect 203904 233918 203932 240040
rect 204168 239488 204220 239494
rect 204168 239430 204220 239436
rect 204076 238128 204128 238134
rect 204076 238070 204128 238076
rect 204088 237726 204116 238070
rect 204076 237720 204128 237726
rect 204076 237662 204128 237668
rect 203892 233912 203944 233918
rect 203892 233854 203944 233860
rect 204088 229094 204116 237662
rect 204180 237386 204208 239430
rect 204904 239216 204956 239222
rect 204904 239158 204956 239164
rect 204168 237380 204220 237386
rect 204168 237322 204220 237328
rect 204088 229066 204208 229094
rect 203616 95260 203668 95266
rect 203616 95202 203668 95208
rect 203524 95192 203576 95198
rect 203524 95134 203576 95140
rect 202420 86964 202472 86970
rect 202420 86906 202472 86912
rect 203628 75818 203656 95202
rect 204180 95130 204208 229066
rect 204916 200802 204944 239158
rect 205836 237726 205864 240040
rect 205824 237720 205876 237726
rect 205824 237662 205876 237668
rect 206282 233880 206338 233889
rect 206282 233815 206338 233824
rect 204904 200796 204956 200802
rect 204904 200738 204956 200744
rect 204996 188624 205048 188630
rect 204996 188566 205048 188572
rect 204902 177304 204958 177313
rect 204902 177239 204958 177248
rect 204168 95124 204220 95130
rect 204168 95066 204220 95072
rect 203616 75812 203668 75818
rect 203616 75754 203668 75760
rect 202236 52284 202288 52290
rect 202236 52226 202288 52232
rect 204916 25634 204944 177239
rect 205008 69834 205036 188566
rect 205088 184952 205140 184958
rect 205088 184894 205140 184900
rect 205100 157350 205128 184894
rect 205088 157344 205140 157350
rect 205088 157286 205140 157292
rect 205088 129872 205140 129878
rect 205088 129814 205140 129820
rect 205100 82822 205128 129814
rect 206296 95062 206324 233815
rect 208412 219298 208440 240040
rect 210298 239816 210326 240040
rect 212230 239816 212258 240040
rect 214806 239816 214834 240040
rect 210252 239788 210326 239816
rect 211908 239788 212258 239816
rect 213932 239788 214834 239816
rect 210252 238785 210280 239788
rect 210238 238776 210294 238785
rect 210238 238711 210294 238720
rect 209136 231192 209188 231198
rect 209136 231134 209188 231140
rect 208400 219292 208452 219298
rect 208400 219234 208452 219240
rect 208412 218074 208440 219234
rect 208400 218068 208452 218074
rect 208400 218010 208452 218016
rect 209044 181552 209096 181558
rect 207662 181520 207718 181529
rect 209044 181494 209096 181500
rect 207662 181455 207718 181464
rect 206376 176316 206428 176322
rect 206376 176258 206428 176264
rect 206284 95056 206336 95062
rect 206284 94998 206336 95004
rect 205088 82816 205140 82822
rect 205088 82758 205140 82764
rect 204996 69828 205048 69834
rect 204996 69770 205048 69776
rect 206388 46918 206416 176258
rect 206468 139460 206520 139466
rect 206468 139402 206520 139408
rect 206480 81326 206508 139402
rect 206560 100836 206612 100842
rect 206560 100778 206612 100784
rect 206572 91050 206600 100778
rect 206560 91044 206612 91050
rect 206560 90986 206612 90992
rect 207676 82210 207704 181455
rect 207756 135380 207808 135386
rect 207756 135322 207808 135328
rect 207768 91633 207796 135322
rect 207848 102264 207900 102270
rect 207848 102206 207900 102212
rect 207754 91624 207810 91633
rect 207754 91559 207810 91568
rect 207860 89729 207888 102206
rect 207846 89720 207902 89729
rect 207846 89655 207902 89664
rect 207664 82204 207716 82210
rect 207664 82146 207716 82152
rect 206468 81320 206520 81326
rect 206468 81262 206520 81268
rect 209056 79490 209084 181494
rect 209148 177410 209176 231134
rect 210252 225622 210280 238711
rect 211908 236745 211936 239788
rect 211894 236736 211950 236745
rect 211894 236671 211950 236680
rect 211804 225752 211856 225758
rect 211804 225694 211856 225700
rect 210240 225616 210292 225622
rect 210240 225558 210292 225564
rect 209228 218068 209280 218074
rect 209228 218010 209280 218016
rect 209240 181529 209268 218010
rect 211816 201006 211844 225694
rect 211908 224233 211936 236671
rect 213184 235544 213236 235550
rect 213184 235486 213236 235492
rect 211894 224224 211950 224233
rect 211894 224159 211950 224168
rect 211804 201000 211856 201006
rect 211804 200942 211856 200948
rect 213196 195294 213224 235486
rect 213932 224874 213960 239788
rect 216784 238474 216812 240040
rect 216772 238468 216824 238474
rect 216772 238410 216824 238416
rect 216784 237454 216812 238410
rect 216772 237448 216824 237454
rect 216772 237390 216824 237396
rect 217324 237448 217376 237454
rect 217324 237390 217376 237396
rect 216126 228304 216182 228313
rect 216126 228239 216182 228248
rect 213920 224868 213972 224874
rect 213920 224810 213972 224816
rect 213932 224466 213960 224810
rect 213920 224460 213972 224466
rect 213920 224402 213972 224408
rect 214564 224460 214616 224466
rect 214564 224402 214616 224408
rect 213276 201068 213328 201074
rect 213276 201010 213328 201016
rect 213184 195288 213236 195294
rect 213184 195230 213236 195236
rect 211804 192772 211856 192778
rect 211804 192714 211856 192720
rect 209226 181520 209282 181529
rect 209226 181455 209282 181464
rect 210424 180124 210476 180130
rect 210424 180066 210476 180072
rect 209136 177404 209188 177410
rect 209136 177346 209188 177352
rect 209136 150544 209188 150550
rect 209136 150486 209188 150492
rect 209148 140078 209176 150486
rect 209228 146396 209280 146402
rect 209228 146338 209280 146344
rect 209136 140072 209188 140078
rect 209136 140014 209188 140020
rect 209136 117972 209188 117978
rect 209136 117914 209188 117920
rect 209044 79484 209096 79490
rect 209044 79426 209096 79432
rect 209148 56098 209176 117914
rect 209240 89622 209268 146338
rect 210436 91050 210464 180066
rect 210516 139528 210568 139534
rect 210516 139470 210568 139476
rect 210424 91044 210476 91050
rect 210424 90986 210476 90992
rect 209228 89616 209280 89622
rect 209228 89558 209280 89564
rect 210528 88330 210556 139470
rect 210516 88324 210568 88330
rect 210516 88266 210568 88272
rect 211816 58886 211844 192714
rect 213184 185904 213236 185910
rect 213184 185846 213236 185852
rect 211896 142316 211948 142322
rect 211896 142258 211948 142264
rect 211908 86902 211936 142258
rect 212448 98048 212500 98054
rect 212448 97990 212500 97996
rect 212460 93906 212488 97990
rect 212448 93900 212500 93906
rect 212448 93842 212500 93848
rect 211896 86896 211948 86902
rect 211896 86838 211948 86844
rect 211804 58880 211856 58886
rect 211804 58822 211856 58828
rect 209136 56092 209188 56098
rect 209136 56034 209188 56040
rect 206376 46912 206428 46918
rect 206376 46854 206428 46860
rect 204904 25628 204956 25634
rect 204904 25570 204956 25576
rect 213196 13190 213224 185846
rect 213288 36718 213316 201010
rect 214576 184278 214604 224402
rect 216036 199572 216088 199578
rect 216036 199514 216088 199520
rect 214564 184272 214616 184278
rect 214564 184214 214616 184220
rect 214656 183592 214708 183598
rect 214656 183534 214708 183540
rect 214564 178152 214616 178158
rect 214564 178094 214616 178100
rect 214196 176724 214248 176730
rect 214196 176666 214248 176672
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 176225 213960 176598
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 214104 176044 214156 176050
rect 214104 175986 214156 175992
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 214012 175160 214064 175166
rect 213918 175128 213974 175137
rect 214012 175102 214064 175108
rect 213918 175063 213974 175072
rect 214024 174729 214052 175102
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 213918 173768 213974 173777
rect 213918 173703 213974 173712
rect 214116 173369 214144 175986
rect 214102 173360 214158 173369
rect 214102 173295 214158 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172417 213960 172450
rect 213918 172408 213974 172417
rect 213918 172343 213974 172352
rect 214208 172009 214236 176666
rect 214194 172000 214250 172009
rect 214194 171935 214250 171944
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170785 213960 171022
rect 214576 170921 214604 178094
rect 214562 170912 214618 170921
rect 214562 170847 214618 170856
rect 213918 170776 213974 170785
rect 213918 170711 213974 170720
rect 213920 169720 213972 169726
rect 214668 169697 214696 183534
rect 215944 183116 215996 183122
rect 215944 183058 215996 183064
rect 213920 169662 213972 169668
rect 214654 169688 214710 169697
rect 213932 169425 213960 169662
rect 214654 169623 214710 169632
rect 213918 169416 213974 169425
rect 213918 169351 213974 169360
rect 214472 169040 214524 169046
rect 214472 168982 214524 168988
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 168065 214052 168302
rect 214010 168056 214066 168065
rect 214010 167991 214066 168000
rect 214104 167000 214156 167006
rect 213918 166968 213974 166977
rect 214104 166942 214156 166948
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 213932 166870 213960 166903
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 214024 166705 214052 166874
rect 214010 166696 214066 166705
rect 214010 166631 214066 166640
rect 214116 166161 214144 166942
rect 214102 166152 214158 166161
rect 214102 166087 214158 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213918 164112 213920 164121
rect 213972 164112 213974 164121
rect 213918 164047 213974 164056
rect 214024 163441 214052 164154
rect 214010 163432 214066 163441
rect 214010 163367 214066 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 214024 162081 214052 162726
rect 214010 162072 214066 162081
rect 214010 162007 214066 162016
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 214024 160857 214052 161298
rect 214010 160848 214066 160857
rect 214010 160783 214066 160792
rect 214012 159384 214064 159390
rect 214012 159326 214064 159332
rect 213920 158704 213972 158710
rect 214024 158681 214052 159326
rect 214484 158817 214512 168982
rect 214470 158808 214526 158817
rect 214470 158743 214526 158752
rect 213920 158646 213972 158652
rect 214010 158672 214066 158681
rect 213932 158137 213960 158646
rect 214010 158607 214066 158616
rect 213918 158128 213974 158137
rect 213918 158063 213974 158072
rect 213920 157344 213972 157350
rect 213918 157312 213920 157321
rect 213972 157312 213974 157321
rect 213918 157247 213974 157256
rect 213918 155952 213974 155961
rect 213918 155887 213974 155896
rect 214012 155916 214064 155922
rect 213932 155854 213960 155887
rect 214012 155858 214064 155864
rect 213920 155848 213972 155854
rect 213920 155790 213972 155796
rect 214024 155553 214052 155858
rect 214010 155544 214066 155553
rect 214010 155479 214066 155488
rect 214564 155236 214616 155242
rect 214564 155178 214616 155184
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153504 213974 153513
rect 213918 153439 213974 153448
rect 213932 153270 213960 153439
rect 214024 153338 214052 153847
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213366 152688 213422 152697
rect 213366 152623 213422 152632
rect 213380 88058 213408 152623
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151842 213960 151943
rect 213920 151836 213972 151842
rect 213920 151778 213972 151784
rect 214010 150920 214066 150929
rect 214010 150855 214066 150864
rect 213918 150648 213974 150657
rect 213918 150583 213974 150592
rect 213932 150482 213960 150583
rect 214024 150550 214052 150855
rect 214012 150544 214064 150550
rect 214012 150486 214064 150492
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 214024 150113 214052 150350
rect 214010 150104 214066 150113
rect 214010 150039 214066 150048
rect 214576 149569 214604 155178
rect 214654 151872 214710 151881
rect 214654 151807 214710 151816
rect 214562 149560 214618 149569
rect 214562 149495 214618 149504
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 214562 148064 214618 148073
rect 214562 147999 214618 148008
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 214024 146402 214052 146639
rect 213918 146367 213974 146376
rect 214012 146396 214064 146402
rect 213932 146334 213960 146367
rect 214012 146338 214064 146344
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213920 144968 213972 144974
rect 213918 144936 213920 144945
rect 213972 144936 213974 144945
rect 213918 144871 213974 144880
rect 213920 143608 213972 143614
rect 213918 143576 213920 143585
rect 213972 143576 213974 143585
rect 213918 143511 213974 143520
rect 213918 142760 213974 142769
rect 213918 142695 213974 142704
rect 213932 142186 213960 142695
rect 214470 142352 214526 142361
rect 214470 142287 214472 142296
rect 214524 142287 214526 142296
rect 214472 142258 214524 142264
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 214024 140894 214052 141335
rect 214012 140888 214064 140894
rect 213918 140856 213974 140865
rect 214012 140830 214064 140836
rect 213918 140791 213920 140800
rect 213972 140791 213974 140800
rect 213920 140762 213972 140768
rect 214010 140040 214066 140049
rect 214010 139975 214066 139984
rect 214024 139534 214052 139975
rect 214012 139528 214064 139534
rect 213918 139496 213974 139505
rect 214012 139470 214064 139476
rect 213918 139431 213920 139440
rect 213972 139431 213974 139440
rect 213920 139402 213972 139408
rect 214010 138816 214066 138825
rect 214010 138751 214066 138760
rect 213918 138136 213974 138145
rect 214024 138106 214052 138751
rect 213918 138071 213974 138080
rect 214012 138100 214064 138106
rect 213932 138038 213960 138071
rect 214012 138042 214064 138048
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 137456 213974 137465
rect 213918 137391 213974 137400
rect 213932 136678 213960 137391
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136096 214066 136105
rect 214010 136031 214066 136040
rect 213918 135688 213974 135697
rect 213918 135623 213974 135632
rect 213932 135318 213960 135623
rect 214024 135386 214052 136031
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 213918 134056 213974 134065
rect 213918 133991 213974 134000
rect 213932 133958 213960 133991
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 214024 131238 214052 131407
rect 214012 131232 214064 131238
rect 213918 131200 213974 131209
rect 214012 131174 214064 131180
rect 213918 131135 213920 131144
rect 213972 131135 213974 131144
rect 213920 131106 213972 131112
rect 214010 130112 214066 130121
rect 214010 130047 214066 130056
rect 214024 129878 214052 130047
rect 214012 129872 214064 129878
rect 213918 129840 213974 129849
rect 214012 129814 214064 129820
rect 213918 129775 213920 129784
rect 213972 129775 213974 129784
rect 213920 129746 213972 129752
rect 213458 128888 213514 128897
rect 213458 128823 213514 128832
rect 213472 128489 213500 128823
rect 213458 128480 213514 128489
rect 213458 128415 213514 128424
rect 213918 127120 213974 127129
rect 213918 127055 213974 127064
rect 213932 127022 213960 127055
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 213918 125695 213920 125704
rect 213972 125695 213974 125704
rect 213920 125666 213972 125672
rect 214024 125662 214052 126103
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 214024 124302 214052 124743
rect 214012 124296 214064 124302
rect 213918 124264 213974 124273
rect 214012 124238 214064 124244
rect 213918 124199 213920 124208
rect 213972 124199 213974 124208
rect 213920 124170 213972 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 214024 122942 214052 123519
rect 214012 122936 214064 122942
rect 213918 122904 213974 122913
rect 214012 122878 214064 122884
rect 213918 122839 213920 122848
rect 213972 122839 213974 122848
rect 213920 122810 213972 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 213918 121816 213974 121825
rect 213918 121751 213974 121760
rect 213932 121582 213960 121751
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122159
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 213918 120456 213974 120465
rect 213918 120391 213974 120400
rect 213932 120222 213960 120391
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 120799
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213458 119096 213514 119105
rect 213458 119031 213514 119040
rect 213368 88052 213420 88058
rect 213368 87994 213420 88000
rect 213472 80034 213500 119031
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118794 213960 118895
rect 214024 118862 214052 119575
rect 214012 118856 214064 118862
rect 214012 118798 214064 118804
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 214024 117434 214052 117535
rect 214012 117428 214064 117434
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 214024 116074 214052 116175
rect 214012 116068 214064 116074
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213918 115968 213920 115977
rect 213972 115968 213974 115977
rect 213918 115903 213974 115912
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 214024 114646 214052 114951
rect 214012 114640 214064 114646
rect 213918 114608 213974 114617
rect 214012 114582 214064 114588
rect 213918 114543 213920 114552
rect 213972 114543 213974 114552
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 213920 113280 213972 113286
rect 213918 113248 213920 113257
rect 213972 113248 213974 113257
rect 214024 113218 214052 113591
rect 213918 113183 213974 113192
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 213920 111920 213972 111926
rect 213918 111888 213920 111897
rect 213972 111888 213974 111897
rect 214024 111858 214052 112231
rect 213918 111823 213974 111832
rect 214012 111852 214064 111858
rect 214012 111794 214064 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 213920 110560 213972 110566
rect 213918 110528 213920 110537
rect 213972 110528 213974 110537
rect 214024 110498 214052 110871
rect 213918 110463 213974 110472
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109168 213974 109177
rect 213918 109103 213920 109112
rect 213972 109103 213974 109112
rect 213920 109074 213972 109080
rect 214024 109070 214052 109647
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107808 213974 107817
rect 213918 107743 213920 107752
rect 213972 107743 213974 107752
rect 213920 107714 213972 107720
rect 214024 107710 214052 108287
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106448 213974 106457
rect 213918 106383 213920 106392
rect 213972 106383 213974 106392
rect 213920 106354 213972 106360
rect 214024 106350 214052 106927
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 213918 105768 213974 105777
rect 213918 105703 213974 105712
rect 213932 104922 213960 105703
rect 213920 104916 213972 104922
rect 213920 104858 213972 104864
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 214010 102504 214066 102513
rect 214010 102439 214066 102448
rect 213918 102368 213974 102377
rect 213918 102303 213974 102312
rect 213932 102270 213960 102303
rect 213920 102264 213972 102270
rect 213920 102206 213972 102212
rect 214024 102202 214052 102439
rect 214012 102196 214064 102202
rect 214012 102138 214064 102144
rect 214010 101280 214066 101289
rect 214010 101215 214066 101224
rect 213918 101144 213974 101153
rect 213918 101079 213974 101088
rect 213932 100774 213960 101079
rect 214024 100842 214052 101215
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214576 100026 214604 147999
rect 214668 144226 214696 151807
rect 214656 144220 214708 144226
rect 214656 144162 214708 144168
rect 214654 143984 214710 143993
rect 214654 143919 214710 143928
rect 214564 100020 214616 100026
rect 214564 99962 214616 99968
rect 213918 99784 213974 99793
rect 213918 99719 213974 99728
rect 213932 99414 213960 99719
rect 214010 99512 214066 99521
rect 214010 99447 214066 99456
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214024 98666 214052 99447
rect 214012 98660 214064 98666
rect 214012 98602 214064 98608
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 213918 95840 213974 95849
rect 213918 95775 213974 95784
rect 213932 95266 213960 95775
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214024 94518 214052 98359
rect 214668 97306 214696 143919
rect 214746 134192 214802 134201
rect 214746 134127 214802 134136
rect 214656 97300 214708 97306
rect 214656 97242 214708 97248
rect 214562 97064 214618 97073
rect 214562 96999 214618 97008
rect 214012 94512 214064 94518
rect 214012 94454 214064 94460
rect 214576 84182 214604 96999
rect 214760 93226 214788 134127
rect 214838 96656 214894 96665
rect 214838 96591 214894 96600
rect 214748 93220 214800 93226
rect 214748 93162 214800 93168
rect 214852 85542 214880 96591
rect 214840 85536 214892 85542
rect 214840 85478 214892 85484
rect 214564 84176 214616 84182
rect 214564 84118 214616 84124
rect 213460 80028 213512 80034
rect 213460 79970 213512 79976
rect 213276 36712 213328 36718
rect 213276 36654 213328 36660
rect 215956 17338 215984 183058
rect 216048 82278 216076 199514
rect 216140 180130 216168 228239
rect 217336 194138 217364 237390
rect 218716 234394 218744 240040
rect 220602 239834 220630 240040
rect 219440 239828 219492 239834
rect 219440 239770 219492 239776
rect 220590 239828 220642 239834
rect 220590 239770 220642 239776
rect 218704 234388 218756 234394
rect 218704 234330 218756 234336
rect 218716 198014 218744 234330
rect 219452 217938 219480 239770
rect 223224 237454 223252 240040
rect 225110 239816 225138 240040
rect 224972 239788 225138 239816
rect 221464 237448 221516 237454
rect 221464 237390 221516 237396
rect 223212 237448 223264 237454
rect 223212 237390 223264 237396
rect 220084 224324 220136 224330
rect 220084 224266 220136 224272
rect 219440 217932 219492 217938
rect 219440 217874 219492 217880
rect 218704 198008 218756 198014
rect 218704 197950 218756 197956
rect 217324 194132 217376 194138
rect 217324 194074 217376 194080
rect 220096 188630 220124 224266
rect 220728 218068 220780 218074
rect 220728 218010 220780 218016
rect 220740 217938 220768 218010
rect 220728 217932 220780 217938
rect 220728 217874 220780 217880
rect 221476 213790 221504 237390
rect 222844 235408 222896 235414
rect 222844 235350 222896 235356
rect 221464 213784 221516 213790
rect 221464 213726 221516 213732
rect 221476 189922 221504 213726
rect 221464 189916 221516 189922
rect 221464 189858 221516 189864
rect 220084 188624 220136 188630
rect 220084 188566 220136 188572
rect 222856 181626 222884 235350
rect 222936 232620 222988 232626
rect 222936 232562 222988 232568
rect 222948 224874 222976 232562
rect 222936 224868 222988 224874
rect 222936 224810 222988 224816
rect 224972 212430 225000 239788
rect 227088 235929 227116 240040
rect 229618 239816 229646 240040
rect 229112 239788 229646 239816
rect 227074 235920 227130 235929
rect 227074 235855 227130 235864
rect 229112 219366 229140 239788
rect 231596 237454 231624 240040
rect 233482 239816 233510 240040
rect 233252 239788 233510 239816
rect 229744 237448 229796 237454
rect 229744 237390 229796 237396
rect 231584 237448 231636 237454
rect 231584 237390 231636 237396
rect 229756 227594 229784 237390
rect 229744 227588 229796 227594
rect 229744 227530 229796 227536
rect 229100 219360 229152 219366
rect 229100 219302 229152 219308
rect 224960 212424 225012 212430
rect 224960 212366 225012 212372
rect 225604 212424 225656 212430
rect 225604 212366 225656 212372
rect 222936 209092 222988 209098
rect 222936 209034 222988 209040
rect 222844 181620 222896 181626
rect 222844 181562 222896 181568
rect 222948 180334 222976 209034
rect 225616 192778 225644 212366
rect 226984 209228 227036 209234
rect 226984 209170 227036 209176
rect 225604 192772 225656 192778
rect 225604 192714 225656 192720
rect 226996 184385 227024 209170
rect 228364 205080 228416 205086
rect 228364 205022 228416 205028
rect 228376 185978 228404 205022
rect 228364 185972 228416 185978
rect 228364 185914 228416 185920
rect 229756 185910 229784 227530
rect 233252 226234 233280 239788
rect 236104 237454 236132 240040
rect 238036 238882 238064 240040
rect 239922 239834 239950 240040
rect 238760 239828 238812 239834
rect 238760 239770 238812 239776
rect 239910 239828 239962 239834
rect 239910 239770 239962 239776
rect 237380 238876 237432 238882
rect 237380 238818 237432 238824
rect 238024 238876 238076 238882
rect 238024 238818 238076 238824
rect 235356 237448 235408 237454
rect 235356 237390 235408 237396
rect 236092 237448 236144 237454
rect 236092 237390 236144 237396
rect 235368 231674 235396 237390
rect 235356 231668 235408 231674
rect 235356 231610 235408 231616
rect 233240 226228 233292 226234
rect 233240 226170 233292 226176
rect 233252 225010 233280 226170
rect 233240 225004 233292 225010
rect 233240 224946 233292 224952
rect 233884 225004 233936 225010
rect 233884 224946 233936 224952
rect 232596 221536 232648 221542
rect 232596 221478 232648 221484
rect 232504 220312 232556 220318
rect 232504 220254 232556 220260
rect 230388 219360 230440 219366
rect 230388 219302 230440 219308
rect 230400 218890 230428 219302
rect 230388 218884 230440 218890
rect 230388 218826 230440 218832
rect 231124 210452 231176 210458
rect 231124 210394 231176 210400
rect 229744 185904 229796 185910
rect 229744 185846 229796 185852
rect 226982 184376 227038 184385
rect 226982 184311 227038 184320
rect 222936 180328 222988 180334
rect 222936 180270 222988 180276
rect 216128 180124 216180 180130
rect 216128 180066 216180 180072
rect 231136 178906 231164 210394
rect 232516 183025 232544 220254
rect 232608 187105 232636 221478
rect 233896 214674 233924 224946
rect 235264 214736 235316 214742
rect 235264 214678 235316 214684
rect 233884 214668 233936 214674
rect 233884 214610 233936 214616
rect 233884 203788 233936 203794
rect 233884 203730 233936 203736
rect 232688 198076 232740 198082
rect 232688 198018 232740 198024
rect 232594 187096 232650 187105
rect 232594 187031 232650 187040
rect 232502 183016 232558 183025
rect 232502 182951 232558 182960
rect 232700 181558 232728 198018
rect 232688 181552 232740 181558
rect 232688 181494 232740 181500
rect 233896 180169 233924 203730
rect 233882 180160 233938 180169
rect 233882 180095 233938 180104
rect 231124 178900 231176 178906
rect 231124 178842 231176 178848
rect 235276 175953 235304 214678
rect 235368 195498 235396 231610
rect 236644 213308 236696 213314
rect 236644 213250 236696 213256
rect 235356 195492 235408 195498
rect 235356 195434 235408 195440
rect 236656 179042 236684 213250
rect 237392 210458 237420 238818
rect 238772 223446 238800 239770
rect 241900 238754 241928 240040
rect 241900 238726 242204 238754
rect 241900 238610 241928 238726
rect 241888 238604 241940 238610
rect 241888 238546 241940 238552
rect 238760 223440 238812 223446
rect 238760 223382 238812 223388
rect 239496 223440 239548 223446
rect 239496 223382 239548 223388
rect 238024 218816 238076 218822
rect 238024 218758 238076 218764
rect 237380 210452 237432 210458
rect 237380 210394 237432 210400
rect 236644 179036 236696 179042
rect 236644 178978 236696 178984
rect 238036 177614 238064 218758
rect 239404 210520 239456 210526
rect 239404 210462 239456 210468
rect 238116 199640 238168 199646
rect 238116 199582 238168 199588
rect 238128 180402 238156 199582
rect 238116 180396 238168 180402
rect 238116 180338 238168 180344
rect 239416 180305 239444 210462
rect 239508 209098 239536 223382
rect 240784 216096 240836 216102
rect 240784 216038 240836 216044
rect 239496 209092 239548 209098
rect 239496 209034 239548 209040
rect 239402 180296 239458 180305
rect 239036 180260 239088 180266
rect 239402 180231 239458 180240
rect 239036 180202 239088 180208
rect 238024 177608 238076 177614
rect 238024 177550 238076 177556
rect 239048 177478 239076 180202
rect 240796 178974 240824 216038
rect 240876 214872 240928 214878
rect 240876 214814 240928 214820
rect 240888 192545 240916 214814
rect 240968 194064 241020 194070
rect 240968 194006 241020 194012
rect 240874 192536 240930 192545
rect 240874 192471 240930 192480
rect 240980 181694 241008 194006
rect 242176 183122 242204 238726
rect 244280 237516 244332 237522
rect 244280 237458 244332 237464
rect 244292 235890 244320 237458
rect 244280 235884 244332 235890
rect 244280 235826 244332 235832
rect 244476 234433 244504 240040
rect 246408 237522 246436 240040
rect 248294 239834 248322 240040
rect 247040 239828 247092 239834
rect 247040 239770 247092 239776
rect 248282 239828 248334 239834
rect 248282 239770 248334 239776
rect 246396 237516 246448 237522
rect 246396 237458 246448 237464
rect 246304 237448 246356 237454
rect 246304 237390 246356 237396
rect 244924 235884 244976 235890
rect 244924 235826 244976 235832
rect 244462 234424 244518 234433
rect 244462 234359 244518 234368
rect 242256 192840 242308 192846
rect 242256 192782 242308 192788
rect 242164 183116 242216 183122
rect 242164 183058 242216 183064
rect 242268 181762 242296 192782
rect 243544 190052 243596 190058
rect 243544 189994 243596 190000
rect 242256 181756 242308 181762
rect 242256 181698 242308 181704
rect 240968 181688 241020 181694
rect 240968 181630 241020 181636
rect 240784 178968 240836 178974
rect 240784 178910 240836 178916
rect 239036 177472 239088 177478
rect 239036 177414 239088 177420
rect 243556 176662 243584 189994
rect 244936 184414 244964 235826
rect 245016 227044 245068 227050
rect 245016 226986 245068 226992
rect 244924 184408 244976 184414
rect 244924 184350 244976 184356
rect 245028 178809 245056 226986
rect 246316 216578 246344 237390
rect 247052 223650 247080 239770
rect 250916 237454 250944 240040
rect 252848 238814 252876 240040
rect 252836 238808 252888 238814
rect 252836 238750 252888 238756
rect 254780 237454 254808 240040
rect 250904 237448 250956 237454
rect 250904 237390 250956 237396
rect 251824 237448 251876 237454
rect 251824 237390 251876 237396
rect 254768 237448 254820 237454
rect 254768 237390 254820 237396
rect 249800 236700 249852 236706
rect 249800 236642 249852 236648
rect 249064 229900 249116 229906
rect 249064 229842 249116 229848
rect 247040 223644 247092 223650
rect 247040 223586 247092 223592
rect 247052 223514 247080 223586
rect 247040 223508 247092 223514
rect 247040 223450 247092 223456
rect 246304 216572 246356 216578
rect 246304 216514 246356 216520
rect 245108 202360 245160 202366
rect 245108 202302 245160 202308
rect 245014 178800 245070 178809
rect 245014 178735 245070 178744
rect 243544 176656 243596 176662
rect 243544 176598 243596 176604
rect 245120 176050 245148 202302
rect 246316 178770 246344 216514
rect 246396 214804 246448 214810
rect 246396 214746 246448 214752
rect 246304 178764 246356 178770
rect 246304 178706 246356 178712
rect 246408 177682 246436 214746
rect 249076 191350 249104 229842
rect 249064 191344 249116 191350
rect 249064 191286 249116 191292
rect 249064 185836 249116 185842
rect 249064 185778 249116 185784
rect 248052 183048 248104 183054
rect 248052 182990 248104 182996
rect 247960 178832 248012 178838
rect 247960 178774 248012 178780
rect 246396 177676 246448 177682
rect 246396 177618 246448 177624
rect 245108 176044 245160 176050
rect 245108 175986 245160 175992
rect 235262 175944 235318 175953
rect 235262 175879 235318 175888
rect 247972 175817 248000 178774
rect 248064 175846 248092 182990
rect 248052 175840 248104 175846
rect 247958 175808 248014 175817
rect 248052 175782 248104 175788
rect 247958 175743 248014 175752
rect 249076 171134 249104 185778
rect 249340 180328 249392 180334
rect 249340 180270 249392 180276
rect 249248 176656 249300 176662
rect 249248 176598 249300 176604
rect 249156 175840 249208 175846
rect 249156 175782 249208 175788
rect 249168 175273 249196 175782
rect 249154 175264 249210 175273
rect 249154 175199 249210 175208
rect 249260 172825 249288 176598
rect 249352 173777 249380 180270
rect 249338 173768 249394 173777
rect 249338 173703 249394 173712
rect 249246 172816 249302 172825
rect 249246 172751 249302 172760
rect 249076 171106 249196 171134
rect 249168 149297 249196 171106
rect 249154 149288 249210 149297
rect 249154 149223 249210 149232
rect 249812 147234 249840 236642
rect 251836 228954 251864 237390
rect 255964 229900 256016 229906
rect 255964 229842 256016 229848
rect 255976 228993 256004 229842
rect 255962 228984 256018 228993
rect 251824 228948 251876 228954
rect 255962 228919 256018 228928
rect 251824 228890 251876 228896
rect 251180 224256 251232 224262
rect 251180 224198 251232 224204
rect 249984 211948 250036 211954
rect 249984 211890 250036 211896
rect 249892 187128 249944 187134
rect 249892 187070 249944 187076
rect 249904 147354 249932 187070
rect 249996 169561 250024 211890
rect 250076 188488 250128 188494
rect 250076 188430 250128 188436
rect 250088 171134 250116 188430
rect 250088 171106 250300 171134
rect 249982 169552 250038 169561
rect 249982 169487 250038 169496
rect 250272 155417 250300 171106
rect 251192 159633 251220 224198
rect 251272 191208 251324 191214
rect 251272 191150 251324 191156
rect 251178 159624 251234 159633
rect 251178 159559 251234 159568
rect 251284 158817 251312 191150
rect 251836 184346 251864 228890
rect 253940 222964 253992 222970
rect 253940 222906 253992 222912
rect 252836 207800 252888 207806
rect 252836 207742 252888 207748
rect 252744 206440 252796 206446
rect 252744 206382 252796 206388
rect 252652 193996 252704 194002
rect 252652 193938 252704 193944
rect 251364 184340 251416 184346
rect 251364 184282 251416 184288
rect 251824 184340 251876 184346
rect 251824 184282 251876 184288
rect 251376 159225 251404 184282
rect 251456 175976 251508 175982
rect 251456 175918 251508 175924
rect 251468 160177 251496 175918
rect 252468 173868 252520 173874
rect 252468 173810 252520 173816
rect 252480 173369 252508 173810
rect 252466 173360 252522 173369
rect 252466 173295 252522 173304
rect 252468 172508 252520 172514
rect 252468 172450 252520 172456
rect 252100 172440 252152 172446
rect 252480 172417 252508 172450
rect 252100 172382 252152 172388
rect 252466 172408 252522 172417
rect 252112 171465 252140 172382
rect 252466 172343 252522 172352
rect 252466 171864 252522 171873
rect 252466 171799 252522 171808
rect 252480 171562 252508 171799
rect 252468 171556 252520 171562
rect 252468 171498 252520 171504
rect 252098 171456 252154 171465
rect 252098 171391 252154 171400
rect 252376 170604 252428 170610
rect 252376 170546 252428 170552
rect 252388 170105 252416 170546
rect 252466 170504 252522 170513
rect 252466 170439 252522 170448
rect 252480 170202 252508 170439
rect 252468 170196 252520 170202
rect 252468 170138 252520 170144
rect 252374 170096 252430 170105
rect 252374 170031 252430 170040
rect 252376 169516 252428 169522
rect 252376 169458 252428 169464
rect 252388 168609 252416 169458
rect 252468 169176 252520 169182
rect 252466 169144 252468 169153
rect 252520 169144 252522 169153
rect 252466 169079 252522 169088
rect 252374 168600 252430 168609
rect 252374 168535 252430 168544
rect 252468 168360 252520 168366
rect 252468 168302 252520 168308
rect 252480 168201 252508 168302
rect 252466 168192 252522 168201
rect 252466 168127 252522 168136
rect 252466 167648 252522 167657
rect 252466 167583 252468 167592
rect 252520 167583 252522 167592
rect 252468 167554 252520 167560
rect 252376 167000 252428 167006
rect 252376 166942 252428 166948
rect 252284 166864 252336 166870
rect 252284 166806 252336 166812
rect 252296 165753 252324 166806
rect 252388 166297 252416 166942
rect 252468 166932 252520 166938
rect 252468 166874 252520 166880
rect 252480 166705 252508 166874
rect 252466 166696 252522 166705
rect 252466 166631 252522 166640
rect 252374 166288 252430 166297
rect 252374 166223 252430 166232
rect 252282 165744 252338 165753
rect 252282 165679 252338 165688
rect 252468 165572 252520 165578
rect 252468 165514 252520 165520
rect 252284 165504 252336 165510
rect 252284 165446 252336 165452
rect 252296 164393 252324 165446
rect 252480 165345 252508 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164792 252430 164801
rect 252374 164727 252430 164736
rect 252282 164384 252338 164393
rect 252282 164319 252338 164328
rect 252388 164286 252416 164727
rect 252376 164280 252428 164286
rect 252376 164222 252428 164228
rect 252468 164212 252520 164218
rect 252468 164154 252520 164160
rect 252376 164144 252428 164150
rect 252376 164086 252428 164092
rect 252388 163033 252416 164086
rect 252480 163985 252508 164154
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 252374 163024 252430 163033
rect 252374 162959 252430 162968
rect 252376 162852 252428 162858
rect 252376 162794 252428 162800
rect 252388 162081 252416 162794
rect 252468 162784 252520 162790
rect 252468 162726 252520 162732
rect 252480 162489 252508 162726
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 252374 162072 252430 162081
rect 252374 162007 252430 162016
rect 252664 161474 252692 193938
rect 252756 167249 252784 206382
rect 252742 167240 252798 167249
rect 252742 167175 252798 167184
rect 252848 161537 252876 207742
rect 252572 161446 252692 161474
rect 252834 161528 252890 161537
rect 252834 161463 252890 161472
rect 252468 161424 252520 161430
rect 252468 161366 252520 161372
rect 252480 160585 252508 161366
rect 252466 160576 252522 160585
rect 252466 160511 252522 160520
rect 251454 160168 251510 160177
rect 251454 160103 251510 160112
rect 251362 159216 251418 159225
rect 251362 159151 251418 159160
rect 251270 158808 251326 158817
rect 251270 158743 251326 158752
rect 251364 158704 251416 158710
rect 251364 158646 251416 158652
rect 251376 157865 251404 158646
rect 252192 158636 252244 158642
rect 252192 158578 252244 158584
rect 252204 158273 252232 158578
rect 252190 158264 252246 158273
rect 252190 158199 252246 158208
rect 251916 158024 251968 158030
rect 251916 157966 251968 157972
rect 251362 157856 251418 157865
rect 251362 157791 251418 157800
rect 250258 155408 250314 155417
rect 250258 155343 250314 155352
rect 251548 154556 251600 154562
rect 251548 154498 251600 154504
rect 251560 153513 251588 154498
rect 251824 153876 251876 153882
rect 251824 153818 251876 153824
rect 251546 153504 251602 153513
rect 251546 153439 251602 153448
rect 249892 147348 249944 147354
rect 249892 147290 249944 147296
rect 249812 147206 250024 147234
rect 249800 147144 249852 147150
rect 249800 147086 249852 147092
rect 249812 139505 249840 147086
rect 249996 142154 250024 147206
rect 249904 142126 250024 142154
rect 249798 139496 249854 139505
rect 249798 139431 249854 139440
rect 249904 137057 249932 142126
rect 250628 138032 250680 138038
rect 250628 137974 250680 137980
rect 249890 137048 249946 137057
rect 249890 136983 249946 136992
rect 250536 136672 250588 136678
rect 250536 136614 250588 136620
rect 217322 135552 217378 135561
rect 217322 135487 217378 135496
rect 216126 105360 216182 105369
rect 216126 105295 216182 105304
rect 216140 94897 216168 105295
rect 216126 94888 216182 94897
rect 216126 94823 216182 94832
rect 216036 82272 216088 82278
rect 216036 82214 216088 82220
rect 217336 80753 217364 135487
rect 250444 110492 250496 110498
rect 250444 110434 250496 110440
rect 249064 106344 249116 106350
rect 249064 106286 249116 106292
rect 247684 95260 247736 95266
rect 247684 95202 247736 95208
rect 242162 84960 242218 84969
rect 242162 84895 242218 84904
rect 239404 82272 239456 82278
rect 239404 82214 239456 82220
rect 232504 82204 232556 82210
rect 232504 82146 232556 82152
rect 217322 80744 217378 80753
rect 217322 80679 217378 80688
rect 215944 17332 215996 17338
rect 215944 17274 215996 17280
rect 213184 13184 213236 13190
rect 213184 13126 213236 13132
rect 198004 10396 198056 10402
rect 198004 10338 198056 10344
rect 232516 7750 232544 82146
rect 238024 79484 238076 79490
rect 238024 79426 238076 79432
rect 238036 31210 238064 79426
rect 239416 38554 239444 82214
rect 240784 72548 240836 72554
rect 240784 72490 240836 72496
rect 240796 51066 240824 72490
rect 240784 51060 240836 51066
rect 240784 51002 240836 51008
rect 240796 50590 240824 51002
rect 240140 50584 240192 50590
rect 240140 50526 240192 50532
rect 240784 50584 240836 50590
rect 240784 50526 240836 50532
rect 239404 38548 239456 38554
rect 239404 38490 239456 38496
rect 238024 31204 238076 31210
rect 238024 31146 238076 31152
rect 238024 10464 238076 10470
rect 238024 10406 238076 10412
rect 232504 7744 232556 7750
rect 232504 7686 232556 7692
rect 191104 4072 191156 4078
rect 191104 4014 191156 4020
rect 187056 3596 187108 3602
rect 187056 3538 187108 3544
rect 178684 3460 178736 3466
rect 178684 3402 178736 3408
rect 238036 3126 238064 10406
rect 239220 4820 239272 4826
rect 239220 4762 239272 4768
rect 239232 4010 239260 4762
rect 239220 4004 239272 4010
rect 239220 3946 239272 3952
rect 235816 3120 235868 3126
rect 235816 3062 235868 3068
rect 238024 3120 238076 3126
rect 238024 3062 238076 3068
rect 171968 3052 172020 3058
rect 171968 2994 172020 3000
rect 177304 3052 177356 3058
rect 177304 2994 177356 3000
rect 171980 480 172008 2994
rect 235828 480 235856 3062
rect 239232 2938 239260 3946
rect 239232 2910 239352 2938
rect 239324 480 239352 2910
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 50526
rect 242176 30326 242204 84895
rect 246304 82136 246356 82142
rect 246304 82078 246356 82084
rect 244924 79416 244976 79422
rect 244924 79358 244976 79364
rect 243542 62928 243598 62937
rect 243542 62863 243598 62872
rect 243556 52426 243584 62863
rect 243544 52420 243596 52426
rect 243544 52362 243596 52368
rect 243556 51134 243584 52362
rect 242900 51128 242952 51134
rect 242900 51070 242952 51076
rect 243544 51128 243596 51134
rect 243544 51070 243596 51076
rect 241520 30320 241572 30326
rect 241520 30262 241572 30268
rect 242164 30320 242216 30326
rect 242164 30262 242216 30268
rect 241532 16574 241560 30262
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 11830 242940 51070
rect 244936 22982 244964 79358
rect 246316 28422 246344 82078
rect 247696 53174 247724 95202
rect 247684 53168 247736 53174
rect 247684 53110 247736 53116
rect 247776 53168 247828 53174
rect 247776 53110 247828 53116
rect 247788 52290 247816 53110
rect 247040 52284 247092 52290
rect 247040 52226 247092 52232
rect 247776 52284 247828 52290
rect 247776 52226 247828 52232
rect 246304 28416 246356 28422
rect 246304 28358 246356 28364
rect 244924 22976 244976 22982
rect 244924 22918 244976 22924
rect 246304 18692 246356 18698
rect 246304 18634 246356 18640
rect 242992 17332 243044 17338
rect 242992 17274 243044 17280
rect 242900 11824 242952 11830
rect 242900 11766 242952 11772
rect 243004 6914 243032 17274
rect 246316 16574 246344 18634
rect 247052 16574 247080 52226
rect 249076 50522 249104 106286
rect 249154 96656 249210 96665
rect 249154 96591 249210 96600
rect 249168 75886 249196 96591
rect 249156 75880 249208 75886
rect 249156 75822 249208 75828
rect 249064 50516 249116 50522
rect 249064 50458 249116 50464
rect 249062 19952 249118 19961
rect 249062 19887 249118 19896
rect 246316 16546 246436 16574
rect 247052 16546 247632 16574
rect 245200 13184 245252 13190
rect 245200 13126 245252 13132
rect 244096 11824 244148 11830
rect 244096 11766 244148 11772
rect 242912 6886 243032 6914
rect 242912 480 242940 6886
rect 244108 480 244136 11766
rect 245212 480 245240 13126
rect 246408 4078 246436 16546
rect 246396 4072 246448 4078
rect 246396 4014 246448 4020
rect 246408 480 246436 4014
rect 247604 480 247632 16546
rect 249076 12374 249104 19887
rect 249064 12368 249116 12374
rect 249064 12310 249116 12316
rect 249076 11966 249104 12310
rect 248420 11960 248472 11966
rect 248420 11902 248472 11908
rect 249064 11960 249116 11966
rect 249064 11902 249116 11908
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 11902
rect 250456 6254 250484 110434
rect 250548 43518 250576 136614
rect 250640 55894 250668 137974
rect 251836 117337 251864 153818
rect 251928 129577 251956 157966
rect 252468 157344 252520 157350
rect 252466 157312 252468 157321
rect 252520 157312 252522 157321
rect 252376 157276 252428 157282
rect 252466 157247 252522 157256
rect 252376 157218 252428 157224
rect 252388 156913 252416 157218
rect 252374 156904 252430 156913
rect 252374 156839 252430 156848
rect 252572 155961 252600 161446
rect 253480 160132 253532 160138
rect 253480 160074 253532 160080
rect 252558 155952 252614 155961
rect 252558 155887 252614 155896
rect 252468 154488 252520 154494
rect 252466 154456 252468 154465
rect 252520 154456 252522 154465
rect 252376 154420 252428 154426
rect 252466 154391 252522 154400
rect 252376 154362 252428 154368
rect 252388 154057 252416 154362
rect 252374 154048 252430 154057
rect 252374 153983 252430 153992
rect 252376 153196 252428 153202
rect 252376 153138 252428 153144
rect 252284 153128 252336 153134
rect 252388 153105 252416 153138
rect 252284 153070 252336 153076
rect 252374 153096 252430 153105
rect 252296 152153 252324 153070
rect 252374 153031 252430 153040
rect 252468 153060 252520 153066
rect 252468 153002 252520 153008
rect 252480 152697 252508 153002
rect 252466 152688 252522 152697
rect 252466 152623 252522 152632
rect 252282 152144 252338 152153
rect 252282 152079 252338 152088
rect 252466 151736 252522 151745
rect 252376 151700 252428 151706
rect 252466 151671 252522 151680
rect 252376 151642 252428 151648
rect 252284 151496 252336 151502
rect 252284 151438 252336 151444
rect 252296 151201 252324 151438
rect 252282 151192 252338 151201
rect 252282 151127 252338 151136
rect 252388 150793 252416 151642
rect 252480 151638 252508 151671
rect 252468 151632 252520 151638
rect 252468 151574 252520 151580
rect 252374 150784 252430 150793
rect 252374 150719 252430 150728
rect 252468 150408 252520 150414
rect 252468 150350 252520 150356
rect 252284 150340 252336 150346
rect 252284 150282 252336 150288
rect 252296 149841 252324 150282
rect 252480 150249 252508 150350
rect 252466 150240 252522 150249
rect 252466 150175 252522 150184
rect 252282 149832 252338 149841
rect 252282 149767 252338 149776
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252376 148980 252428 148986
rect 252376 148922 252428 148928
rect 252388 148889 252416 148922
rect 252374 148880 252430 148889
rect 252374 148815 252430 148824
rect 252480 148345 252508 148990
rect 252466 148336 252522 148345
rect 252466 148271 252522 148280
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 252100 147552 252152 147558
rect 252480 147529 252508 147562
rect 252100 147494 252152 147500
rect 252466 147520 252522 147529
rect 252112 146985 252140 147494
rect 252466 147455 252522 147464
rect 252098 146976 252154 146985
rect 252098 146911 252154 146920
rect 252468 146260 252520 146266
rect 252468 146202 252520 146208
rect 252376 146192 252428 146198
rect 252376 146134 252428 146140
rect 252388 145625 252416 146134
rect 252480 146033 252508 146202
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252374 145616 252430 145625
rect 252374 145551 252430 145560
rect 252376 144900 252428 144906
rect 252376 144842 252428 144848
rect 252388 143721 252416 144842
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 144129 252508 144774
rect 252466 144120 252522 144129
rect 252466 144055 252522 144064
rect 252374 143712 252430 143721
rect 252374 143647 252430 143656
rect 253388 143608 253440 143614
rect 253388 143550 253440 143556
rect 252468 143540 252520 143546
rect 252468 143482 252520 143488
rect 252376 143472 252428 143478
rect 252376 143414 252428 143420
rect 252388 142769 252416 143414
rect 252480 143177 252508 143482
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252374 142760 252430 142769
rect 252374 142695 252430 142704
rect 253204 142180 253256 142186
rect 253204 142122 253256 142128
rect 252376 140752 252428 140758
rect 252376 140694 252428 140700
rect 252388 139913 252416 140694
rect 252468 140684 252520 140690
rect 252468 140626 252520 140632
rect 252480 140457 252508 140626
rect 252466 140448 252522 140457
rect 252466 140383 252522 140392
rect 252374 139904 252430 139913
rect 252374 139839 252430 139848
rect 252008 139800 252060 139806
rect 252008 139742 252060 139748
rect 251914 129568 251970 129577
rect 251914 129503 251970 129512
rect 251916 126880 251968 126886
rect 251916 126822 251968 126828
rect 251928 125769 251956 126822
rect 251914 125760 251970 125769
rect 251914 125695 251970 125704
rect 252020 118833 252048 139742
rect 252468 139392 252520 139398
rect 252468 139334 252520 139340
rect 252480 138553 252508 139334
rect 252466 138544 252522 138553
rect 252466 138479 252522 138488
rect 252466 138000 252522 138009
rect 252376 137964 252428 137970
rect 252466 137935 252522 137944
rect 252376 137906 252428 137912
rect 252388 137601 252416 137906
rect 252480 137902 252508 137935
rect 252468 137896 252520 137902
rect 252468 137838 252520 137844
rect 252374 137592 252430 137601
rect 252374 137527 252430 137536
rect 252100 137284 252152 137290
rect 252100 137226 252152 137232
rect 252112 132841 252140 137226
rect 252466 136640 252522 136649
rect 252192 136604 252244 136610
rect 252466 136575 252522 136584
rect 252192 136546 252244 136552
rect 252204 135697 252232 136546
rect 252376 136536 252428 136542
rect 252376 136478 252428 136484
rect 252284 136400 252336 136406
rect 252284 136342 252336 136348
rect 252190 135688 252246 135697
rect 252190 135623 252246 135632
rect 252296 135289 252324 136342
rect 252388 136241 252416 136478
rect 252480 136474 252508 136575
rect 252468 136468 252520 136474
rect 252468 136410 252520 136416
rect 252374 136232 252430 136241
rect 252374 136167 252430 136176
rect 252282 135280 252338 135289
rect 252282 135215 252338 135224
rect 252468 135244 252520 135250
rect 252468 135186 252520 135192
rect 252376 135176 252428 135182
rect 252376 135118 252428 135124
rect 252388 134337 252416 135118
rect 252480 134745 252508 135186
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252374 134328 252430 134337
rect 252374 134263 252430 134272
rect 252376 133884 252428 133890
rect 252376 133826 252428 133832
rect 252388 133385 252416 133826
rect 252468 133816 252520 133822
rect 252466 133784 252468 133793
rect 252520 133784 252522 133793
rect 252466 133719 252522 133728
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252098 132832 252154 132841
rect 252098 132767 252154 132776
rect 252468 132456 252520 132462
rect 252466 132424 252468 132433
rect 252520 132424 252522 132433
rect 252376 132388 252428 132394
rect 252466 132359 252522 132368
rect 252376 132330 252428 132336
rect 252388 131889 252416 132330
rect 252468 132320 252520 132326
rect 252468 132262 252520 132268
rect 252374 131880 252430 131889
rect 252374 131815 252430 131824
rect 252480 131481 252508 132262
rect 252466 131472 252522 131481
rect 252466 131407 252522 131416
rect 252468 131096 252520 131102
rect 252468 131038 252520 131044
rect 252376 131028 252428 131034
rect 252376 130970 252428 130976
rect 252388 130121 252416 130970
rect 252480 130937 252508 131038
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252466 130520 252522 130529
rect 252466 130455 252468 130464
rect 252520 130455 252522 130464
rect 252468 130426 252520 130432
rect 252374 130112 252430 130121
rect 252374 130047 252430 130056
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252376 129668 252428 129674
rect 252376 129610 252428 129616
rect 252192 129464 252244 129470
rect 252192 129406 252244 129412
rect 252204 126313 252232 129406
rect 252388 129169 252416 129610
rect 252374 129160 252430 129169
rect 252374 129095 252430 129104
rect 252480 128625 252508 129678
rect 252466 128616 252522 128625
rect 252466 128551 252522 128560
rect 252376 128308 252428 128314
rect 252376 128250 252428 128256
rect 252284 128240 252336 128246
rect 252284 128182 252336 128188
rect 252296 127265 252324 128182
rect 252388 127673 252416 128250
rect 252466 128208 252522 128217
rect 252466 128143 252468 128152
rect 252520 128143 252522 128152
rect 252468 128114 252520 128120
rect 252374 127664 252430 127673
rect 252374 127599 252430 127608
rect 252282 127256 252338 127265
rect 252282 127191 252338 127200
rect 252468 126948 252520 126954
rect 252468 126890 252520 126896
rect 252480 126721 252508 126890
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252190 126304 252246 126313
rect 252190 126239 252246 126248
rect 252284 125588 252336 125594
rect 252284 125530 252336 125536
rect 252296 124409 252324 125530
rect 252468 125520 252520 125526
rect 252468 125462 252520 125468
rect 252376 125452 252428 125458
rect 252376 125394 252428 125400
rect 252388 125361 252416 125394
rect 252374 125352 252430 125361
rect 252374 125287 252430 125296
rect 252376 124908 252428 124914
rect 252376 124850 252428 124856
rect 252282 124400 252338 124409
rect 252282 124335 252338 124344
rect 252388 124001 252416 124850
rect 252480 124817 252508 125462
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252374 123992 252430 124001
rect 252374 123927 252430 123936
rect 252480 123457 252508 124102
rect 252466 123448 252522 123457
rect 252466 123383 252522 123392
rect 252100 123208 252152 123214
rect 252100 123150 252152 123156
rect 252006 118824 252062 118833
rect 252006 118759 252062 118768
rect 251916 118720 251968 118726
rect 251916 118662 251968 118668
rect 251822 117328 251878 117337
rect 251822 117263 251878 117272
rect 251824 113824 251876 113830
rect 251824 113766 251876 113772
rect 251836 105641 251864 113766
rect 251822 105632 251878 105641
rect 251822 105567 251878 105576
rect 251928 103514 251956 118662
rect 252008 117972 252060 117978
rect 252008 117914 252060 117920
rect 252020 105097 252048 117914
rect 252112 106593 252140 123150
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252284 122664 252336 122670
rect 252284 122606 252336 122612
rect 252296 121553 252324 122606
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252282 121544 252338 121553
rect 252282 121479 252338 121488
rect 252468 121440 252520 121446
rect 252468 121382 252520 121388
rect 252376 121372 252428 121378
rect 252376 121314 252428 121320
rect 252284 121304 252336 121310
rect 252284 121246 252336 121252
rect 252296 121145 252324 121246
rect 252282 121136 252338 121145
rect 252282 121071 252338 121080
rect 252388 120193 252416 121314
rect 252480 120601 252508 121382
rect 252466 120592 252522 120601
rect 252466 120527 252522 120536
rect 252374 120184 252430 120193
rect 252374 120119 252430 120128
rect 252468 120080 252520 120086
rect 252468 120022 252520 120028
rect 252480 119649 252508 120022
rect 252466 119640 252522 119649
rect 252376 119604 252428 119610
rect 252466 119575 252522 119584
rect 252376 119546 252428 119552
rect 252388 119241 252416 119546
rect 252374 119232 252430 119241
rect 252374 119167 252430 119176
rect 252468 118652 252520 118658
rect 252468 118594 252520 118600
rect 252376 118584 252428 118590
rect 252376 118526 252428 118532
rect 252388 117881 252416 118526
rect 252480 118289 252508 118594
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252374 117872 252430 117881
rect 252374 117807 252430 117816
rect 252284 117292 252336 117298
rect 252284 117234 252336 117240
rect 252296 116385 252324 117234
rect 252468 117224 252520 117230
rect 252468 117166 252520 117172
rect 252376 117156 252428 117162
rect 252376 117098 252428 117104
rect 252282 116376 252338 116385
rect 252282 116311 252338 116320
rect 252388 115977 252416 117098
rect 252480 116929 252508 117166
rect 252466 116920 252522 116929
rect 252466 116855 252522 116864
rect 252374 115968 252430 115977
rect 252374 115903 252430 115912
rect 252468 115932 252520 115938
rect 252468 115874 252520 115880
rect 252376 115864 252428 115870
rect 252376 115806 252428 115812
rect 252388 115025 252416 115806
rect 252480 115433 252508 115874
rect 252466 115424 252522 115433
rect 252466 115359 252522 115368
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252284 114504 252336 114510
rect 252284 114446 252336 114452
rect 252466 114472 252522 114481
rect 252296 113529 252324 114446
rect 252466 114407 252468 114416
rect 252520 114407 252522 114416
rect 252468 114378 252520 114384
rect 252376 114368 252428 114374
rect 252376 114310 252428 114316
rect 252388 114073 252416 114310
rect 252374 114064 252430 114073
rect 252374 113999 252430 114008
rect 252282 113520 252338 113529
rect 252282 113455 252338 113464
rect 252468 113144 252520 113150
rect 252466 113112 252468 113121
rect 252520 113112 252522 113121
rect 252376 113076 252428 113082
rect 252466 113047 252522 113056
rect 252376 113018 252428 113024
rect 252388 112169 252416 113018
rect 252468 112940 252520 112946
rect 252468 112882 252520 112888
rect 252480 112713 252508 112882
rect 252466 112704 252522 112713
rect 252466 112639 252522 112648
rect 252374 112160 252430 112169
rect 252374 112095 252430 112104
rect 252468 111784 252520 111790
rect 252466 111752 252468 111761
rect 252520 111752 252522 111761
rect 252376 111716 252428 111722
rect 252466 111687 252522 111696
rect 252376 111658 252428 111664
rect 252388 111217 252416 111658
rect 252374 111208 252430 111217
rect 252374 111143 252430 111152
rect 252466 110800 252522 110809
rect 252466 110735 252522 110744
rect 252480 110702 252508 110735
rect 252468 110696 252520 110702
rect 252468 110638 252520 110644
rect 252284 110424 252336 110430
rect 252284 110366 252336 110372
rect 252296 109313 252324 110366
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252376 110288 252428 110294
rect 252480 110265 252508 110298
rect 252376 110230 252428 110236
rect 252466 110256 252522 110265
rect 252388 109857 252416 110230
rect 252466 110191 252522 110200
rect 252374 109848 252430 109857
rect 252374 109783 252430 109792
rect 252282 109304 252338 109313
rect 252282 109239 252338 109248
rect 252284 108996 252336 109002
rect 252284 108938 252336 108944
rect 252296 108361 252324 108938
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252376 108860 252428 108866
rect 252466 108831 252522 108840
rect 252376 108802 252428 108808
rect 252282 108352 252338 108361
rect 252282 108287 252338 108296
rect 252388 107953 252416 108802
rect 252374 107944 252430 107953
rect 252374 107879 252430 107888
rect 252468 107636 252520 107642
rect 252468 107578 252520 107584
rect 252376 107568 252428 107574
rect 252480 107545 252508 107578
rect 252376 107510 252428 107516
rect 252466 107536 252522 107545
rect 252388 107001 252416 107510
rect 252466 107471 252522 107480
rect 252374 106992 252430 107001
rect 252374 106927 252430 106936
rect 252098 106584 252154 106593
rect 252098 106519 252154 106528
rect 252468 106276 252520 106282
rect 252468 106218 252520 106224
rect 252480 106049 252508 106218
rect 252466 106040 252522 106049
rect 252466 105975 252522 105984
rect 252192 105664 252244 105670
rect 252192 105606 252244 105612
rect 252006 105088 252062 105097
rect 252006 105023 252062 105032
rect 251836 103486 251956 103514
rect 252204 103514 252232 105606
rect 252284 105596 252336 105602
rect 252284 105538 252336 105544
rect 252296 103737 252324 105538
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252376 104780 252428 104786
rect 252376 104722 252428 104728
rect 252388 104145 252416 104722
rect 252480 104689 252508 104790
rect 252466 104680 252522 104689
rect 252466 104615 252522 104624
rect 252374 104136 252430 104145
rect 252374 104071 252430 104080
rect 252282 103728 252338 103737
rect 252282 103663 252338 103672
rect 252204 103486 252324 103514
rect 251180 102944 251232 102950
rect 251180 102886 251232 102892
rect 251192 102241 251220 102886
rect 251178 102232 251234 102241
rect 251178 102167 251234 102176
rect 251836 98025 251864 103486
rect 252192 101448 252244 101454
rect 252192 101390 252244 101396
rect 251916 99272 251968 99278
rect 251916 99214 251968 99220
rect 251928 98569 251956 99214
rect 251914 98560 251970 98569
rect 251914 98495 251970 98504
rect 251916 98048 251968 98054
rect 251822 98016 251878 98025
rect 251916 97990 251968 97996
rect 251822 97951 251878 97960
rect 251362 97064 251418 97073
rect 251362 96999 251418 97008
rect 251270 96248 251326 96257
rect 251270 96183 251326 96192
rect 251178 80744 251234 80753
rect 251178 80679 251234 80688
rect 250628 55888 250680 55894
rect 250628 55830 250680 55836
rect 250536 43512 250588 43518
rect 250536 43454 250588 43460
rect 250536 20052 250588 20058
rect 250536 19994 250588 20000
rect 250444 6248 250496 6254
rect 250444 6190 250496 6196
rect 250548 4146 250576 19994
rect 249984 4140 250036 4146
rect 249984 4082 250036 4088
rect 250536 4140 250588 4146
rect 250536 4082 250588 4088
rect 249996 480 250024 4082
rect 251192 3534 251220 80679
rect 251284 10470 251312 96183
rect 251376 67590 251404 96999
rect 251928 84194 251956 97990
rect 252204 97617 252232 101390
rect 252296 100881 252324 103486
rect 252468 103420 252520 103426
rect 252468 103362 252520 103368
rect 252376 103352 252428 103358
rect 252376 103294 252428 103300
rect 252388 102785 252416 103294
rect 252480 103193 252508 103362
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252374 102776 252430 102785
rect 252374 102711 252430 102720
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252480 101833 252508 102070
rect 252466 101824 252522 101833
rect 252466 101759 252522 101768
rect 253216 101425 253244 142122
rect 253294 141128 253350 141137
rect 253294 141063 253350 141072
rect 253308 140865 253336 141063
rect 253294 140856 253350 140865
rect 253294 140791 253350 140800
rect 253296 136944 253348 136950
rect 253296 136886 253348 136892
rect 253308 125458 253336 136886
rect 253296 125452 253348 125458
rect 253296 125394 253348 125400
rect 253296 120148 253348 120154
rect 253296 120090 253348 120096
rect 253202 101416 253258 101425
rect 253202 101351 253258 101360
rect 252282 100872 252338 100881
rect 252282 100807 252338 100816
rect 252376 100700 252428 100706
rect 252376 100642 252428 100648
rect 252284 100564 252336 100570
rect 252284 100506 252336 100512
rect 252296 99521 252324 100506
rect 252388 99929 252416 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252480 100473 252508 100574
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252374 99920 252430 99929
rect 252374 99855 252430 99864
rect 252282 99512 252338 99521
rect 252282 99447 252338 99456
rect 252468 99340 252520 99346
rect 252468 99282 252520 99288
rect 252480 98977 252508 99282
rect 252466 98968 252522 98977
rect 252466 98903 252522 98912
rect 252190 97608 252246 97617
rect 252190 97543 252246 97552
rect 252008 97300 252060 97306
rect 252008 97242 252060 97248
rect 252020 96665 252048 97242
rect 252006 96656 252062 96665
rect 252006 96591 252062 96600
rect 253204 86284 253256 86290
rect 253204 86226 253256 86232
rect 251836 84166 251956 84194
rect 251364 67584 251416 67590
rect 251364 67526 251416 67532
rect 251836 18630 251864 84166
rect 253020 54596 253072 54602
rect 253020 54538 253072 54544
rect 253032 52358 253060 54538
rect 252652 52352 252704 52358
rect 252652 52294 252704 52300
rect 253020 52352 253072 52358
rect 253020 52294 253072 52300
rect 252560 21616 252612 21622
rect 252560 21558 252612 21564
rect 251824 18624 251876 18630
rect 251824 18566 251876 18572
rect 251272 10464 251324 10470
rect 251272 10406 251324 10412
rect 251272 3596 251324 3602
rect 251272 3538 251324 3544
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 251284 3346 251312 3538
rect 252376 3528 252428 3534
rect 252376 3470 252428 3476
rect 252572 3482 252600 21558
rect 252664 3602 252692 52294
rect 253216 22098 253244 86226
rect 253308 71058 253336 120090
rect 253400 102950 253428 143550
rect 253492 121310 253520 160074
rect 253952 158710 253980 222906
rect 256712 222154 256740 240040
rect 259242 239834 259270 240040
rect 261174 239850 261202 240040
rect 263106 239850 263134 240040
rect 265682 239850 265710 240040
rect 258080 239828 258132 239834
rect 258080 239770 258132 239776
rect 259230 239828 259282 239834
rect 259230 239770 259282 239776
rect 260852 239822 261202 239850
rect 262968 239822 263134 239850
rect 265636 239822 265710 239850
rect 267614 239834 267642 240040
rect 266360 239828 266412 239834
rect 256700 222148 256752 222154
rect 256700 222090 256752 222096
rect 256712 222018 256740 222090
rect 256700 222012 256752 222018
rect 256700 221954 256752 221960
rect 257344 222012 257396 222018
rect 257344 221954 257396 221960
rect 255320 220244 255372 220250
rect 255320 220186 255372 220192
rect 254032 206372 254084 206378
rect 254032 206314 254084 206320
rect 253940 158704 253992 158710
rect 253940 158646 253992 158652
rect 254044 148986 254072 206314
rect 254124 195356 254176 195362
rect 254124 195298 254176 195304
rect 254136 151502 254164 195298
rect 254216 192568 254268 192574
rect 254216 192510 254268 192516
rect 254228 154562 254256 192510
rect 254216 154556 254268 154562
rect 254216 154498 254268 154504
rect 254124 151496 254176 151502
rect 254124 151438 254176 151444
rect 254032 148980 254084 148986
rect 254032 148922 254084 148928
rect 255332 147558 255360 220186
rect 257356 195362 257384 221954
rect 258092 213926 258120 239770
rect 260852 224942 260880 239822
rect 262968 233034 262996 239822
rect 265636 233102 265664 239822
rect 266360 239770 266412 239776
rect 267602 239828 267654 239834
rect 269546 239816 269574 240040
rect 272122 239816 272150 240040
rect 274054 239816 274082 240040
rect 267602 239770 267654 239776
rect 269132 239788 269574 239816
rect 271892 239788 272150 239816
rect 273272 239788 274082 239816
rect 265624 233096 265676 233102
rect 265624 233038 265676 233044
rect 262956 233028 263008 233034
rect 262956 232970 263008 232976
rect 262864 229832 262916 229838
rect 262864 229774 262916 229780
rect 260840 224936 260892 224942
rect 260840 224878 260892 224884
rect 261484 224936 261536 224942
rect 261484 224878 261536 224884
rect 258172 218748 258224 218754
rect 258172 218690 258224 218696
rect 258080 213920 258132 213926
rect 258080 213862 258132 213868
rect 257344 195356 257396 195362
rect 257344 195298 257396 195304
rect 256976 192704 257028 192710
rect 256976 192646 257028 192652
rect 256792 189848 256844 189854
rect 256792 189790 256844 189796
rect 255412 187196 255464 187202
rect 255412 187138 255464 187144
rect 255424 172446 255452 187138
rect 255504 179036 255556 179042
rect 255504 178978 255556 178984
rect 255412 172440 255464 172446
rect 255412 172382 255464 172388
rect 255516 158642 255544 178978
rect 255596 177676 255648 177682
rect 255596 177618 255648 177624
rect 255504 158636 255556 158642
rect 255504 158578 255556 158584
rect 255608 150346 255636 177618
rect 256804 164150 256832 189790
rect 256882 175944 256938 175953
rect 256882 175879 256938 175888
rect 256896 170610 256924 175879
rect 256884 170604 256936 170610
rect 256884 170546 256936 170552
rect 256988 166870 257016 192646
rect 258080 177540 258132 177546
rect 258080 177482 258132 177488
rect 258092 171562 258120 177482
rect 258080 171556 258132 171562
rect 258080 171498 258132 171504
rect 258184 169522 258212 218690
rect 259368 213920 259420 213926
rect 259368 213862 259420 213868
rect 259380 211954 259408 213862
rect 259368 211948 259420 211954
rect 259368 211890 259420 211896
rect 259460 203720 259512 203726
rect 259460 203662 259512 203668
rect 258356 185632 258408 185638
rect 258356 185574 258408 185580
rect 258264 177608 258316 177614
rect 258264 177550 258316 177556
rect 258172 169516 258224 169522
rect 258172 169458 258224 169464
rect 258276 167618 258304 177550
rect 258264 167612 258316 167618
rect 258264 167554 258316 167560
rect 256976 166864 257028 166870
rect 256976 166806 257028 166812
rect 257436 165640 257488 165646
rect 257436 165582 257488 165588
rect 256792 164144 256844 164150
rect 256792 164086 256844 164092
rect 256148 151088 256200 151094
rect 256148 151030 256200 151036
rect 255596 150340 255648 150346
rect 255596 150282 255648 150288
rect 255320 147552 255372 147558
rect 255320 147494 255372 147500
rect 254768 146328 254820 146334
rect 254768 146270 254820 146276
rect 253570 141808 253626 141817
rect 253570 141743 253626 141752
rect 253584 140865 253612 141743
rect 253664 141432 253716 141438
rect 253664 141374 253716 141380
rect 253570 140856 253626 140865
rect 253570 140791 253626 140800
rect 253676 136950 253704 141374
rect 253664 136944 253716 136950
rect 253664 136886 253716 136892
rect 254676 132524 254728 132530
rect 254676 132466 254728 132472
rect 254584 125656 254636 125662
rect 254584 125598 254636 125604
rect 253480 121304 253532 121310
rect 253480 121246 253532 121252
rect 253388 102944 253440 102950
rect 253388 102886 253440 102892
rect 253388 96688 253440 96694
rect 253388 96630 253440 96636
rect 253296 71052 253348 71058
rect 253296 70994 253348 71000
rect 253400 54534 253428 96630
rect 253940 56092 253992 56098
rect 253940 56034 253992 56040
rect 253952 55894 253980 56034
rect 253940 55888 253992 55894
rect 253940 55830 253992 55836
rect 253388 54528 253440 54534
rect 253388 54470 253440 54476
rect 253204 22092 253256 22098
rect 253204 22034 253256 22040
rect 253216 21622 253244 22034
rect 253204 21616 253256 21622
rect 253204 21558 253256 21564
rect 253952 16574 253980 55830
rect 254596 21486 254624 125598
rect 254688 58818 254716 132466
rect 254780 113830 254808 146270
rect 255964 145648 256016 145654
rect 255964 145590 256016 145596
rect 254952 145580 255004 145586
rect 254952 145522 255004 145528
rect 254860 140820 254912 140826
rect 254860 140762 254912 140768
rect 254872 118726 254900 140762
rect 254964 126886 254992 145522
rect 254952 126880 255004 126886
rect 254952 126822 255004 126828
rect 254950 119368 255006 119377
rect 254950 119303 255006 119312
rect 254860 118720 254912 118726
rect 254860 118662 254912 118668
rect 254768 113824 254820 113830
rect 254768 113766 254820 113772
rect 254768 99544 254820 99550
rect 254768 99486 254820 99492
rect 254780 68338 254808 99486
rect 254964 99278 254992 119303
rect 255976 106282 256004 145590
rect 256056 139460 256108 139466
rect 256056 139402 256108 139408
rect 255964 106276 256016 106282
rect 255964 106218 256016 106224
rect 256068 101454 256096 139402
rect 256160 112946 256188 151030
rect 257344 147756 257396 147762
rect 257344 147698 257396 147704
rect 256240 147688 256292 147694
rect 256240 147630 256292 147636
rect 256252 123214 256280 147630
rect 256240 123208 256292 123214
rect 256240 123150 256292 123156
rect 256148 112940 256200 112946
rect 256148 112882 256200 112888
rect 257356 107574 257384 147698
rect 257448 129470 257476 165582
rect 257528 164892 257580 164898
rect 257528 164834 257580 164840
rect 257540 129674 257568 164834
rect 258368 143478 258396 185574
rect 259472 169182 259500 203662
rect 259552 188352 259604 188358
rect 259552 188294 259604 188300
rect 259460 169176 259512 169182
rect 259460 169118 259512 169124
rect 259368 167680 259420 167686
rect 259368 167622 259420 167628
rect 258816 158772 258868 158778
rect 258816 158714 258868 158720
rect 258724 151836 258776 151842
rect 258724 151778 258776 151784
rect 258356 143472 258408 143478
rect 258356 143414 258408 143420
rect 257620 142860 257672 142866
rect 257620 142802 257672 142808
rect 257528 129668 257580 129674
rect 257528 129610 257580 129616
rect 257436 129464 257488 129470
rect 257436 129406 257488 129412
rect 257632 111722 257660 142802
rect 257620 111716 257672 111722
rect 257620 111658 257672 111664
rect 258736 110702 258764 151778
rect 258828 119610 258856 158714
rect 258816 119604 258868 119610
rect 258816 119546 258868 119552
rect 258724 110696 258776 110702
rect 258724 110638 258776 110644
rect 257436 110560 257488 110566
rect 257436 110502 257488 110508
rect 257344 107568 257396 107574
rect 257344 107510 257396 107516
rect 256056 101448 256108 101454
rect 256056 101390 256108 101396
rect 254952 99272 255004 99278
rect 254952 99214 255004 99220
rect 255318 87544 255374 87553
rect 255318 87479 255374 87488
rect 254768 68332 254820 68338
rect 254768 68274 254820 68280
rect 254676 58812 254728 58818
rect 254676 58754 254728 58760
rect 254584 21480 254636 21486
rect 254584 21422 254636 21428
rect 255332 16574 255360 87479
rect 257448 73982 257476 110502
rect 258724 100768 258776 100774
rect 258724 100710 258776 100716
rect 257436 73976 257488 73982
rect 257436 73918 257488 73924
rect 257344 66972 257396 66978
rect 257344 66914 257396 66920
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252652 3596 252704 3602
rect 252652 3538 252704 3544
rect 251192 3318 251312 3346
rect 251192 480 251220 3318
rect 252388 480 252416 3470
rect 252572 3454 253520 3482
rect 253492 480 253520 3454
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 257356 5506 257384 66914
rect 258736 17270 258764 100710
rect 259380 97306 259408 167622
rect 259564 164286 259592 188294
rect 260932 183184 260984 183190
rect 260932 183126 260984 183132
rect 260840 181756 260892 181762
rect 260840 181698 260892 181704
rect 259644 181552 259696 181558
rect 259644 181494 259696 181500
rect 259656 170202 259684 181494
rect 260380 172576 260432 172582
rect 260380 172518 260432 172524
rect 259644 170196 259696 170202
rect 259644 170138 259696 170144
rect 260288 169788 260340 169794
rect 260288 169730 260340 169736
rect 259552 164280 259604 164286
rect 259552 164222 259604 164228
rect 260196 155984 260248 155990
rect 260196 155926 260248 155932
rect 260104 139528 260156 139534
rect 260104 139470 260156 139476
rect 259368 97300 259420 97306
rect 259368 97242 259420 97248
rect 258816 96756 258868 96762
rect 258816 96698 258868 96704
rect 258828 60042 258856 96698
rect 258816 60036 258868 60042
rect 258816 59978 258868 59984
rect 260116 49162 260144 139470
rect 260208 117162 260236 155926
rect 260300 130490 260328 169730
rect 260392 133822 260420 172518
rect 260472 158840 260524 158846
rect 260472 158782 260524 158788
rect 260484 139806 260512 158782
rect 260852 144838 260880 181698
rect 260944 172514 260972 183126
rect 261024 180396 261076 180402
rect 261024 180338 261076 180344
rect 260932 172508 260984 172514
rect 260932 172450 260984 172456
rect 261036 166938 261064 180338
rect 261496 178838 261524 224878
rect 262220 210588 262272 210594
rect 262220 210530 262272 210536
rect 261484 178832 261536 178838
rect 261484 178774 261536 178780
rect 261116 176044 261168 176050
rect 261116 175986 261168 175992
rect 261024 166932 261076 166938
rect 261024 166874 261076 166880
rect 261128 161430 261156 175986
rect 261668 171828 261720 171834
rect 261668 171770 261720 171776
rect 261484 163532 261536 163538
rect 261484 163474 261536 163480
rect 261116 161424 261168 161430
rect 261116 161366 261168 161372
rect 260840 144832 260892 144838
rect 260840 144774 260892 144780
rect 260472 139800 260524 139806
rect 260472 139742 260524 139748
rect 260380 133816 260432 133822
rect 260380 133758 260432 133764
rect 260472 133204 260524 133210
rect 260472 133146 260524 133152
rect 260288 130484 260340 130490
rect 260288 130426 260340 130432
rect 260196 117156 260248 117162
rect 260196 117098 260248 117104
rect 260196 100836 260248 100842
rect 260196 100778 260248 100784
rect 260104 49156 260156 49162
rect 260104 49098 260156 49104
rect 260208 36650 260236 100778
rect 260484 100570 260512 133146
rect 261496 128178 261524 163474
rect 261576 129804 261628 129810
rect 261576 129746 261628 129752
rect 261484 128172 261536 128178
rect 261484 128114 261536 128120
rect 261484 113212 261536 113218
rect 261484 113154 261536 113160
rect 260472 100564 260524 100570
rect 260472 100506 260524 100512
rect 260286 79384 260342 79393
rect 260286 79319 260342 79328
rect 260196 36644 260248 36650
rect 260196 36586 260248 36592
rect 260300 26217 260328 79319
rect 260840 57724 260892 57730
rect 260840 57666 260892 57672
rect 260286 26208 260342 26217
rect 260286 26143 260342 26152
rect 260300 24993 260328 26143
rect 259458 24984 259514 24993
rect 259458 24919 259514 24928
rect 260286 24984 260342 24993
rect 260286 24919 260342 24928
rect 258724 17264 258776 17270
rect 258724 17206 258776 17212
rect 258264 10396 258316 10402
rect 258264 10338 258316 10344
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257344 5500 257396 5506
rect 257344 5442 257396 5448
rect 257080 480 257108 5442
rect 258276 480 258304 10338
rect 259472 480 259500 24919
rect 260852 16574 260880 57666
rect 261496 35222 261524 113154
rect 261588 57322 261616 129746
rect 261680 99346 261708 171770
rect 262232 168366 262260 210530
rect 262404 185972 262456 185978
rect 262404 185914 262456 185920
rect 262312 181688 262364 181694
rect 262312 181630 262364 181636
rect 262220 168360 262272 168366
rect 262220 168302 262272 168308
rect 261760 154624 261812 154630
rect 261760 154566 261812 154572
rect 261772 114374 261800 154566
rect 262324 144906 262352 181630
rect 262416 165510 262444 185914
rect 262876 181558 262904 229774
rect 262968 206378 262996 232970
rect 263600 217388 263652 217394
rect 263600 217330 263652 217336
rect 262956 206372 263008 206378
rect 262956 206314 263008 206320
rect 262864 181552 262916 181558
rect 262864 181494 262916 181500
rect 263612 173874 263640 217330
rect 263692 205012 263744 205018
rect 263692 204954 263744 204960
rect 263600 173868 263652 173874
rect 263600 173810 263652 173816
rect 263048 172644 263100 172650
rect 263048 172586 263100 172592
rect 262404 165504 262456 165510
rect 262404 165446 262456 165452
rect 262956 161492 263008 161498
rect 262956 161434 263008 161440
rect 262864 154692 262916 154698
rect 262864 154634 262916 154640
rect 262312 144900 262364 144906
rect 262312 144842 262364 144848
rect 262876 115870 262904 154634
rect 262968 122670 262996 161434
rect 263060 135182 263088 172586
rect 263704 167006 263732 204954
rect 265164 196648 265216 196654
rect 265164 196590 265216 196596
rect 264980 189984 265032 189990
rect 264980 189926 265032 189932
rect 263784 185768 263836 185774
rect 263784 185710 263836 185716
rect 263692 167000 263744 167006
rect 263692 166942 263744 166948
rect 263600 157412 263652 157418
rect 263600 157354 263652 157360
rect 263612 153882 263640 157354
rect 263796 157282 263824 185710
rect 264428 168496 264480 168502
rect 264428 168438 264480 168444
rect 264244 168428 264296 168434
rect 264244 168370 264296 168376
rect 264256 158030 264284 168370
rect 264336 160200 264388 160206
rect 264336 160142 264388 160148
rect 264244 158024 264296 158030
rect 264244 157966 264296 157972
rect 263784 157276 263836 157282
rect 263784 157218 263836 157224
rect 263600 153876 263652 153882
rect 263600 153818 263652 153824
rect 264244 150476 264296 150482
rect 264244 150418 264296 150424
rect 263048 135176 263100 135182
rect 263048 135118 263100 135124
rect 262956 122664 263008 122670
rect 262956 122606 263008 122612
rect 262864 115864 262916 115870
rect 262864 115806 262916 115812
rect 261760 114368 261812 114374
rect 261760 114310 261812 114316
rect 264256 110294 264284 150418
rect 264348 121378 264376 160142
rect 264440 131034 264468 168438
rect 264992 150414 265020 189926
rect 265072 178968 265124 178974
rect 265072 178910 265124 178916
rect 264980 150408 265032 150414
rect 264980 150350 265032 150356
rect 264520 144220 264572 144226
rect 264520 144162 264572 144168
rect 264428 131028 264480 131034
rect 264428 130970 264480 130976
rect 264336 121372 264388 121378
rect 264336 121314 264388 121320
rect 264244 110288 264296 110294
rect 264244 110230 264296 110236
rect 264336 104916 264388 104922
rect 264336 104858 264388 104864
rect 264244 103624 264296 103630
rect 264244 103566 264296 103572
rect 262864 102196 262916 102202
rect 262864 102138 262916 102144
rect 261668 99340 261720 99346
rect 261668 99282 261720 99288
rect 261666 83464 261722 83473
rect 261666 83399 261722 83408
rect 261680 57934 261708 83399
rect 262218 67552 262274 67561
rect 262218 67487 262274 67496
rect 262232 66978 262260 67487
rect 262220 66972 262272 66978
rect 262220 66914 262272 66920
rect 261668 57928 261720 57934
rect 261668 57870 261720 57876
rect 261680 57730 261708 57870
rect 261668 57724 261720 57730
rect 261668 57666 261720 57672
rect 261576 57316 261628 57322
rect 261576 57258 261628 57264
rect 261484 35216 261536 35222
rect 261484 35158 261536 35164
rect 260852 16546 261800 16574
rect 260656 3324 260708 3330
rect 260656 3266 260708 3272
rect 260668 480 260696 3266
rect 261772 480 261800 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262232 354 262260 66914
rect 262312 22976 262364 22982
rect 262312 22918 262364 22924
rect 262324 3330 262352 22918
rect 262876 22846 262904 102138
rect 264256 24206 264284 103566
rect 264348 53242 264376 104858
rect 264532 104786 264560 144162
rect 265084 143546 265112 178910
rect 265176 162790 265204 196590
rect 265636 188358 265664 233038
rect 266372 209778 266400 239770
rect 266452 225684 266504 225690
rect 266452 225626 266504 225632
rect 266360 209772 266412 209778
rect 266360 209714 266412 209720
rect 266372 208418 266400 209714
rect 266360 208412 266412 208418
rect 266360 208354 266412 208360
rect 265624 188352 265676 188358
rect 265624 188294 265676 188300
rect 266360 186992 266412 186998
rect 266360 186934 266412 186940
rect 265808 173936 265860 173942
rect 265808 173878 265860 173884
rect 265164 162784 265216 162790
rect 265164 162726 265216 162732
rect 265716 149116 265768 149122
rect 265716 149058 265768 149064
rect 265072 143540 265124 143546
rect 265072 143482 265124 143488
rect 265624 135312 265676 135318
rect 265624 135254 265676 135260
rect 264520 104780 264572 104786
rect 264520 104722 264572 104728
rect 264428 103556 264480 103562
rect 264428 103498 264480 103504
rect 264440 56030 264468 103498
rect 264520 98116 264572 98122
rect 264520 98058 264572 98064
rect 264532 57254 264560 98058
rect 264980 58880 265032 58886
rect 264980 58822 265032 58828
rect 264520 57248 264572 57254
rect 264520 57190 264572 57196
rect 264428 56024 264480 56030
rect 264428 55966 264480 55972
rect 264336 53236 264388 53242
rect 264336 53178 264388 53184
rect 264244 24200 264296 24206
rect 264244 24142 264296 24148
rect 264336 24200 264388 24206
rect 264336 24142 264388 24148
rect 262864 22840 262916 22846
rect 262864 22782 262916 22788
rect 264348 16574 264376 24142
rect 264164 16546 264376 16574
rect 264164 12442 264192 16546
rect 264152 12436 264204 12442
rect 264152 12378 264204 12384
rect 262312 3324 262364 3330
rect 262312 3266 262364 3272
rect 264164 480 264192 12378
rect 262926 354 263038 480
rect 262232 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 58822
rect 265636 32502 265664 135254
rect 265728 108866 265756 149058
rect 265820 136406 265848 173878
rect 266372 162858 266400 186934
rect 266360 162852 266412 162858
rect 266360 162794 266412 162800
rect 266464 153066 266492 225626
rect 267740 213376 267792 213382
rect 267740 213318 267792 213324
rect 267004 208412 267056 208418
rect 267004 208354 267056 208360
rect 267016 175953 267044 208354
rect 267002 175944 267058 175953
rect 267002 175879 267058 175888
rect 267188 171148 267240 171154
rect 267188 171090 267240 171096
rect 267004 157480 267056 157486
rect 267004 157422 267056 157428
rect 266452 153060 266504 153066
rect 266452 153002 266504 153008
rect 265808 136400 265860 136406
rect 265808 136342 265860 136348
rect 267016 118590 267044 157422
rect 267096 153876 267148 153882
rect 267096 153818 267148 153824
rect 267004 118584 267056 118590
rect 267004 118526 267056 118532
rect 267108 114442 267136 153818
rect 267200 137290 267228 171090
rect 267752 137902 267780 213318
rect 269132 208350 269160 239788
rect 270500 233980 270552 233986
rect 270500 233922 270552 233928
rect 269120 208344 269172 208350
rect 269120 208286 269172 208292
rect 269132 207058 269160 208286
rect 269120 207052 269172 207058
rect 269120 206994 269172 207000
rect 269764 207052 269816 207058
rect 269764 206994 269816 207000
rect 269120 202224 269172 202230
rect 269120 202166 269172 202172
rect 267832 199436 267884 199442
rect 267832 199378 267884 199384
rect 267844 154494 267872 199378
rect 268476 169856 268528 169862
rect 268476 169798 268528 169804
rect 267832 154488 267884 154494
rect 267832 154430 267884 154436
rect 267740 137896 267792 137902
rect 267740 137838 267792 137844
rect 267188 137284 267240 137290
rect 267188 137226 267240 137232
rect 268384 136740 268436 136746
rect 268384 136682 268436 136688
rect 267096 114436 267148 114442
rect 267096 114378 267148 114384
rect 267004 113280 267056 113286
rect 267004 113222 267056 113228
rect 265716 108860 265768 108866
rect 265716 108802 265768 108808
rect 266360 42764 266412 42770
rect 266360 42706 266412 42712
rect 266372 42158 266400 42706
rect 266360 42152 266412 42158
rect 266360 42094 266412 42100
rect 265624 32496 265676 32502
rect 265624 32438 265676 32444
rect 266372 16574 266400 42094
rect 267016 21418 267044 113222
rect 267096 103692 267148 103698
rect 267096 103634 267148 103640
rect 267108 33862 267136 103634
rect 267188 49156 267240 49162
rect 267188 49098 267240 49104
rect 267200 42158 267228 49098
rect 267188 42152 267240 42158
rect 267188 42094 267240 42100
rect 268396 39438 268424 136682
rect 268488 132326 268516 169798
rect 269132 164218 269160 202166
rect 269212 181620 269264 181626
rect 269212 181562 269264 181568
rect 269120 164212 269172 164218
rect 269120 164154 269172 164160
rect 268568 163600 268620 163606
rect 268568 163542 268620 163548
rect 268476 132320 268528 132326
rect 268476 132262 268528 132268
rect 268580 126954 268608 163542
rect 269224 153134 269252 181562
rect 269776 175982 269804 206994
rect 269764 175976 269816 175982
rect 269764 175918 269816 175924
rect 269856 167068 269908 167074
rect 269856 167010 269908 167016
rect 269764 164280 269816 164286
rect 269764 164222 269816 164228
rect 269212 153128 269264 153134
rect 269212 153070 269264 153076
rect 268568 126948 268620 126954
rect 268568 126890 268620 126896
rect 268476 125724 268528 125730
rect 268476 125666 268528 125672
rect 268488 47734 268516 125666
rect 269776 125526 269804 164222
rect 269868 129742 269896 167010
rect 270512 165578 270540 233922
rect 271892 213858 271920 239788
rect 273272 223582 273300 239788
rect 276032 224738 276060 240040
rect 277918 239850 277946 240040
rect 280494 239850 280522 240040
rect 282426 239850 282454 240040
rect 284358 239850 284386 240040
rect 277412 239822 277946 239850
rect 280172 239822 280522 239850
rect 282196 239822 282454 239850
rect 284312 239822 284386 239850
rect 286934 239834 286962 240040
rect 285680 239828 285732 239834
rect 277412 228886 277440 239822
rect 280172 230382 280200 239822
rect 282196 238406 282224 239822
rect 282184 238400 282236 238406
rect 282184 238342 282236 238348
rect 280252 235272 280304 235278
rect 280252 235214 280304 235220
rect 280160 230376 280212 230382
rect 280160 230318 280212 230324
rect 277400 228880 277452 228886
rect 277400 228822 277452 228828
rect 277412 227798 277440 228822
rect 277400 227792 277452 227798
rect 277400 227734 277452 227740
rect 278044 227792 278096 227798
rect 278044 227734 278096 227740
rect 276020 224732 276072 224738
rect 276020 224674 276072 224680
rect 276664 224732 276716 224738
rect 276664 224674 276716 224680
rect 276676 224262 276704 224674
rect 276664 224256 276716 224262
rect 276664 224198 276716 224204
rect 273260 223576 273312 223582
rect 273260 223518 273312 223524
rect 273996 223576 274048 223582
rect 273996 223518 274048 223524
rect 271880 213852 271932 213858
rect 271880 213794 271932 213800
rect 272524 213852 272576 213858
rect 272524 213794 272576 213800
rect 272536 207806 272564 213794
rect 273904 209160 273956 209166
rect 273904 209102 273956 209108
rect 272524 207800 272576 207806
rect 272524 207742 272576 207748
rect 273260 200864 273312 200870
rect 273260 200806 273312 200812
rect 271142 195256 271198 195265
rect 271142 195191 271198 195200
rect 270590 184240 270646 184249
rect 270590 184175 270646 184184
rect 270500 165572 270552 165578
rect 270500 165514 270552 165520
rect 269948 146396 270000 146402
rect 269948 146338 270000 146344
rect 269856 129736 269908 129742
rect 269856 129678 269908 129684
rect 269764 125520 269816 125526
rect 269764 125462 269816 125468
rect 269856 116000 269908 116006
rect 269856 115942 269908 115948
rect 269764 106412 269816 106418
rect 269764 106354 269816 106360
rect 269120 66224 269172 66230
rect 269120 66166 269172 66172
rect 268568 60036 268620 60042
rect 268568 59978 268620 59984
rect 268476 47728 268528 47734
rect 268476 47670 268528 47676
rect 268384 39432 268436 39438
rect 268384 39374 268436 39380
rect 267096 33856 267148 33862
rect 267096 33798 267148 33804
rect 267740 25628 267792 25634
rect 267740 25570 267792 25576
rect 267004 21412 267056 21418
rect 267004 21354 267056 21360
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 25570
rect 268580 6905 268608 59978
rect 269132 16574 269160 66166
rect 269776 18766 269804 106354
rect 269868 50386 269896 115942
rect 269960 104854 269988 146338
rect 270604 146198 270632 184175
rect 270592 146192 270644 146198
rect 270592 146134 270644 146140
rect 270040 127628 270092 127634
rect 270040 127570 270092 127576
rect 269948 104848 270000 104854
rect 269948 104790 270000 104796
rect 270052 100638 270080 127570
rect 270040 100632 270092 100638
rect 270040 100574 270092 100580
rect 269948 78124 270000 78130
rect 269948 78066 270000 78072
rect 269960 66230 269988 78066
rect 269948 66224 270000 66230
rect 269948 66166 270000 66172
rect 269856 50380 269908 50386
rect 269856 50322 269908 50328
rect 271156 26246 271184 195191
rect 271880 191344 271932 191350
rect 271880 191286 271932 191292
rect 271328 165708 271380 165714
rect 271328 165650 271380 165656
rect 271340 128246 271368 165650
rect 271892 151706 271920 191286
rect 271972 188556 272024 188562
rect 271972 188498 272024 188504
rect 271984 153202 272012 188498
rect 273272 157350 273300 200806
rect 273352 188624 273404 188630
rect 273352 188566 273404 188572
rect 273260 157344 273312 157350
rect 273260 157286 273312 157292
rect 272708 156052 272760 156058
rect 272708 155994 272760 156000
rect 271972 153196 272024 153202
rect 271972 153138 272024 153144
rect 271880 151700 271932 151706
rect 271880 151642 271932 151648
rect 271328 128240 271380 128246
rect 271328 128182 271380 128188
rect 271236 127016 271288 127022
rect 271236 126958 271288 126964
rect 271248 31074 271276 126958
rect 272616 123004 272668 123010
rect 272616 122946 272668 122952
rect 272524 116068 272576 116074
rect 272524 116010 272576 116016
rect 271880 60784 271932 60790
rect 271880 60726 271932 60732
rect 271236 31068 271288 31074
rect 271236 31010 271288 31016
rect 271144 26240 271196 26246
rect 271144 26182 271196 26188
rect 269764 18760 269816 18766
rect 269764 18702 269816 18708
rect 271156 16574 271184 26182
rect 271892 16574 271920 60726
rect 272536 28354 272564 116010
rect 272628 61538 272656 122946
rect 272720 115938 272748 155994
rect 272800 155236 272852 155242
rect 272800 155178 272852 155184
rect 272812 117230 272840 155178
rect 273364 146266 273392 188566
rect 273352 146260 273404 146266
rect 273352 146202 273404 146208
rect 272800 117224 272852 117230
rect 272800 117166 272852 117172
rect 272708 115932 272760 115938
rect 272708 115874 272760 115880
rect 273260 64864 273312 64870
rect 273260 64806 273312 64812
rect 273272 64462 273300 64806
rect 273260 64456 273312 64462
rect 273260 64398 273312 64404
rect 272616 61532 272668 61538
rect 272616 61474 272668 61480
rect 272524 28348 272576 28354
rect 272524 28290 272576 28296
rect 269132 16546 270080 16574
rect 271156 16546 271276 16574
rect 271892 16546 272472 16574
rect 268566 6896 268622 6905
rect 268566 6831 268622 6840
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268580 354 268608 6831
rect 270052 480 270080 16546
rect 271248 480 271276 16546
rect 272444 480 272472 16546
rect 268814 354 268926 480
rect 268580 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 64398
rect 273916 47734 273944 209102
rect 274008 191214 274036 223518
rect 277400 220176 277452 220182
rect 277400 220118 277452 220124
rect 274732 216028 274784 216034
rect 274732 215970 274784 215976
rect 273996 191208 274048 191214
rect 273996 191150 274048 191156
rect 274640 178900 274692 178906
rect 274640 178842 274692 178848
rect 274088 162172 274140 162178
rect 274088 162114 274140 162120
rect 273996 128376 274048 128382
rect 273996 128318 274048 128324
rect 274008 65550 274036 128318
rect 274100 124166 274128 162114
rect 274088 124160 274140 124166
rect 274088 124102 274140 124108
rect 274086 83464 274142 83473
rect 274086 83399 274142 83408
rect 273996 65544 274048 65550
rect 273996 65486 274048 65492
rect 274100 64462 274128 83399
rect 274088 64456 274140 64462
rect 274088 64398 274140 64404
rect 274652 62082 274680 178842
rect 274744 154426 274772 215970
rect 276020 207732 276072 207738
rect 276020 207674 276072 207680
rect 274732 154420 274784 154426
rect 274732 154362 274784 154368
rect 276032 140690 276060 207674
rect 276112 203652 276164 203658
rect 276112 203594 276164 203600
rect 276124 151638 276152 203594
rect 276664 164348 276716 164354
rect 276664 164290 276716 164296
rect 276112 151632 276164 151638
rect 276112 151574 276164 151580
rect 276020 140684 276072 140690
rect 276020 140626 276072 140632
rect 275284 137284 275336 137290
rect 275284 137226 275336 137232
rect 275296 103426 275324 137226
rect 276676 125594 276704 164290
rect 276848 152516 276900 152522
rect 276848 152458 276900 152464
rect 276664 125588 276716 125594
rect 276664 125530 276716 125536
rect 276664 120216 276716 120222
rect 276664 120158 276716 120164
rect 275284 103420 275336 103426
rect 275284 103362 275336 103368
rect 275284 99476 275336 99482
rect 275284 99418 275336 99424
rect 274640 62076 274692 62082
rect 274640 62018 274692 62024
rect 274652 60790 274680 62018
rect 274640 60784 274692 60790
rect 274640 60726 274692 60732
rect 273904 47728 273956 47734
rect 273904 47670 273956 47676
rect 274640 28416 274692 28422
rect 274640 28358 274692 28364
rect 274652 16574 274680 28358
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 275296 15910 275324 99418
rect 276020 47728 276072 47734
rect 276020 47670 276072 47676
rect 276032 16574 276060 47670
rect 276676 25566 276704 120158
rect 276860 113082 276888 152458
rect 277412 136474 277440 220118
rect 277492 211880 277544 211886
rect 277492 211822 277544 211828
rect 277504 140758 277532 211822
rect 278056 196654 278084 227734
rect 278780 221604 278832 221610
rect 278780 221546 278832 221552
rect 278044 196648 278096 196654
rect 278044 196590 278096 196596
rect 278136 161560 278188 161566
rect 278136 161502 278188 161508
rect 277492 140752 277544 140758
rect 277492 140694 277544 140700
rect 277400 136468 277452 136474
rect 277400 136410 277452 136416
rect 276940 134564 276992 134570
rect 276940 134506 276992 134512
rect 276848 113076 276900 113082
rect 276848 113018 276900 113024
rect 276756 111852 276808 111858
rect 276756 111794 276808 111800
rect 276768 26994 276796 111794
rect 276952 102134 276980 134506
rect 278044 131164 278096 131170
rect 278044 131106 278096 131112
rect 276940 102128 276992 102134
rect 276940 102070 276992 102076
rect 278056 58750 278084 131106
rect 278148 122738 278176 161502
rect 278792 149054 278820 221546
rect 280160 207868 280212 207874
rect 280160 207810 280212 207816
rect 279516 149184 279568 149190
rect 279516 149126 279568 149132
rect 278780 149048 278832 149054
rect 278780 148990 278832 148996
rect 279424 124228 279476 124234
rect 279424 124170 279476 124176
rect 278136 122732 278188 122738
rect 278136 122674 278188 122680
rect 278136 114572 278188 114578
rect 278136 114514 278188 114520
rect 278044 58744 278096 58750
rect 278044 58686 278096 58692
rect 278148 47666 278176 114514
rect 278780 63572 278832 63578
rect 278780 63514 278832 63520
rect 278228 62824 278280 62830
rect 278228 62766 278280 62772
rect 278136 47660 278188 47666
rect 278136 47602 278188 47608
rect 278042 46200 278098 46209
rect 278042 46135 278098 46144
rect 278056 30326 278084 46135
rect 277400 30320 277452 30326
rect 277400 30262 277452 30268
rect 278044 30320 278096 30326
rect 278044 30262 278096 30268
rect 276846 28248 276902 28257
rect 276846 28183 276902 28192
rect 276756 26988 276808 26994
rect 276756 26930 276808 26936
rect 276664 25560 276716 25566
rect 276664 25502 276716 25508
rect 276032 16546 276704 16574
rect 275284 15904 275336 15910
rect 275284 15846 275336 15852
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 276032 480 276060 3470
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 276860 3534 276888 28183
rect 276940 26988 276992 26994
rect 276940 26930 276992 26936
rect 276952 26246 276980 26930
rect 276940 26240 276992 26246
rect 276940 26182 276992 26188
rect 277412 16574 277440 30262
rect 278240 28257 278268 62766
rect 278226 28248 278282 28257
rect 278226 28183 278282 28192
rect 278792 16574 278820 63514
rect 279436 60110 279464 124170
rect 279528 108934 279556 149126
rect 280172 147626 280200 207810
rect 280160 147620 280212 147626
rect 280160 147562 280212 147568
rect 280264 139398 280292 235214
rect 281448 230376 281500 230382
rect 281448 230318 281500 230324
rect 281460 229838 281488 230318
rect 281448 229832 281500 229838
rect 281448 229774 281500 229780
rect 281540 196852 281592 196858
rect 281540 196794 281592 196800
rect 280804 172712 280856 172718
rect 280804 172654 280856 172660
rect 280252 139392 280304 139398
rect 280252 139334 280304 139340
rect 280816 135250 280844 172654
rect 280896 143676 280948 143682
rect 280896 143618 280948 143624
rect 280804 135244 280856 135250
rect 280804 135186 280856 135192
rect 280804 124296 280856 124302
rect 280804 124238 280856 124244
rect 279516 108928 279568 108934
rect 279516 108870 279568 108876
rect 279516 78056 279568 78062
rect 279516 77998 279568 78004
rect 279528 64870 279556 77998
rect 279516 64864 279568 64870
rect 279516 64806 279568 64812
rect 279528 63578 279556 64806
rect 279516 63572 279568 63578
rect 279516 63514 279568 63520
rect 279424 60104 279476 60110
rect 279424 60046 279476 60052
rect 280816 44946 280844 124238
rect 280908 103358 280936 143618
rect 281552 137970 281580 196794
rect 281540 137964 281592 137970
rect 281540 137906 281592 137912
rect 280896 103352 280948 103358
rect 280896 103294 280948 103300
rect 280988 102264 281040 102270
rect 280988 102206 281040 102212
rect 281000 69698 281028 102206
rect 282196 96558 282224 238342
rect 284312 205630 284340 239822
rect 285680 239770 285732 239776
rect 286922 239828 286974 239834
rect 286922 239770 286974 239776
rect 285692 211138 285720 239770
rect 288912 234666 288940 240040
rect 290798 239816 290826 240040
rect 292730 239816 292758 240040
rect 289832 239788 290826 239816
rect 292592 239788 292758 239816
rect 288900 234660 288952 234666
rect 288900 234602 288952 234608
rect 289452 234660 289504 234666
rect 289452 234602 289504 234608
rect 289464 233209 289492 234602
rect 289450 233200 289506 233209
rect 289450 233135 289506 233144
rect 289832 224806 289860 239788
rect 291844 237448 291896 237454
rect 291844 237390 291896 237396
rect 291856 229094 291884 237390
rect 292592 231606 292620 239788
rect 292580 231600 292632 231606
rect 292580 231542 292632 231548
rect 292592 230994 292620 231542
rect 292580 230988 292632 230994
rect 292580 230930 292632 230936
rect 293224 230988 293276 230994
rect 293224 230930 293276 230936
rect 291856 229066 292068 229094
rect 292040 226273 292068 229066
rect 292026 226264 292082 226273
rect 292026 226199 292082 226208
rect 289820 224800 289872 224806
rect 289820 224742 289872 224748
rect 290464 224800 290516 224806
rect 290464 224742 290516 224748
rect 286324 212016 286376 212022
rect 286324 211958 286376 211964
rect 285680 211132 285732 211138
rect 285680 211074 285732 211080
rect 284300 205624 284352 205630
rect 284300 205566 284352 205572
rect 284312 205154 284340 205566
rect 284300 205148 284352 205154
rect 284300 205090 284352 205096
rect 284944 205148 284996 205154
rect 284944 205090 284996 205096
rect 284956 181626 284984 205090
rect 284944 181620 284996 181626
rect 284944 181562 284996 181568
rect 285220 174004 285272 174010
rect 285220 173946 285272 173952
rect 283656 171216 283708 171222
rect 283656 171158 283708 171164
rect 283564 135380 283616 135386
rect 283564 135322 283616 135328
rect 282276 133952 282328 133958
rect 282276 133894 282328 133900
rect 282184 96552 282236 96558
rect 282184 96494 282236 96500
rect 280988 69692 281040 69698
rect 280988 69634 281040 69640
rect 280894 62792 280950 62801
rect 280894 62727 280950 62736
rect 280908 45529 280936 62727
rect 280894 45520 280950 45529
rect 280894 45455 280950 45464
rect 280804 44940 280856 44946
rect 280804 44882 280856 44888
rect 280908 44305 280936 45455
rect 282184 44872 282236 44878
rect 282184 44814 282236 44820
rect 280158 44296 280214 44305
rect 280158 44231 280214 44240
rect 280894 44296 280950 44305
rect 280894 44231 280950 44240
rect 280172 16574 280200 44231
rect 282196 16574 282224 44814
rect 282288 24274 282316 133894
rect 282368 107908 282420 107914
rect 282368 107850 282420 107856
rect 282380 29714 282408 107850
rect 282368 29708 282420 29714
rect 282368 29650 282420 29656
rect 283576 26926 283604 135322
rect 283668 133890 283696 171158
rect 285128 169924 285180 169930
rect 285128 169866 285180 169872
rect 285036 156120 285088 156126
rect 285036 156062 285088 156068
rect 283748 142248 283800 142254
rect 283748 142190 283800 142196
rect 283656 133884 283708 133890
rect 283656 133826 283708 133832
rect 283760 105670 283788 142190
rect 284944 135448 284996 135454
rect 284944 135390 284996 135396
rect 283748 105664 283800 105670
rect 283748 105606 283800 105612
rect 283656 104984 283708 104990
rect 283656 104926 283708 104932
rect 283564 26920 283616 26926
rect 283564 26862 283616 26868
rect 282276 24268 282328 24274
rect 282276 24210 282328 24216
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276848 3528 276900 3534
rect 276848 3470 276900 3476
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281920 16546 282224 16574
rect 281920 6866 281948 16546
rect 282276 15904 282328 15910
rect 282276 15846 282328 15852
rect 281908 6860 281960 6866
rect 281908 6802 281960 6808
rect 281920 480 281948 6802
rect 282288 4010 282316 15846
rect 283104 11756 283156 11762
rect 283104 11698 283156 11704
rect 282276 4004 282328 4010
rect 282276 3946 282328 3952
rect 283116 480 283144 11698
rect 283668 8974 283696 104926
rect 284300 41404 284352 41410
rect 284300 41346 284352 41352
rect 283656 8968 283708 8974
rect 283656 8910 283708 8916
rect 284312 480 284340 41346
rect 284392 31204 284444 31210
rect 284392 31146 284444 31152
rect 284404 31074 284432 31146
rect 284392 31068 284444 31074
rect 284392 31010 284444 31016
rect 284404 6914 284432 31010
rect 284956 16046 284984 135390
rect 285048 117298 285076 156062
rect 285140 132394 285168 169866
rect 285232 136542 285260 173946
rect 285220 136536 285272 136542
rect 285220 136478 285272 136484
rect 285128 132388 285180 132394
rect 285128 132330 285180 132336
rect 285128 121508 285180 121514
rect 285128 121450 285180 121456
rect 285036 117292 285088 117298
rect 285036 117234 285088 117240
rect 285036 109064 285088 109070
rect 285036 109006 285088 109012
rect 285048 40730 285076 109006
rect 285140 76634 285168 121450
rect 285128 76628 285180 76634
rect 285128 76570 285180 76576
rect 286336 66230 286364 211958
rect 289176 198144 289228 198150
rect 289176 198086 289228 198092
rect 287796 166320 287848 166326
rect 287796 166262 287848 166268
rect 286416 162920 286468 162926
rect 286416 162862 286468 162868
rect 286428 149705 286456 162862
rect 286414 149696 286470 149705
rect 286414 149631 286470 149640
rect 286600 147824 286652 147830
rect 286600 147766 286652 147772
rect 286508 138100 286560 138106
rect 286508 138042 286560 138048
rect 286416 111920 286468 111926
rect 286416 111862 286468 111868
rect 285680 66224 285732 66230
rect 285680 66166 285732 66172
rect 286324 66224 286376 66230
rect 286324 66166 286376 66172
rect 285128 61464 285180 61470
rect 285128 61406 285180 61412
rect 285140 41410 285168 61406
rect 285128 41404 285180 41410
rect 285128 41346 285180 41352
rect 285036 40724 285088 40730
rect 285036 40666 285088 40672
rect 284944 16040 284996 16046
rect 284944 15982 284996 15988
rect 285692 6914 285720 66166
rect 286428 7614 286456 111862
rect 286520 40798 286548 138042
rect 286612 107642 286640 147766
rect 287808 128314 287836 166262
rect 287888 157548 287940 157554
rect 287888 157490 287940 157496
rect 287796 128308 287848 128314
rect 287796 128250 287848 128256
rect 287704 127084 287756 127090
rect 287704 127026 287756 127032
rect 286600 107636 286652 107642
rect 286600 107578 286652 107584
rect 287060 76628 287112 76634
rect 287060 76570 287112 76576
rect 286508 40792 286560 40798
rect 286508 40734 286560 40740
rect 287072 16574 287100 76570
rect 287072 16546 287376 16574
rect 286416 7608 286468 7614
rect 286416 7550 286468 7556
rect 284404 6886 284984 6914
rect 285692 6886 286640 6914
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 6886
rect 286612 480 286640 6886
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 6186 287744 127026
rect 287900 118658 287928 157490
rect 287980 149252 288032 149258
rect 287980 149194 288032 149200
rect 287888 118652 287940 118658
rect 287888 118594 287940 118600
rect 287796 117564 287848 117570
rect 287796 117506 287848 117512
rect 287808 10334 287836 117506
rect 287992 109002 288020 149194
rect 289084 131232 289136 131238
rect 289084 131174 289136 131180
rect 287980 108996 288032 109002
rect 287980 108938 288032 108944
rect 287888 107772 287940 107778
rect 287888 107714 287940 107720
rect 287900 43450 287928 107714
rect 287888 43444 287940 43450
rect 287888 43386 287940 43392
rect 288440 33176 288492 33182
rect 288440 33118 288492 33124
rect 288452 16574 288480 33118
rect 289096 22778 289124 131174
rect 289188 90370 289216 198086
rect 290476 185638 290504 224742
rect 291936 218884 291988 218890
rect 291936 218826 291988 218832
rect 291844 196784 291896 196790
rect 291844 196726 291896 196732
rect 290464 185632 290516 185638
rect 290464 185574 290516 185580
rect 290464 184408 290516 184414
rect 290464 184350 290516 184356
rect 289268 150544 289320 150550
rect 289268 150486 289320 150492
rect 289280 110362 289308 150486
rect 289360 110628 289412 110634
rect 289360 110570 289412 110576
rect 289268 110356 289320 110362
rect 289268 110298 289320 110304
rect 289268 96824 289320 96830
rect 289268 96766 289320 96772
rect 289176 90364 289228 90370
rect 289176 90306 289228 90312
rect 289280 46238 289308 96766
rect 289372 72622 289400 110570
rect 290476 94994 290504 184350
rect 290648 140888 290700 140894
rect 290648 140830 290700 140836
rect 290556 106480 290608 106486
rect 290556 106422 290608 106428
rect 290464 94988 290516 94994
rect 290464 94930 290516 94936
rect 289360 72616 289412 72622
rect 289360 72558 289412 72564
rect 289820 69828 289872 69834
rect 289820 69770 289872 69776
rect 289832 67590 289860 69770
rect 289820 67584 289872 67590
rect 289820 67526 289872 67532
rect 289268 46232 289320 46238
rect 289268 46174 289320 46180
rect 289174 42256 289230 42265
rect 289174 42191 289230 42200
rect 289188 34474 289216 42191
rect 289176 34468 289228 34474
rect 289176 34410 289228 34416
rect 289188 33182 289216 34410
rect 289176 33176 289228 33182
rect 289176 33118 289228 33124
rect 289084 22772 289136 22778
rect 289084 22714 289136 22720
rect 288452 16546 289032 16574
rect 287796 10328 287848 10334
rect 287796 10270 287848 10276
rect 287704 6180 287756 6186
rect 287704 6122 287756 6128
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 67526
rect 290568 54738 290596 106422
rect 290660 100706 290688 140830
rect 290648 100700 290700 100706
rect 290648 100642 290700 100648
rect 290556 54732 290608 54738
rect 290556 54674 290608 54680
rect 291200 46300 291252 46306
rect 291200 46242 291252 46248
rect 291212 16574 291240 46242
rect 291856 32502 291884 196726
rect 291948 93770 291976 218826
rect 292040 189689 292068 226199
rect 293236 203658 293264 230930
rect 295352 212498 295380 240040
rect 297284 237454 297312 240040
rect 299216 238754 299244 240040
rect 298756 238726 299244 238754
rect 297272 237448 297324 237454
rect 297272 237390 297324 237396
rect 298756 227730 298784 238726
rect 299216 238513 299244 238726
rect 299202 238504 299258 238513
rect 299202 238439 299258 238448
rect 301792 237454 301820 240040
rect 300124 237448 300176 237454
rect 300124 237390 300176 237396
rect 301780 237448 301832 237454
rect 301780 237390 301832 237396
rect 298744 227724 298796 227730
rect 298744 227666 298796 227672
rect 300136 222086 300164 237390
rect 303724 237182 303752 240040
rect 305656 238649 305684 240040
rect 305642 238640 305698 238649
rect 305642 238575 305698 238584
rect 303712 237176 303764 237182
rect 303712 237118 303764 237124
rect 303724 235278 303752 237118
rect 304906 236600 304962 236609
rect 304906 236535 304962 236544
rect 303712 235272 303764 235278
rect 303712 235214 303764 235220
rect 300124 222080 300176 222086
rect 300124 222022 300176 222028
rect 295340 212492 295392 212498
rect 295340 212434 295392 212440
rect 295352 212090 295380 212434
rect 295340 212084 295392 212090
rect 295340 212026 295392 212032
rect 295984 212084 296036 212090
rect 295984 212026 296036 212032
rect 293224 203652 293276 203658
rect 293224 203594 293276 203600
rect 295996 196790 296024 212026
rect 296076 200932 296128 200938
rect 296076 200874 296128 200880
rect 295984 196784 296036 196790
rect 295984 196726 296036 196732
rect 292026 189680 292082 189689
rect 292026 189615 292082 189624
rect 293408 158908 293460 158914
rect 293408 158850 293460 158856
rect 292028 125792 292080 125798
rect 292028 125734 292080 125740
rect 291936 93764 291988 93770
rect 291936 93706 291988 93712
rect 292040 49026 292068 125734
rect 293316 121576 293368 121582
rect 293316 121518 293368 121524
rect 293224 118720 293276 118726
rect 293224 118662 293276 118668
rect 292120 117428 292172 117434
rect 292120 117370 292172 117376
rect 292132 66910 292160 117370
rect 292580 69760 292632 69766
rect 292580 69702 292632 69708
rect 292592 68950 292620 69702
rect 292580 68944 292632 68950
rect 292580 68886 292632 68892
rect 292120 66904 292172 66910
rect 292120 66846 292172 66852
rect 292028 49020 292080 49026
rect 292028 48962 292080 48968
rect 291844 32496 291896 32502
rect 291844 32438 291896 32444
rect 292592 16574 292620 68886
rect 293236 64190 293264 118662
rect 293328 68406 293356 121518
rect 293420 120086 293448 158850
rect 294788 139596 294840 139602
rect 294788 139538 294840 139544
rect 294604 129872 294656 129878
rect 294604 129814 294656 129820
rect 293408 120080 293460 120086
rect 293408 120022 293460 120028
rect 293316 68400 293368 68406
rect 293316 68342 293368 68348
rect 293224 64184 293276 64190
rect 293224 64126 293276 64132
rect 293960 32496 294012 32502
rect 293960 32438 294012 32444
rect 293972 16574 294000 32438
rect 294616 19990 294644 129814
rect 294696 109132 294748 109138
rect 294696 109074 294748 109080
rect 294708 32434 294736 109074
rect 294800 76566 294828 139538
rect 295984 135516 296036 135522
rect 295984 135458 296036 135464
rect 294788 76560 294840 76566
rect 294788 76502 294840 76508
rect 295340 36712 295392 36718
rect 295340 36654 295392 36660
rect 294696 32428 294748 32434
rect 294696 32370 294748 32376
rect 294604 19984 294656 19990
rect 294604 19926 294656 19932
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 291396 480 291424 16546
rect 292580 3120 292632 3126
rect 292580 3062 292632 3068
rect 292592 480 292620 3062
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295352 354 295380 36654
rect 295432 35216 295484 35222
rect 295430 35184 295432 35193
rect 295484 35184 295486 35193
rect 295430 35119 295486 35128
rect 295444 3126 295472 35119
rect 295996 29646 296024 135458
rect 296088 94926 296116 200874
rect 300136 199442 300164 222022
rect 300124 199436 300176 199442
rect 300124 199378 300176 199384
rect 296260 174072 296312 174078
rect 296260 174014 296312 174020
rect 296168 144968 296220 144974
rect 296168 144910 296220 144916
rect 296180 105602 296208 144910
rect 296272 136610 296300 174014
rect 297364 169040 297416 169046
rect 297364 168982 297416 168988
rect 296260 136604 296312 136610
rect 296260 136546 296312 136552
rect 297376 131102 297404 168982
rect 300216 167748 300268 167754
rect 300216 167690 300268 167696
rect 298744 153264 298796 153270
rect 298744 153206 298796 153212
rect 297456 132592 297508 132598
rect 297456 132534 297508 132540
rect 297364 131096 297416 131102
rect 297364 131038 297416 131044
rect 297364 128444 297416 128450
rect 297364 128386 297416 128392
rect 296260 114640 296312 114646
rect 296260 114582 296312 114588
rect 296168 105596 296220 105602
rect 296168 105538 296220 105544
rect 296168 102332 296220 102338
rect 296168 102274 296220 102280
rect 296076 94920 296128 94926
rect 296076 94862 296128 94868
rect 296180 36582 296208 102274
rect 296272 53106 296300 114582
rect 296260 53100 296312 53106
rect 296260 53042 296312 53048
rect 296720 38616 296772 38622
rect 296720 38558 296772 38564
rect 296168 36576 296220 36582
rect 296168 36518 296220 36524
rect 295984 29640 296036 29646
rect 295984 29582 296036 29588
rect 296732 16574 296760 38558
rect 296732 16546 297312 16574
rect 295432 3120 295484 3126
rect 295432 3062 295484 3068
rect 297284 480 297312 16546
rect 297376 2106 297404 128386
rect 297468 55962 297496 132534
rect 297548 129940 297600 129946
rect 297548 129882 297600 129888
rect 297560 77994 297588 129882
rect 298756 114510 298784 153206
rect 300124 134020 300176 134026
rect 300124 133962 300176 133968
rect 298836 122936 298888 122942
rect 298836 122878 298888 122884
rect 298744 114504 298796 114510
rect 298744 114446 298796 114452
rect 298744 100904 298796 100910
rect 298744 100846 298796 100852
rect 297548 77988 297600 77994
rect 297548 77930 297600 77936
rect 297548 69692 297600 69698
rect 297548 69634 297600 69640
rect 297456 55956 297508 55962
rect 297456 55898 297508 55904
rect 297560 38622 297588 69634
rect 297548 38616 297600 38622
rect 297548 38558 297600 38564
rect 298100 18080 298152 18086
rect 298100 18022 298152 18028
rect 297364 2100 297416 2106
rect 297364 2042 297416 2048
rect 296046 354 296158 480
rect 295352 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 18022
rect 298756 15978 298784 100846
rect 298848 62898 298876 122878
rect 298836 62892 298888 62898
rect 298836 62834 298888 62840
rect 300136 50454 300164 133962
rect 300228 132462 300256 167690
rect 304264 161628 304316 161634
rect 304264 161570 304316 161576
rect 301504 160268 301556 160274
rect 301504 160210 301556 160216
rect 300308 146464 300360 146470
rect 300308 146406 300360 146412
rect 300216 132456 300268 132462
rect 300216 132398 300268 132404
rect 300320 117978 300348 146406
rect 301516 121446 301544 160210
rect 302976 153332 303028 153338
rect 302976 153274 303028 153280
rect 301596 131300 301648 131306
rect 301596 131242 301648 131248
rect 301504 121440 301556 121446
rect 301504 121382 301556 121388
rect 300400 118788 300452 118794
rect 300400 118730 300452 118736
rect 300308 117972 300360 117978
rect 300308 117914 300360 117920
rect 300308 113348 300360 113354
rect 300308 113290 300360 113296
rect 300216 105052 300268 105058
rect 300216 104994 300268 105000
rect 300228 51746 300256 104994
rect 300320 61402 300348 113290
rect 300412 75274 300440 118730
rect 301504 116136 301556 116142
rect 301504 116078 301556 116084
rect 300400 75268 300452 75274
rect 300400 75210 300452 75216
rect 300308 61396 300360 61402
rect 300308 61338 300360 61344
rect 300216 51740 300268 51746
rect 300216 51682 300268 51688
rect 300124 50448 300176 50454
rect 300124 50390 300176 50396
rect 300674 39536 300730 39545
rect 299572 39500 299624 39506
rect 300674 39471 300676 39480
rect 299572 39442 299624 39448
rect 300728 39471 300730 39480
rect 300676 39442 300728 39448
rect 299480 38004 299532 38010
rect 299480 37946 299532 37952
rect 298836 28280 298888 28286
rect 298836 28222 298888 28228
rect 298848 19310 298876 28222
rect 298836 19304 298888 19310
rect 298836 19246 298888 19252
rect 298848 18086 298876 19246
rect 298836 18080 298888 18086
rect 298836 18022 298888 18028
rect 298744 15972 298796 15978
rect 298744 15914 298796 15920
rect 299492 3482 299520 37946
rect 299584 3641 299612 39442
rect 301516 13122 301544 116078
rect 301608 33794 301636 131242
rect 302884 124364 302936 124370
rect 302884 124306 302936 124312
rect 301688 117496 301740 117502
rect 301688 117438 301740 117444
rect 301700 72486 301728 117438
rect 301688 72480 301740 72486
rect 301688 72422 301740 72428
rect 302240 39432 302292 39438
rect 302240 39374 302292 39380
rect 302252 38554 302280 39374
rect 302240 38548 302292 38554
rect 302240 38490 302292 38496
rect 301596 33788 301648 33794
rect 301596 33730 301648 33736
rect 302252 16574 302280 38490
rect 302896 22914 302924 124306
rect 302988 113150 303016 153274
rect 303068 150612 303120 150618
rect 303068 150554 303120 150560
rect 302976 113144 303028 113150
rect 302976 113086 303028 113092
rect 303080 110430 303108 150554
rect 304276 122806 304304 161570
rect 304356 132660 304408 132666
rect 304356 132602 304408 132608
rect 304264 122800 304316 122806
rect 304264 122742 304316 122748
rect 304264 117360 304316 117366
rect 304264 117302 304316 117308
rect 303068 110424 303120 110430
rect 303068 110366 303120 110372
rect 302976 109200 303028 109206
rect 302976 109142 303028 109148
rect 302988 31142 303016 109142
rect 303068 107704 303120 107710
rect 303068 107646 303120 107652
rect 303080 37942 303108 107646
rect 303620 77308 303672 77314
rect 303620 77250 303672 77256
rect 303068 37936 303120 37942
rect 303068 37878 303120 37884
rect 302976 31136 303028 31142
rect 302976 31078 303028 31084
rect 302884 22908 302936 22914
rect 302884 22850 302936 22856
rect 303632 16574 303660 77250
rect 304276 24138 304304 117302
rect 304368 54670 304396 132602
rect 304448 120284 304500 120290
rect 304448 120226 304500 120232
rect 304460 73914 304488 120226
rect 304920 94858 304948 236535
rect 305656 227050 305684 238575
rect 308232 237454 308260 240040
rect 310118 239850 310146 240040
rect 312050 239850 312078 240040
rect 309152 239822 310146 239850
rect 311912 239822 312078 239850
rect 307116 237448 307168 237454
rect 307116 237390 307168 237396
rect 308220 237448 308272 237454
rect 308220 237390 308272 237396
rect 307024 227112 307076 227118
rect 307024 227054 307076 227060
rect 305644 227044 305696 227050
rect 305644 226986 305696 226992
rect 307036 178673 307064 227054
rect 307128 215286 307156 237390
rect 309152 226302 309180 239822
rect 311912 229022 311940 239822
rect 314028 237454 314056 240040
rect 316604 238678 316632 240040
rect 316592 238672 316644 238678
rect 316592 238614 316644 238620
rect 315948 238128 316000 238134
rect 315948 238070 316000 238076
rect 312636 237448 312688 237454
rect 312636 237390 312688 237396
rect 314016 237448 314068 237454
rect 314016 237390 314068 237396
rect 311900 229016 311952 229022
rect 311900 228958 311952 228964
rect 311912 227798 311940 228958
rect 311900 227792 311952 227798
rect 311900 227734 311952 227740
rect 312544 227792 312596 227798
rect 312544 227734 312596 227740
rect 309140 226296 309192 226302
rect 309140 226238 309192 226244
rect 309152 225010 309180 226238
rect 309140 225004 309192 225010
rect 309140 224946 309192 224952
rect 309876 225004 309928 225010
rect 309876 224946 309928 224952
rect 307116 215280 307168 215286
rect 307116 215222 307168 215228
rect 307022 178664 307078 178673
rect 307022 178599 307078 178608
rect 307128 177546 307156 215222
rect 309784 195492 309836 195498
rect 309784 195434 309836 195440
rect 308404 178084 308456 178090
rect 308404 178026 308456 178032
rect 307116 177540 307168 177546
rect 307116 177482 307168 177488
rect 307022 175672 307078 175681
rect 307022 175607 307078 175616
rect 306930 172272 306986 172281
rect 306930 172207 306986 172216
rect 306746 171456 306802 171465
rect 306746 171391 306802 171400
rect 306562 170232 306618 170241
rect 306562 170167 306618 170176
rect 306576 169046 306604 170167
rect 306564 169040 306616 169046
rect 306564 168982 306616 168988
rect 306562 168464 306618 168473
rect 306562 168399 306618 168408
rect 306576 164898 306604 168399
rect 306760 167754 306788 171391
rect 306944 171222 306972 172207
rect 306932 171216 306984 171222
rect 306932 171158 306984 171164
rect 306748 167748 306800 167754
rect 306748 167690 306800 167696
rect 307036 167686 307064 175607
rect 307298 175264 307354 175273
rect 307298 175199 307354 175208
rect 307114 174040 307170 174049
rect 307114 173975 307170 173984
rect 307128 173942 307156 173975
rect 307116 173936 307168 173942
rect 307116 173878 307168 173884
rect 307114 173224 307170 173233
rect 307114 173159 307170 173168
rect 307128 172650 307156 173159
rect 307116 172644 307168 172650
rect 307116 172586 307168 172592
rect 307312 171834 307340 175199
rect 307574 174856 307630 174865
rect 307574 174791 307630 174800
rect 307588 174010 307616 174791
rect 307666 174448 307722 174457
rect 307666 174383 307722 174392
rect 307680 174078 307708 174383
rect 307668 174072 307720 174078
rect 307668 174014 307720 174020
rect 307576 174004 307628 174010
rect 307576 173946 307628 173952
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307588 172718 307616 173567
rect 307576 172712 307628 172718
rect 307576 172654 307628 172660
rect 307666 172680 307722 172689
rect 307666 172615 307722 172624
rect 307680 172582 307708 172615
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 307666 171864 307722 171873
rect 307300 171828 307352 171834
rect 307666 171799 307722 171808
rect 307300 171770 307352 171776
rect 307680 171154 307708 171799
rect 307668 171148 307720 171154
rect 307668 171090 307720 171096
rect 307298 171048 307354 171057
rect 307298 170983 307354 170992
rect 307312 169930 307340 170983
rect 307666 170640 307722 170649
rect 307666 170575 307722 170584
rect 307300 169924 307352 169930
rect 307300 169866 307352 169872
rect 307680 169862 307708 170575
rect 307668 169856 307720 169862
rect 307482 169824 307538 169833
rect 307668 169798 307720 169804
rect 307482 169759 307484 169768
rect 307536 169759 307538 169768
rect 307484 169730 307536 169736
rect 307114 169280 307170 169289
rect 307114 169215 307170 169224
rect 307128 168502 307156 169215
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307116 168496 307168 168502
rect 307116 168438 307168 168444
rect 307680 168434 307708 168807
rect 307668 168428 307720 168434
rect 307668 168370 307720 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307024 167680 307076 167686
rect 307024 167622 307076 167628
rect 307390 167648 307446 167657
rect 307390 167583 307446 167592
rect 307298 167240 307354 167249
rect 307298 167175 307354 167184
rect 307312 166326 307340 167175
rect 307300 166320 307352 166326
rect 307300 166262 307352 166268
rect 306746 165880 306802 165889
rect 306746 165815 306802 165824
rect 306760 165646 306788 165815
rect 306748 165640 306800 165646
rect 306748 165582 306800 165588
rect 307206 165472 307262 165481
rect 307206 165407 307262 165416
rect 307022 165064 307078 165073
rect 307022 164999 307078 165008
rect 306564 164892 306616 164898
rect 306564 164834 306616 164840
rect 306746 163432 306802 163441
rect 306746 163367 306802 163376
rect 305642 162888 305698 162897
rect 305642 162823 305698 162832
rect 305656 124914 305684 162823
rect 306760 162178 306788 163367
rect 306748 162172 306800 162178
rect 306748 162114 306800 162120
rect 306562 160032 306618 160041
rect 306562 159967 306618 159976
rect 306576 158914 306604 159967
rect 306564 158908 306616 158914
rect 306564 158850 306616 158856
rect 306562 158672 306618 158681
rect 306562 158607 306618 158616
rect 306576 157554 306604 158607
rect 306564 157548 306616 157554
rect 306564 157490 306616 157496
rect 306562 156224 306618 156233
rect 306562 156159 306618 156168
rect 306576 156058 306604 156159
rect 306564 156052 306616 156058
rect 306564 155994 306616 156000
rect 306562 154456 306618 154465
rect 306562 154391 306618 154400
rect 306576 153270 306604 154391
rect 306654 153640 306710 153649
rect 306654 153575 306710 153584
rect 306564 153264 306616 153270
rect 306564 153206 306616 153212
rect 306668 151094 306696 153575
rect 306656 151088 306708 151094
rect 306656 151030 306708 151036
rect 306930 151056 306986 151065
rect 306930 150991 306986 151000
rect 306944 150482 306972 150991
rect 306932 150476 306984 150482
rect 306932 150418 306984 150424
rect 306562 150240 306618 150249
rect 306562 150175 306618 150184
rect 306576 149190 306604 150175
rect 306930 149832 306986 149841
rect 306930 149767 306986 149776
rect 306944 149258 306972 149767
rect 306932 149252 306984 149258
rect 306932 149194 306984 149200
rect 306564 149184 306616 149190
rect 306564 149126 306616 149132
rect 306930 147656 306986 147665
rect 306930 147591 306986 147600
rect 306944 145654 306972 147591
rect 306932 145648 306984 145654
rect 306932 145590 306984 145596
rect 306930 145480 306986 145489
rect 306930 145415 306986 145424
rect 306944 144974 306972 145415
rect 306932 144968 306984 144974
rect 306932 144910 306984 144916
rect 306562 144664 306618 144673
rect 306562 144599 306618 144608
rect 306576 143682 306604 144599
rect 306564 143676 306616 143682
rect 306564 143618 306616 143624
rect 306838 141672 306894 141681
rect 306838 141607 306894 141616
rect 306852 133210 306880 141607
rect 307036 141438 307064 164999
rect 307116 164348 307168 164354
rect 307116 164290 307168 164296
rect 307128 164257 307156 164290
rect 307114 164248 307170 164257
rect 307114 164183 307170 164192
rect 307114 152280 307170 152289
rect 307114 152215 307170 152224
rect 307128 142866 307156 152215
rect 307220 145586 307248 165407
rect 307404 163538 307432 167583
rect 307496 167074 307524 167991
rect 307484 167068 307536 167074
rect 307484 167010 307536 167016
rect 307666 166832 307722 166841
rect 307666 166767 307722 166776
rect 307482 166424 307538 166433
rect 307482 166359 307538 166368
rect 307496 163606 307524 166359
rect 307680 165714 307708 166767
rect 307668 165708 307720 165714
rect 307668 165650 307720 165656
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307680 164286 307708 164591
rect 307668 164280 307720 164286
rect 307668 164222 307720 164228
rect 307574 163840 307630 163849
rect 307574 163775 307630 163784
rect 307484 163600 307536 163606
rect 307484 163542 307536 163548
rect 307392 163532 307444 163538
rect 307392 163474 307444 163480
rect 307588 162897 307616 163775
rect 307666 163024 307722 163033
rect 307666 162959 307722 162968
rect 307680 162926 307708 162959
rect 307668 162920 307720 162926
rect 307574 162888 307630 162897
rect 307668 162862 307720 162868
rect 307574 162823 307630 162832
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307496 161634 307524 162415
rect 307574 162072 307630 162081
rect 307574 162007 307630 162016
rect 307484 161628 307536 161634
rect 307484 161570 307536 161576
rect 307588 161566 307616 162007
rect 307666 161664 307722 161673
rect 307666 161599 307722 161608
rect 307576 161560 307628 161566
rect 307576 161502 307628 161508
rect 307680 161498 307708 161599
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307482 161256 307538 161265
rect 307482 161191 307538 161200
rect 307496 160138 307524 161191
rect 307574 160848 307630 160857
rect 307574 160783 307630 160792
rect 307588 160274 307616 160783
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307576 160268 307628 160274
rect 307576 160210 307628 160216
rect 307680 160206 307708 160375
rect 307668 160200 307720 160206
rect 307668 160142 307720 160148
rect 307484 160132 307536 160138
rect 307484 160074 307536 160080
rect 307574 159624 307630 159633
rect 307574 159559 307630 159568
rect 307588 158778 307616 159559
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307680 158846 307708 159015
rect 307668 158840 307720 158846
rect 307668 158782 307720 158788
rect 307576 158772 307628 158778
rect 307576 158714 307628 158720
rect 307666 158264 307722 158273
rect 307666 158199 307722 158208
rect 307482 157856 307538 157865
rect 307482 157791 307538 157800
rect 307390 157448 307446 157457
rect 307496 157418 307524 157791
rect 307680 157486 307708 158199
rect 307668 157480 307720 157486
rect 307668 157422 307720 157428
rect 307390 157383 307446 157392
rect 307484 157412 307536 157418
rect 307404 155242 307432 157383
rect 307484 157354 307536 157360
rect 307666 157040 307722 157049
rect 307666 156975 307722 156984
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307588 155990 307616 156567
rect 307680 156126 307708 156975
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307574 155680 307630 155689
rect 307574 155615 307630 155624
rect 307482 155272 307538 155281
rect 307392 155236 307444 155242
rect 307482 155207 307538 155216
rect 307392 155178 307444 155184
rect 307496 153882 307524 155207
rect 307588 154698 307616 155615
rect 307666 154864 307722 154873
rect 307666 154799 307722 154808
rect 307576 154692 307628 154698
rect 307576 154634 307628 154640
rect 307680 154630 307708 154799
rect 307668 154624 307720 154630
rect 307668 154566 307720 154572
rect 307666 154048 307722 154057
rect 307666 153983 307722 153992
rect 307484 153876 307536 153882
rect 307484 153818 307536 153824
rect 307680 153338 307708 153983
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307666 153232 307722 153241
rect 307666 153167 307722 153176
rect 307680 152522 307708 153167
rect 307668 152516 307720 152522
rect 307668 152458 307720 152464
rect 307666 151872 307722 151881
rect 307666 151807 307668 151816
rect 307720 151807 307722 151816
rect 307668 151778 307720 151784
rect 307298 151464 307354 151473
rect 307298 151399 307354 151408
rect 307312 150550 307340 151399
rect 307666 150648 307722 150657
rect 307666 150583 307668 150592
rect 307720 150583 307722 150592
rect 307668 150554 307720 150560
rect 307300 150544 307352 150550
rect 307300 150486 307352 150492
rect 307298 149288 307354 149297
rect 307298 149223 307354 149232
rect 307312 149122 307340 149223
rect 307300 149116 307352 149122
rect 307300 149058 307352 149064
rect 307482 148880 307538 148889
rect 307482 148815 307538 148824
rect 307496 147830 307524 148815
rect 307574 148472 307630 148481
rect 307574 148407 307630 148416
rect 307484 147824 307536 147830
rect 307484 147766 307536 147772
rect 307588 147762 307616 148407
rect 307666 148064 307722 148073
rect 307666 147999 307722 148008
rect 307576 147756 307628 147762
rect 307576 147698 307628 147704
rect 307680 147694 307708 147999
rect 307668 147688 307720 147694
rect 307668 147630 307720 147636
rect 307482 147248 307538 147257
rect 307482 147183 307538 147192
rect 307496 146334 307524 147183
rect 307574 146840 307630 146849
rect 307574 146775 307630 146784
rect 307588 146470 307616 146775
rect 307576 146464 307628 146470
rect 307576 146406 307628 146412
rect 307666 146432 307722 146441
rect 307666 146367 307668 146376
rect 307720 146367 307722 146376
rect 307668 146338 307720 146344
rect 307484 146328 307536 146334
rect 307484 146270 307536 146276
rect 307482 145888 307538 145897
rect 307482 145823 307538 145832
rect 307208 145580 307260 145586
rect 307208 145522 307260 145528
rect 307390 145072 307446 145081
rect 307390 145007 307446 145016
rect 307298 143848 307354 143857
rect 307298 143783 307354 143792
rect 307116 142860 307168 142866
rect 307116 142802 307168 142808
rect 307206 142488 307262 142497
rect 307206 142423 307262 142432
rect 307024 141432 307076 141438
rect 307024 141374 307076 141380
rect 307114 137456 307170 137465
rect 307114 137391 307170 137400
rect 307022 137048 307078 137057
rect 307022 136983 307078 136992
rect 306930 133240 306986 133249
rect 306840 133204 306892 133210
rect 306930 133175 306986 133184
rect 306840 133146 306892 133152
rect 306944 132666 306972 133175
rect 306932 132660 306984 132666
rect 306932 132602 306984 132608
rect 307036 132494 307064 136983
rect 307128 136678 307156 137391
rect 307116 136672 307168 136678
rect 307116 136614 307168 136620
rect 307114 136232 307170 136241
rect 307114 136167 307170 136176
rect 307128 135522 307156 136167
rect 307116 135516 307168 135522
rect 307116 135458 307168 135464
rect 307036 132466 307156 132494
rect 306562 132288 306618 132297
rect 306562 132223 306618 132232
rect 306576 131238 306604 132223
rect 306564 131232 306616 131238
rect 306564 131174 306616 131180
rect 306562 128072 306618 128081
rect 306562 128007 306618 128016
rect 306576 127090 306604 128007
rect 306564 127084 306616 127090
rect 306564 127026 306616 127032
rect 306562 126848 306618 126857
rect 306562 126783 306618 126792
rect 306576 125662 306604 126783
rect 306564 125656 306616 125662
rect 306564 125598 306616 125604
rect 305644 124908 305696 124914
rect 305644 124850 305696 124856
rect 305826 123312 305882 123321
rect 305826 123247 305882 123256
rect 305734 107808 305790 107817
rect 305734 107743 305790 107752
rect 305642 99648 305698 99657
rect 305642 99583 305698 99592
rect 304908 94852 304960 94858
rect 304908 94794 304960 94800
rect 304448 73908 304500 73914
rect 304448 73850 304500 73856
rect 304356 54664 304408 54670
rect 304356 54606 304408 54612
rect 305000 42152 305052 42158
rect 305000 42094 305052 42100
rect 304264 24132 304316 24138
rect 304264 24074 304316 24080
rect 305012 16574 305040 42094
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301504 13116 301556 13122
rect 301504 13058 301556 13064
rect 301504 7676 301556 7682
rect 301504 7618 301556 7624
rect 301516 6798 301544 7618
rect 301504 6792 301556 6798
rect 301504 6734 301556 6740
rect 299570 3632 299626 3641
rect 299570 3567 299626 3576
rect 300766 3632 300822 3641
rect 300766 3567 300822 3576
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3567
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 6734
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 305656 14482 305684 99583
rect 305748 39370 305776 107743
rect 305840 57390 305868 123247
rect 307022 122088 307078 122097
rect 307022 122023 307078 122032
rect 306746 117872 306802 117881
rect 306746 117807 306802 117816
rect 306760 117570 306788 117807
rect 306748 117564 306800 117570
rect 306748 117506 306800 117512
rect 306748 113280 306800 113286
rect 306746 113248 306748 113257
rect 306800 113248 306802 113257
rect 306746 113183 306802 113192
rect 305918 112024 305974 112033
rect 305918 111959 305974 111968
rect 305932 65618 305960 111959
rect 306746 109848 306802 109857
rect 306746 109783 306802 109792
rect 306760 109206 306788 109783
rect 306748 109200 306800 109206
rect 306748 109142 306800 109148
rect 306930 108896 306986 108905
rect 306930 108831 306986 108840
rect 306944 107710 306972 108831
rect 306932 107704 306984 107710
rect 306932 107646 306984 107652
rect 306746 104272 306802 104281
rect 306746 104207 306802 104216
rect 306760 103698 306788 104207
rect 306748 103692 306800 103698
rect 306748 103634 306800 103640
rect 306746 103048 306802 103057
rect 306746 102983 306802 102992
rect 306760 102338 306788 102983
rect 306748 102332 306800 102338
rect 306748 102274 306800 102280
rect 306930 100872 306986 100881
rect 306930 100807 306986 100816
rect 306944 100774 306972 100807
rect 306932 100768 306984 100774
rect 306932 100710 306984 100716
rect 306746 98696 306802 98705
rect 306746 98631 306802 98640
rect 306760 98054 306788 98631
rect 306748 98048 306800 98054
rect 306748 97990 306800 97996
rect 306930 97880 306986 97889
rect 306930 97815 306986 97824
rect 306944 96762 306972 97815
rect 306932 96756 306984 96762
rect 306932 96698 306984 96704
rect 305920 65612 305972 65618
rect 305920 65554 305972 65560
rect 305828 57384 305880 57390
rect 305828 57326 305880 57332
rect 305736 39364 305788 39370
rect 305736 39306 305788 39312
rect 305644 14476 305696 14482
rect 305644 14418 305696 14424
rect 307036 9042 307064 122023
rect 307128 80714 307156 132466
rect 307220 127634 307248 142423
rect 307312 134570 307340 143783
rect 307404 137290 307432 145007
rect 307496 144226 307524 145823
rect 307666 144256 307722 144265
rect 307484 144220 307536 144226
rect 307666 144191 307722 144200
rect 307484 144162 307536 144168
rect 307680 143614 307708 144191
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 307574 143440 307630 143449
rect 307574 143375 307630 143384
rect 307588 142186 307616 143375
rect 307666 143032 307722 143041
rect 307666 142967 307722 142976
rect 307680 142254 307708 142967
rect 307668 142248 307720 142254
rect 307668 142190 307720 142196
rect 307576 142180 307628 142186
rect 307576 142122 307628 142128
rect 307574 142080 307630 142089
rect 307574 142015 307630 142024
rect 307588 140894 307616 142015
rect 307576 140888 307628 140894
rect 307576 140830 307628 140836
rect 307666 140856 307722 140865
rect 307666 140791 307668 140800
rect 307720 140791 307722 140800
rect 307668 140762 307720 140768
rect 307482 140448 307538 140457
rect 307482 140383 307538 140392
rect 307496 139466 307524 140383
rect 307574 140040 307630 140049
rect 307574 139975 307630 139984
rect 307588 139602 307616 139975
rect 307666 139632 307722 139641
rect 307576 139596 307628 139602
rect 307666 139567 307722 139576
rect 307576 139538 307628 139544
rect 307680 139534 307708 139567
rect 307668 139528 307720 139534
rect 307668 139470 307720 139476
rect 307484 139460 307536 139466
rect 307484 139402 307536 139408
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307574 138136 307630 138145
rect 307680 138106 307708 138207
rect 307574 138071 307630 138080
rect 307668 138100 307720 138106
rect 307588 138038 307616 138071
rect 307668 138042 307720 138048
rect 307576 138032 307628 138038
rect 307576 137974 307628 137980
rect 307666 137864 307722 137873
rect 307666 137799 307722 137808
rect 307392 137284 307444 137290
rect 307392 137226 307444 137232
rect 307680 136746 307708 137799
rect 307668 136740 307720 136746
rect 307668 136682 307720 136688
rect 307482 136640 307538 136649
rect 307482 136575 307538 136584
rect 307496 135318 307524 136575
rect 307574 135688 307630 135697
rect 307574 135623 307630 135632
rect 307588 135386 307616 135623
rect 307668 135448 307720 135454
rect 307668 135390 307720 135396
rect 307576 135380 307628 135386
rect 307576 135322 307628 135328
rect 307484 135312 307536 135318
rect 307680 135289 307708 135390
rect 307484 135254 307536 135260
rect 307666 135280 307722 135289
rect 307666 135215 307722 135224
rect 307574 134872 307630 134881
rect 307574 134807 307630 134816
rect 307300 134564 307352 134570
rect 307300 134506 307352 134512
rect 307588 134026 307616 134807
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307576 134020 307628 134026
rect 307576 133962 307628 133968
rect 307680 133958 307708 134399
rect 307668 133952 307720 133958
rect 307668 133894 307720 133900
rect 307574 133648 307630 133657
rect 307574 133583 307630 133592
rect 307588 132530 307616 133583
rect 307666 132696 307722 132705
rect 307666 132631 307722 132640
rect 307680 132598 307708 132631
rect 307668 132592 307720 132598
rect 307668 132534 307720 132540
rect 307576 132524 307628 132530
rect 307576 132466 307628 132472
rect 307666 131880 307722 131889
rect 307666 131815 307722 131824
rect 307574 131472 307630 131481
rect 307574 131407 307630 131416
rect 307588 131170 307616 131407
rect 307680 131306 307708 131815
rect 307668 131300 307720 131306
rect 307668 131242 307720 131248
rect 307576 131164 307628 131170
rect 307576 131106 307628 131112
rect 307298 131064 307354 131073
rect 307298 130999 307354 131008
rect 307312 129810 307340 130999
rect 307574 130656 307630 130665
rect 307574 130591 307630 130600
rect 307588 129878 307616 130591
rect 307666 130248 307722 130257
rect 307666 130183 307722 130192
rect 307680 129946 307708 130183
rect 307668 129940 307720 129946
rect 307668 129882 307720 129888
rect 307576 129872 307628 129878
rect 307576 129814 307628 129820
rect 307300 129804 307352 129810
rect 307300 129746 307352 129752
rect 307574 128616 307630 128625
rect 307574 128551 307630 128560
rect 307588 128450 307616 128551
rect 307666 128480 307722 128489
rect 307576 128444 307628 128450
rect 307666 128415 307722 128424
rect 307576 128386 307628 128392
rect 307680 128382 307708 128415
rect 307668 128376 307720 128382
rect 307668 128318 307720 128324
rect 307208 127628 307260 127634
rect 307208 127570 307260 127576
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307680 127022 307708 127191
rect 307668 127016 307720 127022
rect 307668 126958 307720 126964
rect 307574 126440 307630 126449
rect 307574 126375 307630 126384
rect 307588 125798 307616 126375
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307576 125792 307628 125798
rect 307576 125734 307628 125740
rect 307680 125730 307708 125831
rect 307668 125724 307720 125730
rect 307668 125666 307720 125672
rect 307298 125488 307354 125497
rect 307298 125423 307354 125432
rect 307206 124264 307262 124273
rect 307312 124234 307340 125423
rect 307574 125080 307630 125089
rect 307574 125015 307630 125024
rect 307588 124302 307616 125015
rect 307666 124672 307722 124681
rect 307666 124607 307722 124616
rect 307680 124370 307708 124607
rect 307668 124364 307720 124370
rect 307668 124306 307720 124312
rect 307576 124296 307628 124302
rect 307576 124238 307628 124244
rect 307206 124199 307262 124208
rect 307300 124228 307352 124234
rect 307116 80708 307168 80714
rect 307116 80650 307168 80656
rect 307220 79354 307248 124199
rect 307300 124170 307352 124176
rect 307574 123856 307630 123865
rect 307574 123791 307630 123800
rect 307588 123010 307616 123791
rect 308416 123457 308444 178026
rect 308494 152688 308550 152697
rect 308494 152623 308550 152632
rect 308402 123448 308458 123457
rect 308402 123383 308458 123392
rect 307666 123040 307722 123049
rect 307576 123004 307628 123010
rect 307666 122975 307722 122984
rect 307576 122946 307628 122952
rect 307680 122942 307708 122975
rect 307668 122936 307720 122942
rect 307668 122878 307720 122884
rect 307574 122496 307630 122505
rect 307574 122431 307630 122440
rect 307588 121582 307616 122431
rect 307666 121680 307722 121689
rect 307666 121615 307722 121624
rect 307576 121576 307628 121582
rect 307576 121518 307628 121524
rect 307680 121514 307708 121615
rect 307668 121508 307720 121514
rect 307668 121450 307720 121456
rect 307482 121272 307538 121281
rect 307482 121207 307538 121216
rect 307496 120154 307524 121207
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120290 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307576 120284 307628 120290
rect 307576 120226 307628 120232
rect 307680 120222 307708 120391
rect 307668 120216 307720 120222
rect 307668 120158 307720 120164
rect 307484 120148 307536 120154
rect 307484 120090 307536 120096
rect 307574 120048 307630 120057
rect 307574 119983 307630 119992
rect 307298 119096 307354 119105
rect 307298 119031 307354 119040
rect 307312 89010 307340 119031
rect 307588 118726 307616 119983
rect 307666 119640 307722 119649
rect 307666 119575 307722 119584
rect 307680 118794 307708 119575
rect 307668 118788 307720 118794
rect 307668 118730 307720 118736
rect 307576 118720 307628 118726
rect 307482 118688 307538 118697
rect 307576 118662 307628 118668
rect 307482 118623 307538 118632
rect 307496 117434 307524 118623
rect 307574 118280 307630 118289
rect 307574 118215 307630 118224
rect 307588 117502 307616 118215
rect 307576 117496 307628 117502
rect 307576 117438 307628 117444
rect 307666 117464 307722 117473
rect 307484 117428 307536 117434
rect 307666 117399 307722 117408
rect 307484 117370 307536 117376
rect 307680 117366 307708 117399
rect 307668 117360 307720 117366
rect 307668 117302 307720 117308
rect 307482 117056 307538 117065
rect 307482 116991 307538 117000
rect 307496 116142 307524 116991
rect 307574 116648 307630 116657
rect 307574 116583 307630 116592
rect 307484 116136 307536 116142
rect 307484 116078 307536 116084
rect 307588 116074 307616 116583
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307576 116068 307628 116074
rect 307576 116010 307628 116016
rect 307680 116006 307708 116175
rect 307668 116000 307720 116006
rect 307668 115942 307720 115948
rect 307574 115696 307630 115705
rect 307574 115631 307630 115640
rect 307588 114646 307616 115631
rect 307666 115288 307722 115297
rect 307666 115223 307722 115232
rect 307576 114640 307628 114646
rect 307576 114582 307628 114588
rect 307680 114578 307708 115223
rect 307668 114572 307720 114578
rect 307668 114514 307720 114520
rect 307574 114064 307630 114073
rect 307574 113999 307630 114008
rect 307588 113218 307616 113999
rect 307666 113656 307722 113665
rect 307666 113591 307722 113600
rect 307680 113354 307708 113591
rect 307668 113348 307720 113354
rect 307668 113290 307720 113296
rect 307576 113212 307628 113218
rect 307576 113154 307628 113160
rect 307574 112704 307630 112713
rect 307574 112639 307630 112648
rect 307588 111926 307616 112639
rect 307576 111920 307628 111926
rect 307576 111862 307628 111868
rect 307666 111888 307722 111897
rect 307666 111823 307668 111832
rect 307720 111823 307722 111832
rect 307668 111794 307720 111800
rect 308508 111790 308536 152623
rect 309690 138680 309746 138689
rect 309690 138615 309746 138624
rect 309704 138145 309732 138615
rect 309690 138136 309746 138145
rect 309690 138071 309746 138080
rect 308496 111784 308548 111790
rect 308496 111726 308548 111732
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110634 307524 111415
rect 307574 111072 307630 111081
rect 307574 111007 307630 111016
rect 307484 110628 307536 110634
rect 307484 110570 307536 110576
rect 307588 110566 307616 111007
rect 307666 110664 307722 110673
rect 307666 110599 307722 110608
rect 307576 110560 307628 110566
rect 307576 110502 307628 110508
rect 307680 110498 307708 110599
rect 307668 110492 307720 110498
rect 307668 110434 307720 110440
rect 307574 110256 307630 110265
rect 307574 110191 307630 110200
rect 307588 109138 307616 110191
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307574 108488 307630 108497
rect 307574 108423 307630 108432
rect 307484 107908 307536 107914
rect 307484 107850 307536 107856
rect 307496 107681 307524 107850
rect 307588 107817 307616 108423
rect 307666 108080 307722 108089
rect 307666 108015 307722 108024
rect 307574 107808 307630 107817
rect 307680 107778 307708 108015
rect 307574 107743 307630 107752
rect 307668 107772 307720 107778
rect 307668 107714 307720 107720
rect 307482 107672 307538 107681
rect 307482 107607 307538 107616
rect 307574 107264 307630 107273
rect 307574 107199 307630 107208
rect 307482 106856 307538 106865
rect 307482 106791 307538 106800
rect 307496 106418 307524 106791
rect 307588 106486 307616 107199
rect 307576 106480 307628 106486
rect 307576 106422 307628 106428
rect 307666 106448 307722 106457
rect 307484 106412 307536 106418
rect 307666 106383 307722 106392
rect 307484 106354 307536 106360
rect 307680 106350 307708 106383
rect 307668 106344 307720 106350
rect 307668 106286 307720 106292
rect 307482 105904 307538 105913
rect 307482 105839 307538 105848
rect 307496 105058 307524 105839
rect 307574 105496 307630 105505
rect 307574 105431 307630 105440
rect 307484 105052 307536 105058
rect 307484 104994 307536 105000
rect 307588 104990 307616 105431
rect 307666 105088 307722 105097
rect 307666 105023 307722 105032
rect 307576 104984 307628 104990
rect 307576 104926 307628 104932
rect 307680 104922 307708 105023
rect 307668 104916 307720 104922
rect 307668 104858 307720 104864
rect 307574 104680 307630 104689
rect 307574 104615 307630 104624
rect 307588 103630 307616 104615
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307576 103624 307628 103630
rect 307576 103566 307628 103572
rect 307680 103562 307708 103799
rect 307668 103556 307720 103562
rect 307668 103498 307720 103504
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307588 102202 307616 103391
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307680 102270 307708 102439
rect 307668 102264 307720 102270
rect 307668 102206 307720 102212
rect 307576 102196 307628 102202
rect 307576 102138 307628 102144
rect 307574 102096 307630 102105
rect 307574 102031 307630 102040
rect 307588 100910 307616 102031
rect 307666 101008 307722 101017
rect 307666 100943 307722 100952
rect 307576 100904 307628 100910
rect 307576 100846 307628 100852
rect 307680 100842 307708 100943
rect 307668 100836 307720 100842
rect 307668 100778 307720 100784
rect 307574 100464 307630 100473
rect 307574 100399 307630 100408
rect 307588 99550 307616 100399
rect 307576 99544 307628 99550
rect 307576 99486 307628 99492
rect 307666 99512 307722 99521
rect 307666 99447 307668 99456
rect 307720 99447 307722 99456
rect 307668 99418 307720 99424
rect 307666 99104 307722 99113
rect 307666 99039 307722 99048
rect 307680 98122 307708 99039
rect 307668 98116 307720 98122
rect 307668 98058 307720 98064
rect 307574 97472 307630 97481
rect 307574 97407 307630 97416
rect 307588 96694 307616 97407
rect 308404 97300 308456 97306
rect 308404 97242 308456 97248
rect 307668 96824 307720 96830
rect 307668 96766 307720 96772
rect 307576 96688 307628 96694
rect 307680 96665 307708 96766
rect 307576 96630 307628 96636
rect 307666 96656 307722 96665
rect 307666 96591 307722 96600
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 308416 93838 308444 97242
rect 309796 96490 309824 195434
rect 309888 180266 309916 224946
rect 309876 180260 309928 180266
rect 309876 180202 309928 180208
rect 312556 178906 312584 227734
rect 312648 216646 312676 237390
rect 315960 229906 315988 238070
rect 316604 238066 316632 238614
rect 316592 238060 316644 238066
rect 316592 238002 316644 238008
rect 318536 237454 318564 240094
rect 319364 238754 319392 244287
rect 319272 238726 319392 238754
rect 318064 237448 318116 237454
rect 318064 237390 318116 237396
rect 318524 237448 318576 237454
rect 318524 237390 318576 237396
rect 316684 236020 316736 236026
rect 316684 235962 316736 235968
rect 315948 229900 316000 229906
rect 315948 229842 316000 229848
rect 315960 229158 315988 229842
rect 315948 229152 316000 229158
rect 315948 229094 316000 229100
rect 312636 216640 312688 216646
rect 312636 216582 312688 216588
rect 312544 178900 312596 178906
rect 312544 178842 312596 178848
rect 312648 177614 312676 216582
rect 313924 201000 313976 201006
rect 313924 200942 313976 200948
rect 312636 177608 312688 177614
rect 312636 177550 312688 177556
rect 313936 175681 313964 200942
rect 314016 195424 314068 195430
rect 314016 195366 314068 195372
rect 314028 177682 314056 195366
rect 316696 180794 316724 235962
rect 316776 229152 316828 229158
rect 316776 229094 316828 229100
rect 316420 180766 316724 180794
rect 316420 178090 316448 180766
rect 316040 178084 316092 178090
rect 316040 178026 316092 178032
rect 316408 178084 316460 178090
rect 316408 178026 316460 178032
rect 314016 177676 314068 177682
rect 314016 177618 314068 177624
rect 316052 175930 316080 178026
rect 316788 177313 316816 229094
rect 318076 229090 318104 237390
rect 319272 231810 319300 238726
rect 319260 231804 319312 231810
rect 319260 231746 319312 231752
rect 318064 229084 318116 229090
rect 318064 229026 318116 229032
rect 318064 226364 318116 226370
rect 318064 226306 318116 226312
rect 316774 177304 316830 177313
rect 316774 177239 316830 177248
rect 318076 176050 318104 226306
rect 318156 223644 318208 223650
rect 318156 223586 318208 223592
rect 318168 176118 318196 223586
rect 319456 177449 319484 360334
rect 319548 307737 319576 375974
rect 320088 374196 320140 374202
rect 320088 374138 320140 374144
rect 320100 373994 320128 374138
rect 320836 373994 320864 683130
rect 327080 401668 327132 401674
rect 327080 401610 327132 401616
rect 324320 392012 324372 392018
rect 324320 391954 324372 391960
rect 323124 378208 323176 378214
rect 323124 378150 323176 378156
rect 320100 373966 320864 373994
rect 320100 361729 320128 373966
rect 321744 372700 321796 372706
rect 321744 372642 321796 372648
rect 321652 367124 321704 367130
rect 321652 367066 321704 367072
rect 320180 366104 320232 366110
rect 320180 366046 320232 366052
rect 320086 361720 320142 361729
rect 320086 361655 320142 361664
rect 319628 359508 319680 359514
rect 319628 359450 319680 359456
rect 319640 347070 319668 359450
rect 319628 347064 319680 347070
rect 319628 347006 319680 347012
rect 319534 307728 319590 307737
rect 319534 307663 319590 307672
rect 319534 298208 319590 298217
rect 319534 298143 319590 298152
rect 319548 297430 319576 298143
rect 319536 297424 319588 297430
rect 319536 297366 319588 297372
rect 319548 239494 319576 297366
rect 320086 240000 320142 240009
rect 320086 239935 320142 239944
rect 319536 239488 319588 239494
rect 319536 239430 319588 239436
rect 320100 239426 320128 239935
rect 320088 239420 320140 239426
rect 320088 239362 320140 239368
rect 320192 238134 320220 366046
rect 320824 361820 320876 361826
rect 320824 361762 320876 361768
rect 320364 358828 320416 358834
rect 320364 358770 320416 358776
rect 320270 356960 320326 356969
rect 320270 356895 320326 356904
rect 320180 238128 320232 238134
rect 320180 238070 320232 238076
rect 320284 236026 320312 356895
rect 320376 325009 320404 358770
rect 320836 348430 320864 361762
rect 321560 358964 321612 358970
rect 321560 358906 321612 358912
rect 320824 348424 320876 348430
rect 320824 348366 320876 348372
rect 321572 331809 321600 358906
rect 321664 347585 321692 367066
rect 321756 359009 321784 372642
rect 322112 363044 322164 363050
rect 322112 362986 322164 362992
rect 321742 359000 321798 359009
rect 321742 358935 321798 358944
rect 322124 354674 322152 362986
rect 323032 360460 323084 360466
rect 323032 360402 323084 360408
rect 322202 359000 322258 359009
rect 322202 358935 322258 358944
rect 322216 358057 322244 358935
rect 322202 358048 322258 358057
rect 322202 357983 322258 357992
rect 322124 354646 322244 354674
rect 322110 352200 322166 352209
rect 322110 352135 322166 352144
rect 322124 351218 322152 352135
rect 322112 351212 322164 351218
rect 322112 351154 322164 351160
rect 321650 347576 321706 347585
rect 321650 347511 321706 347520
rect 321664 344350 321692 347511
rect 322216 345014 322244 354646
rect 322754 350160 322810 350169
rect 322754 350095 322810 350104
rect 322768 349858 322796 350095
rect 322756 349852 322808 349858
rect 322756 349794 322808 349800
rect 322480 345704 322532 345710
rect 322480 345646 322532 345652
rect 322492 345545 322520 345646
rect 322478 345536 322534 345545
rect 322478 345471 322534 345480
rect 322216 344986 322428 345014
rect 321652 344344 321704 344350
rect 321652 344286 321704 344292
rect 322400 339522 322428 344986
rect 322478 343360 322534 343369
rect 322478 343295 322534 343304
rect 322492 342922 322520 343295
rect 322480 342916 322532 342922
rect 322480 342858 322532 342864
rect 322572 341556 322624 341562
rect 322572 341498 322624 341504
rect 322848 341556 322900 341562
rect 322848 341498 322900 341504
rect 322584 341465 322612 341498
rect 322570 341456 322626 341465
rect 322570 341391 322626 341400
rect 322388 339516 322440 339522
rect 322388 339458 322440 339464
rect 322400 338745 322428 339458
rect 322386 338736 322442 338745
rect 322386 338671 322442 338680
rect 322478 336560 322534 336569
rect 322478 336495 322534 336504
rect 322492 336054 322520 336495
rect 322480 336048 322532 336054
rect 322480 335990 322532 335996
rect 322478 334656 322534 334665
rect 322478 334591 322480 334600
rect 322532 334591 322534 334600
rect 322480 334562 322532 334568
rect 321558 331800 321614 331809
rect 321558 331735 321614 331744
rect 322202 331800 322258 331809
rect 322202 331735 322204 331744
rect 322256 331735 322258 331744
rect 322204 331706 322256 331712
rect 322756 331084 322808 331090
rect 322756 331026 322808 331032
rect 322768 329905 322796 331026
rect 322754 329896 322810 329905
rect 322754 329831 322810 329840
rect 322756 327752 322808 327758
rect 322754 327720 322756 327729
rect 322808 327720 322810 327729
rect 322754 327655 322810 327664
rect 322860 326398 322888 341498
rect 322848 326392 322900 326398
rect 322848 326334 322900 326340
rect 320362 325000 320418 325009
rect 320362 324935 320418 324944
rect 320376 324358 320404 324935
rect 320364 324352 320416 324358
rect 320364 324294 320416 324300
rect 322848 324352 322900 324358
rect 322848 324294 322900 324300
rect 322480 322992 322532 322998
rect 322478 322960 322480 322969
rect 322532 322960 322534 322969
rect 322478 322895 322534 322904
rect 322860 322810 322888 324294
rect 322860 322782 322980 322810
rect 322846 320920 322902 320929
rect 322846 320855 322902 320864
rect 322860 320210 322888 320855
rect 322848 320204 322900 320210
rect 322848 320146 322900 320152
rect 322480 317416 322532 317422
rect 322480 317358 322532 317364
rect 322492 316305 322520 317358
rect 322478 316296 322534 316305
rect 322478 316231 322534 316240
rect 322480 314628 322532 314634
rect 322480 314570 322532 314576
rect 322492 314265 322520 314570
rect 322478 314256 322534 314265
rect 322478 314191 322534 314200
rect 322848 312588 322900 312594
rect 322848 312530 322900 312536
rect 322860 312225 322888 312530
rect 322846 312216 322902 312225
rect 322846 312151 322902 312160
rect 322480 309800 322532 309806
rect 322480 309742 322532 309748
rect 322492 309505 322520 309742
rect 322478 309496 322534 309505
rect 322478 309431 322534 309440
rect 321742 307728 321798 307737
rect 321742 307663 321798 307672
rect 321756 307086 321784 307663
rect 321744 307080 321796 307086
rect 321744 307022 321796 307028
rect 322478 305280 322534 305289
rect 322478 305215 322534 305224
rect 322492 305046 322520 305215
rect 322480 305040 322532 305046
rect 322480 304982 322532 304988
rect 322478 303240 322534 303249
rect 322478 303175 322534 303184
rect 322492 302258 322520 303175
rect 322480 302252 322532 302258
rect 322480 302194 322532 302200
rect 322570 300520 322626 300529
rect 322570 300455 322626 300464
rect 322584 300150 322612 300455
rect 322572 300144 322624 300150
rect 322572 300086 322624 300092
rect 322756 300144 322808 300150
rect 322756 300086 322808 300092
rect 322478 296440 322534 296449
rect 322478 296375 322534 296384
rect 322492 295390 322520 296375
rect 322480 295384 322532 295390
rect 322480 295326 322532 295332
rect 322768 294642 322796 300086
rect 322756 294636 322808 294642
rect 322756 294578 322808 294584
rect 322846 293720 322902 293729
rect 322846 293655 322902 293664
rect 322860 293282 322888 293655
rect 322848 293276 322900 293282
rect 322848 293218 322900 293224
rect 322478 291680 322534 291689
rect 322478 291615 322534 291624
rect 322492 291242 322520 291615
rect 322480 291236 322532 291242
rect 322480 291178 322532 291184
rect 321558 289640 321614 289649
rect 321558 289575 321614 289584
rect 320824 276072 320876 276078
rect 320824 276014 320876 276020
rect 320362 242856 320418 242865
rect 320362 242791 320418 242800
rect 320272 236020 320324 236026
rect 320272 235962 320324 235968
rect 320376 230489 320404 242791
rect 320836 239873 320864 276014
rect 321468 242956 321520 242962
rect 321468 242898 321520 242904
rect 321480 242865 321508 242898
rect 321466 242856 321522 242865
rect 321466 242791 321522 242800
rect 320822 239864 320878 239873
rect 320822 239799 320878 239808
rect 321572 234546 321600 289575
rect 322756 287700 322808 287706
rect 322756 287642 322808 287648
rect 322478 286920 322534 286929
rect 322478 286855 322534 286864
rect 322492 285734 322520 286855
rect 322480 285728 322532 285734
rect 322480 285670 322532 285676
rect 322768 285025 322796 287642
rect 322754 285016 322810 285025
rect 322754 284951 322810 284960
rect 322478 282976 322534 282985
rect 322478 282911 322480 282920
rect 322532 282911 322534 282920
rect 322480 282882 322532 282888
rect 322478 280800 322534 280809
rect 322478 280735 322534 280744
rect 322492 280226 322520 280735
rect 322480 280220 322532 280226
rect 322480 280162 322532 280168
rect 321834 278080 321890 278089
rect 321834 278015 321890 278024
rect 321848 276690 321876 278015
rect 321836 276684 321888 276690
rect 321836 276626 321888 276632
rect 321848 276078 321876 276626
rect 321836 276072 321888 276078
rect 321836 276014 321888 276020
rect 322202 276040 322258 276049
rect 322202 275975 322258 275984
rect 321650 271280 321706 271289
rect 321650 271215 321706 271224
rect 321480 234530 321600 234546
rect 321468 234524 321600 234530
rect 321520 234518 321600 234524
rect 321468 234466 321520 234472
rect 321560 234456 321612 234462
rect 321560 234398 321612 234404
rect 321572 233918 321600 234398
rect 321560 233912 321612 233918
rect 321560 233854 321612 233860
rect 320362 230480 320418 230489
rect 320362 230415 320418 230424
rect 321664 224874 321692 271215
rect 321834 255640 321890 255649
rect 321834 255575 321890 255584
rect 321742 244760 321798 244769
rect 321742 244695 321798 244704
rect 321756 244322 321784 244695
rect 321744 244316 321796 244322
rect 321744 244258 321796 244264
rect 321744 239420 321796 239426
rect 321744 239362 321796 239368
rect 321652 224868 321704 224874
rect 321652 224810 321704 224816
rect 321664 224505 321692 224810
rect 321650 224496 321706 224505
rect 321650 224431 321706 224440
rect 319536 211200 319588 211206
rect 319536 211142 319588 211148
rect 319442 177440 319498 177449
rect 319442 177375 319498 177384
rect 319548 176662 319576 211142
rect 321560 202428 321612 202434
rect 321560 202370 321612 202376
rect 321284 178832 321336 178838
rect 321284 178774 321336 178780
rect 319536 176656 319588 176662
rect 319536 176598 319588 176604
rect 318156 176112 318208 176118
rect 318156 176054 318208 176060
rect 318064 176044 318116 176050
rect 318064 175986 318116 175992
rect 316020 175902 316080 175930
rect 313922 175672 313978 175681
rect 313922 175607 313978 175616
rect 321296 172689 321324 178774
rect 321374 175808 321430 175817
rect 321374 175743 321430 175752
rect 321388 173777 321416 175743
rect 321374 173768 321430 173777
rect 321374 173703 321430 173712
rect 321282 172680 321338 172689
rect 321282 172615 321338 172624
rect 321572 132705 321600 202370
rect 321652 194132 321704 194138
rect 321652 194074 321704 194080
rect 321558 132696 321614 132705
rect 321558 132631 321614 132640
rect 321664 129713 321692 194074
rect 321756 162217 321784 239362
rect 321848 234462 321876 255575
rect 322216 241466 322244 275975
rect 322388 274644 322440 274650
rect 322388 274586 322440 274592
rect 322400 274145 322428 274586
rect 322386 274136 322442 274145
rect 322386 274071 322442 274080
rect 322846 269240 322902 269249
rect 322846 269175 322902 269184
rect 322860 269142 322888 269175
rect 322848 269136 322900 269142
rect 322848 269078 322900 269084
rect 322480 267708 322532 267714
rect 322480 267650 322532 267656
rect 322492 267345 322520 267650
rect 322478 267336 322534 267345
rect 322478 267271 322534 267280
rect 322478 265160 322534 265169
rect 322478 265095 322534 265104
rect 322492 264994 322520 265095
rect 322480 264988 322532 264994
rect 322480 264930 322532 264936
rect 322478 262440 322534 262449
rect 322478 262375 322534 262384
rect 322492 262274 322520 262375
rect 322480 262268 322532 262274
rect 322480 262210 322532 262216
rect 322478 260400 322534 260409
rect 322478 260335 322534 260344
rect 322492 259486 322520 260335
rect 322480 259480 322532 259486
rect 322480 259422 322532 259428
rect 322846 258360 322902 258369
rect 322846 258295 322902 258304
rect 322860 258194 322888 258295
rect 322848 258188 322900 258194
rect 322848 258130 322900 258136
rect 322846 253600 322902 253609
rect 322846 253535 322902 253544
rect 322860 252618 322888 253535
rect 322848 252612 322900 252618
rect 322848 252554 322900 252560
rect 322478 248840 322534 248849
rect 322478 248775 322534 248784
rect 322492 248470 322520 248775
rect 322480 248464 322532 248470
rect 322480 248406 322532 248412
rect 322478 246800 322534 246809
rect 322478 246735 322534 246744
rect 322492 245682 322520 246735
rect 322480 245676 322532 245682
rect 322480 245618 322532 245624
rect 322204 241460 322256 241466
rect 322204 241402 322256 241408
rect 322204 234524 322256 234530
rect 322204 234466 322256 234472
rect 321836 234456 321888 234462
rect 321836 234398 321888 234404
rect 321742 162208 321798 162217
rect 321742 162143 321798 162152
rect 322216 158681 322244 234466
rect 322952 174729 322980 322782
rect 322938 174720 322994 174729
rect 322938 174655 322994 174664
rect 323044 160857 323072 360402
rect 323136 354385 323164 378150
rect 323216 369980 323268 369986
rect 323216 369922 323268 369928
rect 323122 354376 323178 354385
rect 323122 354311 323178 354320
rect 323228 349858 323256 369922
rect 323308 363248 323360 363254
rect 323308 363190 323360 363196
rect 323216 349852 323268 349858
rect 323216 349794 323268 349800
rect 323124 177336 323176 177342
rect 323124 177278 323176 177284
rect 323136 163169 323164 177278
rect 323122 163160 323178 163169
rect 323122 163095 323178 163104
rect 323030 160848 323086 160857
rect 323030 160783 323086 160792
rect 322202 158672 322258 158681
rect 322202 158607 322258 158616
rect 323320 135561 323348 363190
rect 324332 331242 324360 391954
rect 324504 371408 324556 371414
rect 324504 371350 324556 371356
rect 324412 364540 324464 364546
rect 324412 364482 324464 364488
rect 324240 331214 324360 331242
rect 324240 330970 324268 331214
rect 324318 331120 324374 331129
rect 324318 331055 324320 331064
rect 324372 331055 324374 331064
rect 324320 331026 324372 331032
rect 324240 330942 324360 330970
rect 324332 327758 324360 330942
rect 324320 327752 324372 327758
rect 324320 327694 324372 327700
rect 324320 320204 324372 320210
rect 324320 320146 324372 320152
rect 323582 251560 323638 251569
rect 323582 251495 323638 251504
rect 323596 220862 323624 251495
rect 324332 235249 324360 320146
rect 324424 293282 324452 364482
rect 324516 312594 324544 371350
rect 325792 367328 325844 367334
rect 325792 367270 325844 367276
rect 325698 363080 325754 363089
rect 325698 363015 325754 363024
rect 324596 358896 324648 358902
rect 324596 358838 324648 358844
rect 324608 331129 324636 358838
rect 324594 331120 324650 331129
rect 324594 331055 324650 331064
rect 324504 312588 324556 312594
rect 324504 312530 324556 312536
rect 325712 309806 325740 363015
rect 325804 334626 325832 367270
rect 327092 345710 327120 401610
rect 328550 386472 328606 386481
rect 328550 386407 328606 386416
rect 327172 374128 327224 374134
rect 327172 374070 327224 374076
rect 327080 345704 327132 345710
rect 327080 345646 327132 345652
rect 327184 342922 327212 374070
rect 328460 344344 328512 344350
rect 328460 344286 328512 344292
rect 327172 342916 327224 342922
rect 327172 342858 327224 342864
rect 325792 334620 325844 334626
rect 325792 334562 325844 334568
rect 327448 331764 327500 331770
rect 327448 331706 327500 331712
rect 325700 309800 325752 309806
rect 325700 309742 325752 309748
rect 327172 305040 327224 305046
rect 327172 304982 327224 304988
rect 325700 302252 325752 302258
rect 325700 302194 325752 302200
rect 324412 293276 324464 293282
rect 324412 293218 324464 293224
rect 324504 258188 324556 258194
rect 324504 258130 324556 258136
rect 324412 252612 324464 252618
rect 324412 252554 324464 252560
rect 324318 235240 324374 235249
rect 324318 235175 324374 235184
rect 324424 227633 324452 252554
rect 324516 237289 324544 258130
rect 324596 241460 324648 241466
rect 324596 241402 324648 241408
rect 324608 240174 324636 241402
rect 324596 240168 324648 240174
rect 324596 240110 324648 240116
rect 324502 237280 324558 237289
rect 324502 237215 324558 237224
rect 324608 234569 324636 240110
rect 324688 235340 324740 235346
rect 324688 235282 324740 235288
rect 324594 234560 324650 234569
rect 324594 234495 324650 234504
rect 324410 227624 324466 227633
rect 324410 227559 324466 227568
rect 323584 220856 323636 220862
rect 323584 220798 323636 220804
rect 324504 217456 324556 217462
rect 324504 217398 324556 217404
rect 324412 175976 324464 175982
rect 324412 175918 324464 175924
rect 324320 172508 324372 172514
rect 324320 172450 324372 172456
rect 324332 171737 324360 172450
rect 324318 171728 324374 171737
rect 324318 171663 324374 171672
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170921 324360 171022
rect 324318 170912 324374 170921
rect 324318 170847 324374 170856
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 169425 324360 169662
rect 324318 169416 324374 169425
rect 324318 169351 324374 169360
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167793 324360 168302
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324320 165572 324372 165578
rect 324320 165514 324372 165520
rect 324332 165481 324360 165514
rect 324318 165472 324374 165481
rect 324318 165407 324374 165416
rect 324320 164212 324372 164218
rect 324320 164154 324372 164160
rect 324332 163985 324360 164154
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 162489 324360 162794
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324320 160268 324372 160274
rect 324320 160210 324372 160216
rect 324332 160177 324360 160210
rect 324318 160168 324374 160177
rect 324318 160103 324374 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324320 158704 324372 158710
rect 324320 158646 324372 158652
rect 324332 157865 324360 158646
rect 324318 157856 324374 157865
rect 324318 157791 324374 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 157049 324360 157286
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324424 156369 324452 175918
rect 324516 174049 324544 217398
rect 324502 174040 324558 174049
rect 324502 173975 324558 173984
rect 324504 169652 324556 169658
rect 324504 169594 324556 169600
rect 324516 168609 324544 169594
rect 324502 168600 324558 168609
rect 324502 168535 324558 168544
rect 324504 168292 324556 168298
rect 324504 168234 324556 168240
rect 324516 167113 324544 168234
rect 324502 167104 324558 167113
rect 324502 167039 324558 167048
rect 324504 165504 324556 165510
rect 324504 165446 324556 165452
rect 324516 164801 324544 165446
rect 324502 164792 324558 164801
rect 324502 164727 324558 164736
rect 324410 156360 324466 156369
rect 324410 156295 324466 156304
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 155553 324360 155858
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324412 154488 324464 154494
rect 324412 154430 324464 154436
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324424 153241 324452 154430
rect 324410 153232 324466 153241
rect 324320 153196 324372 153202
rect 324410 153167 324466 153176
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 324320 151768 324372 151774
rect 324320 151710 324372 151716
rect 324332 150929 324360 151710
rect 324318 150920 324374 150929
rect 324318 150855 324374 150864
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150340 324464 150346
rect 324412 150282 324464 150288
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150282
rect 324502 149696 324558 149705
rect 324502 149631 324558 149640
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324412 149048 324464 149054
rect 324412 148990 324464 148996
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 324332 148617 324360 148922
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324424 147801 324452 148990
rect 324410 147792 324466 147801
rect 324410 147727 324466 147736
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324374 146240
rect 324412 146260 324464 146266
rect 324332 146198 324360 146231
rect 324412 146202 324464 146208
rect 324320 146192 324372 146198
rect 324320 146134 324372 146140
rect 324424 145489 324452 146202
rect 324410 145480 324466 145489
rect 324410 145415 324466 145424
rect 324320 143540 324372 143546
rect 324320 143482 324372 143488
rect 324332 143177 324360 143482
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324516 142497 324544 149631
rect 324502 142488 324558 142497
rect 324502 142423 324558 142432
rect 324412 142112 324464 142118
rect 324412 142054 324464 142060
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324424 140865 324452 142054
rect 324410 140856 324466 140865
rect 324410 140791 324466 140800
rect 324320 139120 324372 139126
rect 324320 139062 324372 139068
rect 324332 138553 324360 139062
rect 324318 138544 324374 138553
rect 324318 138479 324374 138488
rect 324412 137964 324464 137970
rect 324412 137906 324464 137912
rect 324320 137896 324372 137902
rect 324318 137864 324320 137873
rect 324372 137864 324374 137873
rect 324318 137799 324374 137808
rect 324424 137057 324452 137906
rect 324410 137048 324466 137057
rect 324410 136983 324466 136992
rect 324320 136604 324372 136610
rect 324320 136546 324372 136552
rect 324332 136377 324360 136546
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 323306 135552 323362 135561
rect 323306 135487 323362 135496
rect 324320 135176 324372 135182
rect 324320 135118 324372 135124
rect 324332 134745 324360 135118
rect 324412 135108 324464 135114
rect 324412 135050 324464 135056
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324424 134065 324452 135050
rect 324410 134056 324466 134065
rect 324410 133991 324466 134000
rect 324320 133612 324372 133618
rect 324320 133554 324372 133560
rect 324332 133249 324360 133554
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130121 324360 131038
rect 324318 130112 324374 130121
rect 324318 130047 324374 130056
rect 324320 129736 324372 129742
rect 321650 129704 321706 129713
rect 324320 129678 324372 129684
rect 321650 129639 321706 129648
rect 324332 128625 324360 129678
rect 324318 128616 324374 128625
rect 324318 128551 324374 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324412 128240 324464 128246
rect 324412 128182 324464 128188
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 128182
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 125497 324360 125530
rect 324412 125520 324464 125526
rect 324318 125488 324374 125497
rect 324412 125462 324464 125468
rect 324318 125423 324374 125432
rect 324424 124817 324452 125462
rect 324410 124808 324466 124817
rect 324410 124743 324466 124752
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 124001 324360 124102
rect 324412 124092 324464 124098
rect 324412 124034 324464 124040
rect 324318 123992 324374 124001
rect 324318 123927 324374 123936
rect 324424 123185 324452 124034
rect 324410 123176 324466 123185
rect 324410 123111 324466 123120
rect 324412 122800 324464 122806
rect 324412 122742 324464 122748
rect 324320 122732 324372 122738
rect 324320 122674 324372 122680
rect 324332 122505 324360 122674
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 324424 121689 324452 122742
rect 324410 121680 324466 121689
rect 324410 121615 324466 121624
rect 324412 121440 324464 121446
rect 324412 121382 324464 121388
rect 324320 121372 324372 121378
rect 324320 121314 324372 121320
rect 324332 120873 324360 121314
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121382
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324412 117292 324464 117298
rect 324412 117234 324464 117240
rect 324320 117224 324372 117230
rect 324320 117166 324372 117172
rect 324332 117065 324360 117166
rect 324318 117056 324374 117065
rect 324318 116991 324374 117000
rect 324424 116385 324452 117234
rect 324410 116376 324466 116385
rect 324410 116311 324466 116320
rect 324320 115932 324372 115938
rect 324320 115874 324372 115880
rect 324332 115569 324360 115874
rect 324412 115864 324464 115870
rect 324412 115806 324464 115812
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324424 114753 324452 115806
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324320 114504 324372 114510
rect 324320 114446 324372 114452
rect 324332 114073 324360 114446
rect 324412 114436 324464 114442
rect 324412 114378 324464 114384
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114378
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 322940 112464 322992 112470
rect 324332 112441 324360 113086
rect 322940 112406 322992 112412
rect 324318 112432 324374 112441
rect 321834 110528 321890 110537
rect 321834 110463 321890 110472
rect 321650 102776 321706 102785
rect 321650 102711 321706 102720
rect 321558 99648 321614 99657
rect 321558 99583 321614 99592
rect 321374 98832 321430 98841
rect 321374 98767 321430 98776
rect 309784 96484 309836 96490
rect 309784 96426 309836 96432
rect 321388 95198 321416 98767
rect 321466 96656 321522 96665
rect 321466 96591 321468 96600
rect 321520 96591 321522 96600
rect 321468 96562 321520 96568
rect 321572 96558 321600 99583
rect 321560 96552 321612 96558
rect 321560 96494 321612 96500
rect 321664 96490 321692 102711
rect 321742 102232 321798 102241
rect 321742 102167 321798 102176
rect 321652 96484 321704 96490
rect 321652 96426 321704 96432
rect 321376 95192 321428 95198
rect 321376 95134 321428 95140
rect 321756 95062 321784 102167
rect 321848 95130 321876 110463
rect 321836 95124 321888 95130
rect 321836 95066 321888 95072
rect 321744 95056 321796 95062
rect 321744 94998 321796 95004
rect 308404 93832 308456 93838
rect 308404 93774 308456 93780
rect 320824 93220 320876 93226
rect 320824 93162 320876 93168
rect 313280 91792 313332 91798
rect 313280 91734 313332 91740
rect 307300 89004 307352 89010
rect 307300 88946 307352 88952
rect 311900 86284 311952 86290
rect 311900 86226 311952 86232
rect 307208 79348 307260 79354
rect 307208 79290 307260 79296
rect 309784 79348 309836 79354
rect 309784 79290 309836 79296
rect 308402 59936 308458 59945
rect 308402 59871 308458 59880
rect 308416 9654 308444 59871
rect 308494 40624 308550 40633
rect 308494 40559 308550 40568
rect 308404 9648 308456 9654
rect 308404 9590 308456 9596
rect 307024 9036 307076 9042
rect 307024 8978 307076 8984
rect 306748 7608 306800 7614
rect 306748 7550 306800 7556
rect 306760 480 306788 7550
rect 308508 6730 308536 40559
rect 309048 9648 309100 9654
rect 309048 9590 309100 9596
rect 308496 6724 308548 6730
rect 308496 6666 308548 6672
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 354 308026 480
rect 308508 354 308536 6666
rect 309060 480 309088 9590
rect 309796 6730 309824 79290
rect 309876 75200 309928 75206
rect 309876 75142 309928 75148
rect 309888 40730 309916 75142
rect 311164 49700 311216 49706
rect 311164 49642 311216 49648
rect 311176 49094 311204 49642
rect 311164 49088 311216 49094
rect 311164 49030 311216 49036
rect 309876 40724 309928 40730
rect 309876 40666 309928 40672
rect 309784 6724 309836 6730
rect 309784 6666 309836 6672
rect 307914 326 308536 354
rect 307914 -960 308026 326
rect 309018 -960 309130 480
rect 309888 354 309916 40666
rect 311176 16574 311204 49030
rect 311912 16574 311940 86226
rect 312544 75200 312596 75206
rect 312544 75142 312596 75148
rect 312556 49706 312584 75142
rect 312544 49700 312596 49706
rect 312544 49642 312596 49648
rect 313292 38554 313320 91734
rect 316040 89004 316092 89010
rect 316040 88946 316092 88952
rect 315304 83496 315356 83502
rect 315304 83438 315356 83444
rect 313924 42084 313976 42090
rect 313924 42026 313976 42032
rect 313280 38548 313332 38554
rect 313280 38490 313332 38496
rect 313292 38010 313320 38490
rect 313280 38004 313332 38010
rect 313280 37946 313332 37952
rect 313936 33114 313964 42026
rect 313924 33108 313976 33114
rect 313924 33050 313976 33056
rect 313936 32094 313964 33050
rect 313280 32088 313332 32094
rect 313280 32030 313332 32036
rect 313924 32088 313976 32094
rect 313924 32030 313976 32036
rect 313292 16574 313320 32030
rect 311176 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309888 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 13802 315344 83438
rect 316052 16574 316080 88946
rect 318800 87712 318852 87718
rect 318800 87654 318852 87660
rect 317420 80708 317472 80714
rect 317420 80650 317472 80656
rect 316682 43480 316738 43489
rect 316682 43415 316738 43424
rect 317326 43480 317382 43489
rect 317326 43415 317328 43424
rect 316052 16546 316264 16574
rect 314660 13796 314712 13802
rect 314660 13738 314712 13744
rect 315304 13796 315356 13802
rect 315304 13738 315356 13744
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 13738
rect 316236 480 316264 16546
rect 316696 3534 316724 43415
rect 317380 43415 317382 43424
rect 317328 43386 317380 43392
rect 317432 16574 317460 80650
rect 318812 16574 318840 87654
rect 320180 45552 320232 45558
rect 320180 45494 320232 45500
rect 320192 45286 320220 45494
rect 320836 45286 320864 93162
rect 321560 90364 321612 90370
rect 321560 90306 321612 90312
rect 320180 45280 320232 45286
rect 320180 45222 320232 45228
rect 320824 45280 320876 45286
rect 320824 45222 320876 45228
rect 320192 16574 320220 45222
rect 321572 16574 321600 90306
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316684 3528 316736 3534
rect 316684 3470 316736 3476
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 317340 480 317368 3470
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 112406
rect 324318 112367 324374 112376
rect 323030 111752 323086 111761
rect 323030 111687 323086 111696
rect 323044 94994 323072 111687
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 109449 324360 110366
rect 324412 109744 324464 109750
rect 324412 109686 324464 109692
rect 324318 109440 324374 109449
rect 324318 109375 324374 109384
rect 324320 108792 324372 108798
rect 324320 108734 324372 108740
rect 324332 107817 324360 108734
rect 324318 107808 324374 107817
rect 324318 107743 324374 107752
rect 324320 107636 324372 107642
rect 324320 107578 324372 107584
rect 324332 107137 324360 107578
rect 324318 107128 324374 107137
rect 324318 107063 324374 107072
rect 323122 106312 323178 106321
rect 323122 106247 323178 106256
rect 323032 94988 323084 94994
rect 323032 94930 323084 94936
rect 323136 93770 323164 106247
rect 323214 105496 323270 105505
rect 323214 105431 323270 105440
rect 323228 94926 323256 105431
rect 324424 104825 324452 109686
rect 324700 108633 324728 235282
rect 325712 230314 325740 302194
rect 327184 238754 327212 304982
rect 327264 269136 327316 269142
rect 327264 269078 327316 269084
rect 327092 238726 327212 238754
rect 327092 233238 327120 238726
rect 327276 234598 327304 269078
rect 327356 259480 327408 259486
rect 327356 259422 327408 259428
rect 327264 234592 327316 234598
rect 327264 234534 327316 234540
rect 327080 233232 327132 233238
rect 327080 233174 327132 233180
rect 327368 230450 327396 259422
rect 327356 230444 327408 230450
rect 327356 230386 327408 230392
rect 325700 230308 325752 230314
rect 325700 230250 325752 230256
rect 325712 229094 325740 230250
rect 325712 229066 325832 229094
rect 325700 207800 325752 207806
rect 325700 207742 325752 207748
rect 324964 169788 325016 169794
rect 324964 169730 325016 169736
rect 324976 151745 325004 169730
rect 324962 151736 325018 151745
rect 324962 151671 325018 151680
rect 324686 108624 324742 108633
rect 324686 108559 324742 108568
rect 324410 104816 324466 104825
rect 324410 104751 324466 104760
rect 325606 104000 325662 104009
rect 325712 103986 325740 207742
rect 325804 143993 325832 229066
rect 327172 196784 327224 196790
rect 327172 196726 327224 196732
rect 325976 195356 326028 195362
rect 325976 195298 326028 195304
rect 325884 180260 325936 180266
rect 325884 180202 325936 180208
rect 325790 143984 325846 143993
rect 325790 143919 325846 143928
rect 325896 119377 325924 180202
rect 325988 139126 326016 195298
rect 327080 176656 327132 176662
rect 327080 176598 327132 176604
rect 327092 169794 327120 176598
rect 327080 169788 327132 169794
rect 327080 169730 327132 169736
rect 325976 139120 326028 139126
rect 325976 139062 326028 139068
rect 325882 119368 325938 119377
rect 325882 119303 325938 119312
rect 327184 108798 327212 196726
rect 327264 178900 327316 178906
rect 327264 178842 327316 178848
rect 327276 133618 327304 178842
rect 327460 160274 327488 331706
rect 328368 234592 328420 234598
rect 328368 234534 328420 234540
rect 328380 233986 328408 234534
rect 328368 233980 328420 233986
rect 328368 233922 328420 233928
rect 328368 233232 328420 233238
rect 328368 233174 328420 233180
rect 328380 232626 328408 233174
rect 328368 232620 328420 232626
rect 328368 232562 328420 232568
rect 328368 230444 328420 230450
rect 328368 230386 328420 230392
rect 328380 229906 328408 230386
rect 328368 229900 328420 229906
rect 328368 229842 328420 229848
rect 327448 160268 327500 160274
rect 327448 160210 327500 160216
rect 328472 146198 328500 344286
rect 328564 342242 328592 386407
rect 334636 372774 334664 696934
rect 356704 577516 356756 577522
rect 356704 577458 356756 577464
rect 342260 405748 342312 405754
rect 342260 405690 342312 405696
rect 335450 390688 335506 390697
rect 335450 390623 335506 390632
rect 333980 372768 334032 372774
rect 333980 372710 334032 372716
rect 334624 372768 334676 372774
rect 334624 372710 334676 372716
rect 331312 365900 331364 365906
rect 331312 365842 331364 365848
rect 328552 342236 328604 342242
rect 328552 342178 328604 342184
rect 328564 341562 328592 342178
rect 328552 341556 328604 341562
rect 328552 341498 328604 341504
rect 329840 334620 329892 334626
rect 329840 334562 329892 334568
rect 328552 282940 328604 282946
rect 328552 282882 328604 282888
rect 328564 237250 328592 282882
rect 328552 237244 328604 237250
rect 328552 237186 328604 237192
rect 328460 146192 328512 146198
rect 328460 146134 328512 146140
rect 328564 142050 328592 237186
rect 328736 192772 328788 192778
rect 328736 192714 328788 192720
rect 328644 176112 328696 176118
rect 328644 176054 328696 176060
rect 328552 142044 328604 142050
rect 328552 141986 328604 141992
rect 327264 133612 327316 133618
rect 327264 133554 327316 133560
rect 328656 121378 328684 176054
rect 328748 154494 328776 192714
rect 328736 154488 328788 154494
rect 328736 154430 328788 154436
rect 328644 121372 328696 121378
rect 328644 121314 328696 121320
rect 329852 109750 329880 334562
rect 331220 322992 331272 322998
rect 331220 322934 331272 322940
rect 329932 285728 329984 285734
rect 329932 285670 329984 285676
rect 329944 235958 329972 285670
rect 330024 264988 330076 264994
rect 330024 264930 330076 264936
rect 329932 235952 329984 235958
rect 329932 235894 329984 235900
rect 329944 148986 329972 235894
rect 330036 226166 330064 264930
rect 331232 238754 331260 322934
rect 331324 314634 331352 365842
rect 332876 339516 332928 339522
rect 332876 339458 332928 339464
rect 331312 314628 331364 314634
rect 331312 314570 331364 314576
rect 331324 313954 331352 314570
rect 331312 313948 331364 313954
rect 331312 313890 331364 313896
rect 331312 295384 331364 295390
rect 331312 295326 331364 295332
rect 331324 248414 331352 295326
rect 331324 248386 331628 248414
rect 331232 238726 331352 238754
rect 331324 237318 331352 238726
rect 331600 238542 331628 248386
rect 332692 245676 332744 245682
rect 332692 245618 332744 245624
rect 331588 238536 331640 238542
rect 331588 238478 331640 238484
rect 331312 237312 331364 237318
rect 331312 237254 331364 237260
rect 330024 226160 330076 226166
rect 330024 226102 330076 226108
rect 330036 153202 330064 226102
rect 330116 184272 330168 184278
rect 330116 184214 330168 184220
rect 330024 153196 330076 153202
rect 330024 153138 330076 153144
rect 329932 148980 329984 148986
rect 329932 148922 329984 148928
rect 330128 128246 330156 184214
rect 331324 155922 331352 237254
rect 331404 191208 331456 191214
rect 331404 191150 331456 191156
rect 331416 165510 331444 191150
rect 331496 176044 331548 176050
rect 331496 175986 331548 175992
rect 331404 165504 331456 165510
rect 331404 165446 331456 165452
rect 331508 160070 331536 175986
rect 331496 160064 331548 160070
rect 331496 160006 331548 160012
rect 331312 155916 331364 155922
rect 331312 155858 331364 155864
rect 330116 128240 330168 128246
rect 330116 128182 330168 128188
rect 329840 109744 329892 109750
rect 329840 109686 329892 109692
rect 327172 108792 327224 108798
rect 327172 108734 327224 108740
rect 325662 103958 325740 103986
rect 325606 103935 325662 103944
rect 330484 102808 330536 102814
rect 330484 102750 330536 102756
rect 324502 101688 324558 101697
rect 324502 101623 324558 101632
rect 324412 98660 324464 98666
rect 324412 98602 324464 98608
rect 324320 97980 324372 97986
rect 324320 97922 324372 97928
rect 324332 97073 324360 97922
rect 324424 97889 324452 98602
rect 324410 97880 324466 97889
rect 324410 97815 324466 97824
rect 324318 97064 324374 97073
rect 324318 96999 324374 97008
rect 323216 94920 323268 94926
rect 323216 94862 323268 94868
rect 324516 94858 324544 101623
rect 324594 100872 324650 100881
rect 324594 100807 324650 100816
rect 324504 94852 324556 94858
rect 324504 94794 324556 94800
rect 323124 93764 323176 93770
rect 323124 93706 323176 93712
rect 324608 92478 324636 100807
rect 325700 100020 325752 100026
rect 325700 99962 325752 99968
rect 324596 92472 324648 92478
rect 324596 92414 324648 92420
rect 324320 82136 324372 82142
rect 324318 82104 324320 82113
rect 324372 82104 324374 82113
rect 324318 82039 324374 82048
rect 324332 3534 324360 82039
rect 325712 16574 325740 99962
rect 327724 47592 327776 47598
rect 327724 47534 327776 47540
rect 327736 33114 327764 47534
rect 327724 33108 327776 33114
rect 327724 33050 327776 33056
rect 327736 31822 327764 33050
rect 327080 31816 327132 31822
rect 327080 31758 327132 31764
rect 327724 31816 327776 31822
rect 327724 31758 327776 31764
rect 327092 16574 327120 31758
rect 330496 27606 330524 102750
rect 331600 98666 331628 238478
rect 332704 220726 332732 245618
rect 332692 220720 332744 220726
rect 332692 220662 332744 220668
rect 332690 185600 332746 185609
rect 332690 185535 332746 185544
rect 332600 177404 332652 177410
rect 332600 177346 332652 177352
rect 332612 169658 332640 177346
rect 332600 169652 332652 169658
rect 332600 169594 332652 169600
rect 331864 157412 331916 157418
rect 331864 157354 331916 157360
rect 331588 98660 331640 98666
rect 331588 98602 331640 98608
rect 331312 70576 331364 70582
rect 331312 70518 331364 70524
rect 329840 27600 329892 27606
rect 329840 27542 329892 27548
rect 330484 27600 330536 27606
rect 330484 27542 330536 27548
rect 329852 16574 329880 27542
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 324412 3460 324464 3466
rect 324412 3402 324464 3408
rect 324424 480 324452 3402
rect 325620 480 325648 3470
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 329196 3528 329248 3534
rect 329196 3470 329248 3476
rect 329208 480 329236 3470
rect 330404 480 330432 16546
rect 331324 3534 331352 70518
rect 331876 41410 331904 157354
rect 332704 143546 332732 185535
rect 332784 177676 332836 177682
rect 332784 177618 332836 177624
rect 332796 164218 332824 177618
rect 332784 164212 332836 164218
rect 332784 164154 332836 164160
rect 332692 143540 332744 143546
rect 332692 143482 332744 143488
rect 332888 110430 332916 339458
rect 333992 336054 334020 372710
rect 335360 368620 335412 368626
rect 335360 368562 335412 368568
rect 333980 336048 334032 336054
rect 333980 335990 334032 335996
rect 333992 333266 334020 335990
rect 333980 333260 334032 333266
rect 333980 333202 334032 333208
rect 335372 267714 335400 368562
rect 335464 317422 335492 390623
rect 340880 374264 340932 374270
rect 340880 374206 340932 374212
rect 339500 372632 339552 372638
rect 339500 372574 339552 372580
rect 338764 371272 338816 371278
rect 338764 371214 338816 371220
rect 337384 370524 337436 370530
rect 337384 370466 337436 370472
rect 335452 317416 335504 317422
rect 335452 317358 335504 317364
rect 336648 317416 336700 317422
rect 336648 317358 336700 317364
rect 336660 316742 336688 317358
rect 336648 316736 336700 316742
rect 336648 316678 336700 316684
rect 336004 280220 336056 280226
rect 336004 280162 336056 280168
rect 336016 273290 336044 280162
rect 336004 273284 336056 273290
rect 336004 273226 336056 273232
rect 335360 267708 335412 267714
rect 335360 267650 335412 267656
rect 334348 262880 334400 262886
rect 334348 262822 334400 262828
rect 334360 262274 334388 262822
rect 334072 262268 334124 262274
rect 334072 262210 334124 262216
rect 334348 262268 334400 262274
rect 334348 262210 334400 262216
rect 333980 233912 334032 233918
rect 333980 233854 334032 233860
rect 333992 150346 334020 233854
rect 334084 231742 334112 262210
rect 335452 248464 335504 248470
rect 335452 248406 335504 248412
rect 335360 233980 335412 233986
rect 335360 233922 335412 233928
rect 334072 231736 334124 231742
rect 334072 231678 334124 231684
rect 334072 188420 334124 188426
rect 334072 188362 334124 188368
rect 333980 150340 334032 150346
rect 333980 150282 334032 150288
rect 333244 142860 333296 142866
rect 333244 142802 333296 142808
rect 332876 110424 332928 110430
rect 332876 110366 332928 110372
rect 333256 89010 333284 142802
rect 334084 117298 334112 188362
rect 334164 177540 334216 177546
rect 334164 177482 334216 177488
rect 334176 129742 334204 177482
rect 334256 177472 334308 177478
rect 334256 177414 334308 177420
rect 334268 167006 334296 177414
rect 334256 167000 334308 167006
rect 334256 166942 334308 166948
rect 334624 164280 334676 164286
rect 334624 164222 334676 164228
rect 334164 129736 334216 129742
rect 334164 129678 334216 129684
rect 334072 117292 334124 117298
rect 334072 117234 334124 117240
rect 333980 94512 334032 94518
rect 333980 94454 334032 94460
rect 333992 91050 334020 94454
rect 333980 91044 334032 91050
rect 333980 90986 334032 90992
rect 333244 89004 333296 89010
rect 333244 88946 333296 88952
rect 331954 86184 332010 86193
rect 331954 86119 332010 86128
rect 331864 41404 331916 41410
rect 331864 41346 331916 41352
rect 331968 12434 331996 86119
rect 332048 83496 332100 83502
rect 332048 83438 332100 83444
rect 332060 71670 332088 83438
rect 332048 71664 332100 71670
rect 332048 71606 332100 71612
rect 332060 70582 332088 71606
rect 333244 71120 333296 71126
rect 333244 71062 333296 71068
rect 332048 70576 332100 70582
rect 332048 70518 332100 70524
rect 333256 70446 333284 71062
rect 333244 70440 333296 70446
rect 333244 70382 333296 70388
rect 332600 58676 332652 58682
rect 332600 58618 332652 58624
rect 332612 57798 332640 58618
rect 332600 57792 332652 57798
rect 332600 57734 332652 57740
rect 331600 12406 331996 12434
rect 331600 9654 331628 12406
rect 331588 9648 331640 9654
rect 331588 9590 331640 9596
rect 331312 3528 331364 3534
rect 331312 3470 331364 3476
rect 331600 480 331628 9590
rect 332612 8906 332640 57734
rect 332600 8900 332652 8906
rect 332600 8842 332652 8848
rect 333256 4146 333284 70382
rect 333992 16574 334020 90986
rect 334636 78130 334664 164222
rect 335372 113150 335400 233922
rect 335464 219434 335492 248406
rect 335452 219428 335504 219434
rect 335452 219370 335504 219376
rect 336016 218006 336044 273226
rect 336648 267708 336700 267714
rect 336648 267650 336700 267656
rect 336660 267034 336688 267650
rect 336648 267028 336700 267034
rect 336648 266970 336700 266976
rect 336740 229900 336792 229906
rect 336740 229842 336792 229848
rect 336004 218000 336056 218006
rect 336004 217942 336056 217948
rect 335544 191276 335596 191282
rect 335544 191218 335596 191224
rect 335452 180192 335504 180198
rect 335452 180134 335504 180140
rect 335464 150414 335492 180134
rect 335556 165578 335584 191218
rect 335636 189916 335688 189922
rect 335636 189858 335688 189864
rect 335648 169726 335676 189858
rect 335636 169720 335688 169726
rect 335636 169662 335688 169668
rect 335544 165572 335596 165578
rect 335544 165514 335596 165520
rect 336004 155984 336056 155990
rect 336004 155926 336056 155932
rect 335452 150408 335504 150414
rect 335452 150350 335504 150356
rect 335360 113144 335412 113150
rect 335360 113086 335412 113092
rect 334716 89004 334768 89010
rect 334716 88946 334768 88952
rect 334624 78124 334676 78130
rect 334624 78066 334676 78072
rect 334728 70446 334756 88946
rect 336016 76634 336044 155926
rect 336752 115870 336780 229842
rect 336830 177304 336886 177313
rect 336830 177239 336886 177248
rect 336740 115864 336792 115870
rect 336740 115806 336792 115812
rect 336844 114442 336872 177239
rect 336922 175264 336978 175273
rect 336922 175199 336978 175208
rect 336936 158710 336964 175199
rect 336924 158704 336976 158710
rect 336924 158646 336976 158652
rect 336832 114436 336884 114442
rect 336832 114378 336884 114384
rect 336096 84856 336148 84862
rect 336096 84798 336148 84804
rect 336004 76628 336056 76634
rect 336004 76570 336056 76576
rect 334716 70440 334768 70446
rect 334716 70382 334768 70388
rect 336108 69018 336136 84798
rect 335360 69012 335412 69018
rect 335360 68954 335412 68960
rect 336096 69012 336148 69018
rect 336096 68954 336148 68960
rect 335372 16574 335400 68954
rect 337396 16574 337424 370466
rect 338120 199504 338172 199510
rect 338120 199446 338172 199452
rect 338132 137902 338160 199446
rect 338212 181620 338264 181626
rect 338212 181562 338264 181568
rect 338120 137896 338172 137902
rect 338120 137838 338172 137844
rect 338224 128314 338252 181562
rect 338302 177440 338358 177449
rect 338302 177375 338358 177384
rect 338316 157350 338344 177375
rect 338776 174554 338804 371214
rect 339512 274650 339540 372574
rect 340144 291236 340196 291242
rect 340144 291178 340196 291184
rect 340156 288454 340184 291178
rect 340144 288448 340196 288454
rect 340144 288390 340196 288396
rect 339500 274644 339552 274650
rect 339500 274586 339552 274592
rect 339512 273970 339540 274586
rect 339500 273964 339552 273970
rect 339500 273906 339552 273912
rect 340156 227662 340184 288390
rect 340236 229832 340288 229838
rect 340236 229774 340288 229780
rect 340144 227656 340196 227662
rect 340144 227598 340196 227604
rect 339592 185700 339644 185706
rect 339592 185642 339644 185648
rect 339500 177608 339552 177614
rect 339500 177550 339552 177556
rect 338764 174548 338816 174554
rect 338764 174490 338816 174496
rect 338764 168428 338816 168434
rect 338764 168370 338816 168376
rect 338304 157344 338356 157350
rect 338304 157286 338356 157292
rect 338212 128308 338264 128314
rect 338212 128250 338264 128256
rect 338776 66978 338804 168370
rect 339512 115938 339540 177550
rect 339604 151774 339632 185642
rect 340144 176724 340196 176730
rect 340144 176666 340196 176672
rect 339592 151768 339644 151774
rect 339592 151710 339644 151716
rect 339500 115932 339552 115938
rect 339500 115874 339552 115880
rect 339408 78668 339460 78674
rect 339408 78610 339460 78616
rect 339420 78577 339448 78610
rect 339406 78568 339462 78577
rect 339406 78503 339462 78512
rect 339420 77314 339448 78503
rect 339408 77308 339460 77314
rect 339408 77250 339460 77256
rect 338856 73840 338908 73846
rect 338856 73782 338908 73788
rect 338764 66972 338816 66978
rect 338764 66914 338816 66920
rect 338868 45490 338896 73782
rect 339500 73228 339552 73234
rect 339500 73170 339552 73176
rect 338856 45484 338908 45490
rect 338856 45426 338908 45432
rect 338868 44198 338896 45426
rect 338120 44192 338172 44198
rect 338120 44134 338172 44140
rect 338856 44192 338908 44198
rect 338856 44134 338908 44140
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 333888 8900 333940 8906
rect 333888 8842 333940 8848
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 332704 480 332732 4082
rect 333900 480 333928 8842
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 337028 16546 337424 16574
rect 338132 16574 338160 44134
rect 338132 16546 338712 16574
rect 337028 15201 337056 16546
rect 337014 15192 337070 15201
rect 337014 15127 337070 15136
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 15127
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 73170
rect 340156 13190 340184 176666
rect 340248 135250 340276 229774
rect 340236 135244 340288 135250
rect 340236 135186 340288 135192
rect 340892 107642 340920 374206
rect 341524 211948 341576 211954
rect 341524 211890 341576 211896
rect 340972 184340 341024 184346
rect 340972 184282 341024 184288
rect 340984 114510 341012 184282
rect 341064 183116 341116 183122
rect 341064 183058 341116 183064
rect 341076 154562 341104 183058
rect 341064 154556 341116 154562
rect 341064 154498 341116 154504
rect 340972 114504 341024 114510
rect 340972 114446 341024 114452
rect 340880 107636 340932 107642
rect 340880 107578 340932 107584
rect 341536 106282 341564 211890
rect 342272 143546 342300 405690
rect 353300 403640 353352 403646
rect 353300 403582 353352 403588
rect 351920 400920 351972 400926
rect 351920 400862 351972 400868
rect 349804 381540 349856 381546
rect 349804 381482 349856 381488
rect 347780 378276 347832 378282
rect 347780 378218 347832 378224
rect 345020 367396 345072 367402
rect 345020 367338 345072 367344
rect 342352 364676 342404 364682
rect 342352 364618 342404 364624
rect 342364 162858 342392 364618
rect 343640 364608 343692 364614
rect 343640 364550 343692 364556
rect 342904 227044 342956 227050
rect 342904 226986 342956 226992
rect 342444 185904 342496 185910
rect 342444 185846 342496 185852
rect 342352 162852 342404 162858
rect 342352 162794 342404 162800
rect 342456 149054 342484 185846
rect 342444 149048 342496 149054
rect 342444 148990 342496 148996
rect 342350 144800 342406 144809
rect 342350 144735 342406 144744
rect 342364 143614 342392 144735
rect 342352 143608 342404 143614
rect 342352 143550 342404 143556
rect 342260 143540 342312 143546
rect 342260 143482 342312 143488
rect 342272 142866 342300 143482
rect 342260 142860 342312 142866
rect 342260 142802 342312 142808
rect 341524 106276 341576 106282
rect 341524 106218 341576 106224
rect 342260 86352 342312 86358
rect 342260 86294 342312 86300
rect 340880 46232 340932 46238
rect 340878 46200 340880 46209
rect 340932 46200 340934 46209
rect 340878 46135 340934 46144
rect 342272 16574 342300 86294
rect 342364 86290 342392 143550
rect 342916 117298 342944 226986
rect 343652 125526 343680 364550
rect 343824 192636 343876 192642
rect 343824 192578 343876 192584
rect 343730 183016 343786 183025
rect 343730 182951 343786 182960
rect 343640 125520 343692 125526
rect 343640 125462 343692 125468
rect 342904 117292 342956 117298
rect 342904 117234 342956 117240
rect 342352 86284 342404 86290
rect 342352 86226 342404 86232
rect 343744 74526 343772 182951
rect 343836 118590 343864 192578
rect 343916 182844 343968 182850
rect 343916 182786 343968 182792
rect 343928 124098 343956 182786
rect 345032 168298 345060 367338
rect 346400 365832 346452 365838
rect 346400 365774 346452 365780
rect 345112 232620 345164 232626
rect 345112 232562 345164 232568
rect 345020 168292 345072 168298
rect 345020 168234 345072 168240
rect 343916 124092 343968 124098
rect 343916 124034 343968 124040
rect 343824 118584 343876 118590
rect 343824 118526 343876 118532
rect 345124 117230 345152 232562
rect 345204 189780 345256 189786
rect 345204 189722 345256 189728
rect 345216 118658 345244 189722
rect 345296 182912 345348 182918
rect 345296 182854 345348 182860
rect 345308 122738 345336 182854
rect 345664 161492 345716 161498
rect 345664 161434 345716 161440
rect 345296 122732 345348 122738
rect 345296 122674 345348 122680
rect 345204 118652 345256 118658
rect 345204 118594 345256 118600
rect 345112 117224 345164 117230
rect 345112 117166 345164 117172
rect 343732 74520 343784 74526
rect 343732 74462 343784 74468
rect 343744 73234 343772 74462
rect 343732 73228 343784 73234
rect 343732 73170 343784 73176
rect 345676 47734 345704 161434
rect 346412 97986 346440 365774
rect 346492 218068 346544 218074
rect 346492 218010 346544 218016
rect 346504 137970 346532 218010
rect 347042 182880 347098 182889
rect 347042 182815 347098 182824
rect 346582 180024 346638 180033
rect 346582 179959 346638 179968
rect 346492 137964 346544 137970
rect 346492 137906 346544 137912
rect 346596 135114 346624 179959
rect 346584 135108 346636 135114
rect 346584 135050 346636 135056
rect 346400 97980 346452 97986
rect 346400 97922 346452 97928
rect 345756 71800 345808 71806
rect 345756 71742 345808 71748
rect 345664 47728 345716 47734
rect 345664 47670 345716 47676
rect 345020 47592 345072 47598
rect 345020 47534 345072 47540
rect 343640 44872 343692 44878
rect 343640 44814 343692 44820
rect 343652 16574 343680 44814
rect 345032 16574 345060 47534
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 340144 13184 340196 13190
rect 340144 13126 340196 13132
rect 342166 11792 342222 11801
rect 342166 11727 342222 11736
rect 340970 7576 341026 7585
rect 340970 7511 341026 7520
rect 340984 480 341012 7511
rect 342180 480 342208 11727
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 345768 3466 345796 71742
rect 347056 6914 347084 182815
rect 347792 168366 347820 378218
rect 349160 366036 349212 366042
rect 349160 365978 349212 365984
rect 347872 222216 347924 222222
rect 347872 222158 347924 222164
rect 347780 168360 347832 168366
rect 347780 168302 347832 168308
rect 347884 122806 347912 222158
rect 347964 220856 348016 220862
rect 347964 220798 348016 220804
rect 347976 125594 348004 220798
rect 348424 174548 348476 174554
rect 348424 174490 348476 174496
rect 347964 125588 348016 125594
rect 347964 125530 348016 125536
rect 347872 122800 347924 122806
rect 347872 122742 347924 122748
rect 346964 6886 347084 6914
rect 346964 4146 346992 6886
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 345756 3460 345808 3466
rect 345756 3402 345808 3408
rect 346964 480 346992 4082
rect 348436 4049 348464 174490
rect 349172 142118 349200 365978
rect 349252 202292 349304 202298
rect 349252 202234 349304 202240
rect 349160 142112 349212 142118
rect 349160 142054 349212 142060
rect 349264 113150 349292 202234
rect 349344 178764 349396 178770
rect 349344 178706 349396 178712
rect 349356 131102 349384 178706
rect 349344 131096 349396 131102
rect 349344 131038 349396 131044
rect 349252 113144 349304 113150
rect 349252 113086 349304 113092
rect 349264 112470 349292 113086
rect 349252 112464 349304 112470
rect 349252 112406 349304 112412
rect 349816 86290 349844 381482
rect 350540 365968 350592 365974
rect 350540 365910 350592 365916
rect 350552 135182 350580 365910
rect 350632 229764 350684 229770
rect 350632 229706 350684 229712
rect 350644 146266 350672 229706
rect 351184 196716 351236 196722
rect 351184 196658 351236 196664
rect 350632 146260 350684 146266
rect 350632 146202 350684 146208
rect 350540 135176 350592 135182
rect 350540 135118 350592 135124
rect 351196 96626 351224 196658
rect 350540 96620 350592 96626
rect 350540 96562 350592 96568
rect 351184 96620 351236 96626
rect 351184 96562 351236 96568
rect 349804 86284 349856 86290
rect 349804 86226 349856 86232
rect 349160 49020 349212 49026
rect 349160 48962 349212 48968
rect 349172 46918 349200 48962
rect 349160 46912 349212 46918
rect 349160 46854 349212 46860
rect 349172 16574 349200 46854
rect 349172 16546 349292 16574
rect 348422 4040 348478 4049
rect 348422 3975 348478 3984
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 354 348138 480
rect 348436 354 348464 3975
rect 349264 480 349292 16546
rect 349816 3534 349844 86226
rect 350552 16574 350580 96562
rect 351932 81394 351960 400862
rect 352012 368824 352064 368830
rect 352012 368766 352064 368772
rect 352024 147626 352052 368766
rect 352104 187060 352156 187066
rect 352104 187002 352156 187008
rect 352012 147620 352064 147626
rect 352012 147562 352064 147568
rect 351920 81388 351972 81394
rect 351920 81330 351972 81336
rect 351932 80714 351960 81330
rect 351920 80708 351972 80714
rect 351920 80650 351972 80656
rect 352116 73098 352144 187002
rect 352196 182980 352248 182986
rect 352196 182922 352248 182928
rect 352208 136610 352236 182922
rect 353312 142118 353340 403582
rect 353944 378208 353996 378214
rect 353944 378150 353996 378156
rect 353956 297430 353984 378150
rect 354680 371476 354732 371482
rect 354680 371418 354732 371424
rect 353944 297424 353996 297430
rect 353944 297366 353996 297372
rect 353390 222864 353446 222873
rect 353390 222799 353446 222808
rect 353300 142112 353352 142118
rect 353300 142054 353352 142060
rect 353312 140826 353340 142054
rect 352656 140820 352708 140826
rect 352656 140762 352708 140768
rect 353300 140820 353352 140826
rect 353300 140762 353352 140768
rect 352196 136604 352248 136610
rect 352196 136546 352248 136552
rect 352668 87718 352696 140762
rect 353404 93854 353432 222799
rect 354692 171086 354720 371418
rect 356060 363112 356112 363118
rect 356060 363054 356112 363060
rect 354772 193928 354824 193934
rect 354772 193870 354824 193876
rect 354680 171080 354732 171086
rect 354680 171022 354732 171028
rect 353944 165640 353996 165646
rect 353944 165582 353996 165588
rect 353312 93826 353432 93854
rect 352656 87712 352708 87718
rect 352656 87654 352708 87660
rect 352564 87644 352616 87650
rect 352564 87586 352616 87592
rect 352104 73092 352156 73098
rect 352104 73034 352156 73040
rect 352116 71806 352144 73034
rect 352104 71800 352156 71806
rect 352104 71742 352156 71748
rect 350552 16546 351224 16574
rect 349804 3528 349856 3534
rect 349804 3470 349856 3476
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 348026 326 348464 354
rect 348026 -960 348138 326
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352576 4146 352604 87586
rect 353312 86970 353340 93826
rect 353300 86964 353352 86970
rect 353300 86906 353352 86912
rect 353312 86358 353340 86906
rect 353300 86352 353352 86358
rect 353300 86294 353352 86300
rect 353956 49162 353984 165582
rect 353944 49156 353996 49162
rect 353944 49098 353996 49104
rect 354784 8265 354812 193870
rect 356072 121446 356100 363054
rect 356716 300150 356744 577458
rect 357440 378344 357492 378350
rect 357440 378286 357492 378292
rect 356704 300144 356756 300150
rect 356704 300086 356756 300092
rect 356796 154624 356848 154630
rect 356796 154566 356848 154572
rect 356704 146328 356756 146334
rect 356704 146270 356756 146276
rect 356060 121440 356112 121446
rect 356060 121382 356112 121388
rect 356716 9586 356744 146270
rect 356808 46306 356836 154566
rect 357452 124166 357480 378286
rect 358740 287706 358768 702986
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429200 702840 429252 702846
rect 429200 702782 429252 702788
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 425704 702704 425756 702710
rect 425704 702646 425756 702652
rect 425716 700330 425744 702646
rect 425704 700324 425756 700330
rect 425704 700266 425756 700272
rect 385684 590708 385736 590714
rect 385684 590650 385736 590656
rect 370504 418192 370556 418198
rect 370504 418134 370556 418140
rect 360200 392080 360252 392086
rect 360200 392022 360252 392028
rect 358820 376848 358872 376854
rect 358820 376790 358872 376796
rect 358728 287700 358780 287706
rect 358728 287642 358780 287648
rect 358084 173936 358136 173942
rect 358084 173878 358136 173884
rect 357440 124160 357492 124166
rect 357440 124102 357492 124108
rect 356796 46300 356848 46306
rect 356796 46242 356848 46248
rect 358096 12374 358124 173878
rect 358832 172514 358860 376790
rect 359464 360324 359516 360330
rect 359464 360266 359516 360272
rect 358820 172508 358872 172514
rect 358820 172450 358872 172456
rect 359476 104854 359504 360266
rect 359556 150476 359608 150482
rect 359556 150418 359608 150424
rect 359464 104848 359516 104854
rect 359464 104790 359516 104796
rect 359568 19310 359596 150418
rect 360212 100706 360240 392022
rect 360844 351212 360896 351218
rect 360844 351154 360896 351160
rect 360856 324970 360884 351154
rect 370516 342242 370544 418134
rect 385696 395350 385724 590650
rect 385684 395344 385736 395350
rect 385684 395286 385736 395292
rect 403624 375420 403676 375426
rect 403624 375362 403676 375368
rect 385684 367260 385736 367266
rect 385684 367202 385736 367208
rect 370504 342236 370556 342242
rect 370504 342178 370556 342184
rect 371884 333260 371936 333266
rect 371884 333202 371936 333208
rect 360844 324964 360896 324970
rect 360844 324906 360896 324912
rect 361488 300144 361540 300150
rect 361488 300086 361540 300092
rect 361500 263634 361528 300086
rect 370504 293276 370556 293282
rect 370504 293218 370556 293224
rect 360292 263628 360344 263634
rect 360292 263570 360344 263576
rect 361488 263628 361540 263634
rect 361488 263570 361540 263576
rect 360304 262886 360332 263570
rect 360292 262880 360344 262886
rect 360292 262822 360344 262828
rect 370516 260166 370544 293218
rect 370504 260160 370556 260166
rect 370504 260102 370556 260108
rect 362958 221504 363014 221513
rect 362958 221439 363014 221448
rect 360844 153264 360896 153270
rect 360844 153206 360896 153212
rect 360200 100700 360252 100706
rect 360200 100642 360252 100648
rect 360212 100026 360240 100642
rect 360200 100020 360252 100026
rect 360200 99962 360252 99968
rect 360856 32502 360884 153206
rect 362972 45558 363000 221439
rect 367100 217320 367152 217326
rect 367100 217262 367152 217268
rect 363604 149116 363656 149122
rect 363604 149058 363656 149064
rect 362960 45552 363012 45558
rect 362960 45494 363012 45500
rect 362972 44878 363000 45494
rect 362960 44872 363012 44878
rect 362960 44814 363012 44820
rect 360844 32496 360896 32502
rect 360844 32438 360896 32444
rect 359556 19304 359608 19310
rect 359556 19246 359608 19252
rect 358084 12368 358136 12374
rect 358084 12310 358136 12316
rect 356704 9580 356756 9586
rect 356704 9522 356756 9528
rect 354770 8256 354826 8265
rect 354770 8191 354826 8200
rect 354784 7585 354812 8191
rect 354770 7576 354826 7585
rect 354770 7511 354826 7520
rect 363616 6798 363644 149058
rect 367112 47598 367140 217262
rect 369858 148336 369914 148345
rect 369858 148271 369914 148280
rect 369872 147694 369900 148271
rect 369860 147688 369912 147694
rect 369860 147630 369912 147636
rect 367744 139460 367796 139466
rect 367744 139402 367796 139408
rect 367756 113150 367784 139402
rect 367744 113144 367796 113150
rect 367744 113086 367796 113092
rect 367836 48272 367888 48278
rect 367836 48214 367888 48220
rect 367848 47598 367876 48214
rect 367100 47592 367152 47598
rect 367100 47534 367152 47540
rect 367836 47592 367888 47598
rect 367836 47534 367888 47540
rect 369872 42158 369900 147630
rect 370504 136672 370556 136678
rect 370504 136614 370556 136620
rect 370516 100706 370544 136614
rect 371896 111790 371924 333202
rect 380900 324964 380952 324970
rect 380900 324906 380952 324912
rect 380912 324358 380940 324906
rect 380900 324352 380952 324358
rect 380900 324294 380952 324300
rect 382188 324352 382240 324358
rect 382188 324294 382240 324300
rect 377404 309800 377456 309806
rect 377404 309742 377456 309748
rect 374644 245676 374696 245682
rect 374644 245618 374696 245624
rect 374656 133890 374684 245618
rect 376024 135312 376076 135318
rect 376024 135254 376076 135260
rect 374644 133884 374696 133890
rect 374644 133826 374696 133832
rect 371884 111784 371936 111790
rect 371884 111726 371936 111732
rect 376036 102814 376064 135254
rect 377416 110430 377444 309742
rect 378784 244316 378836 244322
rect 378784 244258 378836 244264
rect 377404 110424 377456 110430
rect 377404 110366 377456 110372
rect 376024 102808 376076 102814
rect 376024 102750 376076 102756
rect 378796 100706 378824 244258
rect 382200 122806 382228 324294
rect 382924 273964 382976 273970
rect 382924 273906 382976 273912
rect 382936 128314 382964 273906
rect 385696 180062 385724 367202
rect 389824 360256 389876 360262
rect 389824 360198 389876 360204
rect 388444 297424 388496 297430
rect 388444 297366 388496 297372
rect 385684 180056 385736 180062
rect 385684 179998 385736 180004
rect 386328 180056 386380 180062
rect 386328 179998 386380 180004
rect 386340 179450 386368 179998
rect 386328 179444 386380 179450
rect 386328 179386 386380 179392
rect 386340 133210 386368 179386
rect 386328 133204 386380 133210
rect 386328 133146 386380 133152
rect 382924 128308 382976 128314
rect 382924 128250 382976 128256
rect 382188 122800 382240 122806
rect 382188 122742 382240 122748
rect 388456 121446 388484 297366
rect 388444 121440 388496 121446
rect 388444 121382 388496 121388
rect 370504 100700 370556 100706
rect 370504 100642 370556 100648
rect 378784 100700 378836 100706
rect 378784 100642 378836 100648
rect 389836 95198 389864 360198
rect 395344 312588 395396 312594
rect 395344 312530 395396 312536
rect 393964 258120 394016 258126
rect 393964 258062 394016 258068
rect 393976 185706 394004 258062
rect 393964 185700 394016 185706
rect 393964 185642 394016 185648
rect 395356 113150 395384 312530
rect 400864 204944 400916 204950
rect 400864 204886 400916 204892
rect 399484 203584 399536 203590
rect 399484 203526 399536 203532
rect 396724 202156 396776 202162
rect 396724 202098 396776 202104
rect 395344 113144 395396 113150
rect 395344 113086 395396 113092
rect 396736 96529 396764 202098
rect 399496 97986 399524 203526
rect 400876 99278 400904 204886
rect 403636 181626 403664 375362
rect 417424 371340 417476 371346
rect 417424 371282 417476 371288
rect 413284 363180 413336 363186
rect 413284 363122 413336 363128
rect 406384 362228 406436 362234
rect 406384 362170 406436 362176
rect 403714 192536 403770 192545
rect 403714 192471 403770 192480
rect 403624 181620 403676 181626
rect 403624 181562 403676 181568
rect 403728 107642 403756 192471
rect 403716 107636 403768 107642
rect 403716 107578 403768 107584
rect 406396 100638 406424 362170
rect 410522 359408 410578 359417
rect 410522 359343 410578 359352
rect 407764 213240 407816 213246
rect 407764 213182 407816 213188
rect 407776 103494 407804 213182
rect 410536 181694 410564 359343
rect 410616 193860 410668 193866
rect 410616 193802 410668 193808
rect 410524 181688 410576 181694
rect 410524 181630 410576 181636
rect 407764 103488 407816 103494
rect 407764 103430 407816 103436
rect 406384 100632 406436 100638
rect 406384 100574 406436 100580
rect 400864 99272 400916 99278
rect 400864 99214 400916 99220
rect 410628 99210 410656 193802
rect 411904 192500 411956 192506
rect 411904 192442 411956 192448
rect 411916 132462 411944 192442
rect 411904 132456 411956 132462
rect 411904 132398 411956 132404
rect 410616 99204 410668 99210
rect 410616 99146 410668 99152
rect 399484 97980 399536 97986
rect 399484 97922 399536 97928
rect 413296 97918 413324 363122
rect 414662 360224 414718 360233
rect 414662 360159 414718 360168
rect 414676 182918 414704 360159
rect 417436 271930 417464 371282
rect 420920 294636 420972 294642
rect 420920 294578 420972 294584
rect 417424 271924 417476 271930
rect 417424 271866 417476 271872
rect 419540 271924 419592 271930
rect 419540 271866 419592 271872
rect 418160 232552 418212 232558
rect 418160 232494 418212 232500
rect 418172 231878 418200 232494
rect 418160 231872 418212 231878
rect 418160 231814 418212 231820
rect 419448 231872 419500 231878
rect 419448 231814 419500 231820
rect 417424 220108 417476 220114
rect 417424 220050 417476 220056
rect 414664 182912 414716 182918
rect 414664 182854 414716 182860
rect 414664 179512 414716 179518
rect 414664 179454 414716 179460
rect 413284 97912 413336 97918
rect 413284 97854 413336 97860
rect 396722 96520 396778 96529
rect 396722 96455 396778 96464
rect 389824 95192 389876 95198
rect 389824 95134 389876 95140
rect 414676 57866 414704 179454
rect 416778 177032 416834 177041
rect 416778 176967 416834 176976
rect 416792 176730 416820 176967
rect 416780 176724 416832 176730
rect 416780 176666 416832 176672
rect 416778 175264 416834 175273
rect 416778 175199 416834 175208
rect 416792 173942 416820 175199
rect 416780 173936 416832 173942
rect 416780 173878 416832 173884
rect 416778 168464 416834 168473
rect 416778 168399 416780 168408
rect 416832 168399 416834 168408
rect 416780 168370 416832 168376
rect 416778 166832 416834 166841
rect 416778 166767 416834 166776
rect 416792 165646 416820 166767
rect 416780 165640 416832 165646
rect 416780 165582 416832 165588
rect 416778 165064 416834 165073
rect 416778 164999 416834 165008
rect 416792 164286 416820 164999
rect 416780 164280 416832 164286
rect 416780 164222 416832 164228
rect 416778 161800 416834 161809
rect 416778 161735 416834 161744
rect 416792 161498 416820 161735
rect 416780 161492 416832 161498
rect 416780 161434 416832 161440
rect 416778 158400 416834 158409
rect 416778 158335 416834 158344
rect 416792 157418 416820 158335
rect 416780 157412 416832 157418
rect 416780 157354 416832 157360
rect 416778 156632 416834 156641
rect 416778 156567 416834 156576
rect 416792 155990 416820 156567
rect 416780 155984 416832 155990
rect 416780 155926 416832 155932
rect 416778 155000 416834 155009
rect 416778 154935 416834 154944
rect 416792 154630 416820 154935
rect 416780 154624 416832 154630
rect 416780 154566 416832 154572
rect 416780 153264 416832 153270
rect 416778 153232 416780 153241
rect 416832 153232 416834 153241
rect 416778 153167 416834 153176
rect 416778 151600 416834 151609
rect 416778 151535 416834 151544
rect 416792 150482 416820 151535
rect 416780 150476 416832 150482
rect 416780 150418 416832 150424
rect 416778 149832 416834 149841
rect 416778 149767 416834 149776
rect 416792 149122 416820 149767
rect 416780 149116 416832 149122
rect 416780 149058 416832 149064
rect 416778 148200 416834 148209
rect 416778 148135 416834 148144
rect 416792 147694 416820 148135
rect 416780 147688 416832 147694
rect 416780 147630 416832 147636
rect 416778 146568 416834 146577
rect 416778 146503 416834 146512
rect 416792 146334 416820 146503
rect 416780 146328 416832 146334
rect 416780 146270 416832 146276
rect 416870 144800 416926 144809
rect 416870 144735 416926 144744
rect 416884 143614 416912 144735
rect 416872 143608 416924 143614
rect 416872 143550 416924 143556
rect 416780 143540 416832 143546
rect 416780 143482 416832 143488
rect 416792 143177 416820 143482
rect 416778 143168 416834 143177
rect 416778 143103 416834 143112
rect 416780 142112 416832 142118
rect 416780 142054 416832 142060
rect 416792 141409 416820 142054
rect 416778 141400 416834 141409
rect 416778 141335 416834 141344
rect 416778 139768 416834 139777
rect 416778 139703 416834 139712
rect 416792 139466 416820 139703
rect 416780 139460 416832 139466
rect 416780 139402 416832 139408
rect 416778 138000 416834 138009
rect 416778 137935 416834 137944
rect 416792 136678 416820 137935
rect 416780 136672 416832 136678
rect 416780 136614 416832 136620
rect 416778 136368 416834 136377
rect 416778 136303 416834 136312
rect 416792 135318 416820 136303
rect 416780 135312 416832 135318
rect 416780 135254 416832 135260
rect 417332 135244 417384 135250
rect 417332 135186 417384 135192
rect 417344 134609 417372 135186
rect 417330 134600 417386 134609
rect 417330 134535 417386 134544
rect 417332 132456 417384 132462
rect 417332 132398 417384 132404
rect 417344 131345 417372 132398
rect 417330 131336 417386 131345
rect 417330 131271 417386 131280
rect 416780 122800 416832 122806
rect 416778 122768 416780 122777
rect 416832 122768 416834 122777
rect 416778 122703 416834 122712
rect 416780 121440 416832 121446
rect 416780 121382 416832 121388
rect 416792 121145 416820 121382
rect 416778 121136 416834 121145
rect 416778 121071 416834 121080
rect 417436 119377 417464 220050
rect 419264 182844 419316 182850
rect 419264 182786 419316 182792
rect 417516 178696 417568 178702
rect 417516 178638 417568 178644
rect 417422 119368 417478 119377
rect 417422 119303 417478 119312
rect 416780 117292 416832 117298
rect 416780 117234 416832 117240
rect 416792 116113 416820 117234
rect 416778 116104 416834 116113
rect 416778 116039 416834 116048
rect 416780 113144 416832 113150
rect 416780 113086 416832 113092
rect 416792 112713 416820 113086
rect 416778 112704 416834 112713
rect 416778 112639 416834 112648
rect 416780 111784 416832 111790
rect 416780 111726 416832 111732
rect 416792 110945 416820 111726
rect 416778 110936 416834 110945
rect 416778 110871 416834 110880
rect 416780 110424 416832 110430
rect 416780 110366 416832 110372
rect 416792 109313 416820 110366
rect 416778 109304 416834 109313
rect 416778 109239 416834 109248
rect 416780 107636 416832 107642
rect 416780 107578 416832 107584
rect 416792 107545 416820 107578
rect 416778 107536 416834 107545
rect 416778 107471 416834 107480
rect 416780 106276 416832 106282
rect 416780 106218 416832 106224
rect 416792 105913 416820 106218
rect 416778 105904 416834 105913
rect 416778 105839 416834 105848
rect 416780 104848 416832 104854
rect 416780 104790 416832 104796
rect 416792 104145 416820 104790
rect 416778 104136 416834 104145
rect 416778 104071 416834 104080
rect 416780 103488 416832 103494
rect 416780 103430 416832 103436
rect 416792 102513 416820 103430
rect 416778 102504 416834 102513
rect 416778 102439 416834 102448
rect 417528 100881 417556 178638
rect 419170 134600 419226 134609
rect 419170 134535 419226 134544
rect 417608 128308 417660 128314
rect 417608 128250 417660 128256
rect 417620 127945 417648 128250
rect 417606 127936 417662 127945
rect 417606 127871 417662 127880
rect 417514 100872 417570 100881
rect 417514 100807 417570 100816
rect 417424 96824 417476 96830
rect 417424 96766 417476 96772
rect 414664 57860 414716 57866
rect 414664 57802 414716 57808
rect 369860 42152 369912 42158
rect 369860 42094 369912 42100
rect 417436 14550 417464 96766
rect 419184 93158 419212 134535
rect 419276 127945 419304 182786
rect 419356 133884 419408 133890
rect 419356 133826 419408 133832
rect 419368 132977 419396 133826
rect 419354 132968 419410 132977
rect 419354 132903 419410 132912
rect 419262 127936 419318 127945
rect 419262 127871 419318 127880
rect 419172 93152 419224 93158
rect 419172 93094 419224 93100
rect 419368 73166 419396 132903
rect 419460 126177 419488 231814
rect 419446 126168 419502 126177
rect 419446 126103 419502 126112
rect 419552 124545 419580 271866
rect 420932 179466 420960 294578
rect 425716 210050 425744 700266
rect 429212 577522 429240 702782
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 492588 702704 492640 702710
rect 492588 702646 492640 702652
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 492600 700330 492628 702646
rect 527192 702642 527220 703520
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 521568 702568 521620 702574
rect 521568 702510 521620 702516
rect 521580 701010 521608 702510
rect 543476 702506 543504 703520
rect 559668 702574 559696 703520
rect 550548 702568 550600 702574
rect 550548 702510 550600 702516
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 519544 701004 519596 701010
rect 519544 700946 519596 700952
rect 521568 701004 521620 701010
rect 521568 700946 521620 700952
rect 492588 700324 492640 700330
rect 492588 700266 492640 700272
rect 429200 577516 429252 577522
rect 429200 577458 429252 577464
rect 429844 575544 429896 575550
rect 429844 575486 429896 575492
rect 429856 565146 429884 575486
rect 429844 565140 429896 565146
rect 429844 565082 429896 565088
rect 497464 565140 497516 565146
rect 497464 565082 497516 565088
rect 504364 565140 504416 565146
rect 504364 565082 504416 565088
rect 431224 510672 431276 510678
rect 431224 510614 431276 510620
rect 427820 340196 427872 340202
rect 427820 340138 427872 340144
rect 422300 210044 422352 210050
rect 422300 209986 422352 209992
rect 425704 210044 425756 210050
rect 425704 209986 425756 209992
rect 422312 190454 422340 209986
rect 422312 190426 422984 190454
rect 422956 179466 422984 190426
rect 425336 185700 425388 185706
rect 425336 185642 425388 185648
rect 425348 179466 425376 185642
rect 427832 179466 427860 340138
rect 431236 204270 431264 510614
rect 446404 456816 446456 456822
rect 446404 456758 446456 456764
rect 434720 248464 434772 248470
rect 434720 248406 434772 248412
rect 432604 234660 432656 234666
rect 432604 234602 432656 234608
rect 432616 211138 432644 234602
rect 432604 211132 432656 211138
rect 432604 211074 432656 211080
rect 432616 210730 432644 211074
rect 431960 210724 432012 210730
rect 431960 210666 432012 210672
rect 432604 210724 432656 210730
rect 432604 210666 432656 210672
rect 429844 204264 429896 204270
rect 429844 204206 429896 204212
rect 431224 204264 431276 204270
rect 431224 204206 431276 204212
rect 429856 203658 429884 204206
rect 429844 203652 429896 203658
rect 429844 203594 429896 203600
rect 429856 190454 429884 203594
rect 431972 190454 432000 210666
rect 429856 190426 429976 190454
rect 431972 190426 432368 190454
rect 429948 179466 429976 190426
rect 432340 179466 432368 190426
rect 434732 179466 434760 248406
rect 443644 242956 443696 242962
rect 443644 242898 443696 242904
rect 438860 238060 438912 238066
rect 438860 238002 438912 238008
rect 436100 206304 436152 206310
rect 436100 206246 436152 206252
rect 436112 190454 436140 206246
rect 438872 190454 438900 238002
rect 436112 190426 436968 190454
rect 438872 190426 439360 190454
rect 436940 179466 436968 190426
rect 439332 179466 439360 190426
rect 443656 181626 443684 242898
rect 446416 211138 446444 456758
rect 483664 379568 483716 379574
rect 483664 379510 483716 379516
rect 471980 374060 472032 374066
rect 471980 374002 472032 374008
rect 464344 368688 464396 368694
rect 464344 368630 464396 368636
rect 447784 364472 447836 364478
rect 447784 364414 447836 364420
rect 446496 215960 446548 215966
rect 446496 215902 446548 215908
rect 446404 211132 446456 211138
rect 446404 211074 446456 211080
rect 446508 181694 446536 215902
rect 444012 181688 444064 181694
rect 444012 181630 444064 181636
rect 446496 181688 446548 181694
rect 446496 181630 446548 181636
rect 441620 181620 441672 181626
rect 441620 181562 441672 181568
rect 443644 181620 443696 181626
rect 443644 181562 443696 181568
rect 441632 179466 441660 181562
rect 444024 179466 444052 181630
rect 447796 181558 447824 364414
rect 452660 360936 452712 360942
rect 452660 360878 452712 360884
rect 448520 348424 448572 348430
rect 448520 348366 448572 348372
rect 446404 181552 446456 181558
rect 446404 181494 446456 181500
rect 447784 181552 447836 181558
rect 447784 181494 447836 181500
rect 446416 179466 446444 181494
rect 448532 179466 448560 348366
rect 452672 190454 452700 360878
rect 458178 355328 458234 355337
rect 458178 355263 458234 355272
rect 454684 316736 454736 316742
rect 454684 316678 454736 316684
rect 452672 190426 453160 190454
rect 451372 181484 451424 181490
rect 451372 181426 451424 181432
rect 451384 179466 451412 181426
rect 420932 179438 421130 179466
rect 422956 179438 423430 179466
rect 425348 179438 425730 179466
rect 427832 179438 428030 179466
rect 429948 179438 430422 179466
rect 432340 179438 432722 179466
rect 434732 179438 435022 179466
rect 436940 179438 437322 179466
rect 439332 179438 439714 179466
rect 441632 179438 442014 179466
rect 444024 179438 444314 179466
rect 446416 179438 446706 179466
rect 448532 179438 449006 179466
rect 451306 179438 451412 179466
rect 453132 179466 453160 190426
rect 454696 182170 454724 316678
rect 457444 273284 457496 273290
rect 457444 273226 457496 273232
rect 457456 184278 457484 273226
rect 457444 184272 457496 184278
rect 457444 184214 457496 184220
rect 454684 182164 454736 182170
rect 454684 182106 454736 182112
rect 455604 182164 455656 182170
rect 455604 182106 455656 182112
rect 455616 179466 455644 182106
rect 458192 179466 458220 355263
rect 461584 345704 461636 345710
rect 461584 345646 461636 345652
rect 461596 182170 461624 345646
rect 461584 182164 461636 182170
rect 461584 182106 461636 182112
rect 462596 182164 462648 182170
rect 462596 182106 462648 182112
rect 460204 181688 460256 181694
rect 460204 181630 460256 181636
rect 460216 179466 460244 181630
rect 462608 179466 462636 182106
rect 464356 181694 464384 368630
rect 468484 368552 468536 368558
rect 468484 368494 468536 368500
rect 466460 362976 466512 362982
rect 466460 362918 466512 362924
rect 465080 342916 465132 342922
rect 465080 342858 465132 342864
rect 464344 181688 464396 181694
rect 464344 181630 464396 181636
rect 465092 179466 465120 342858
rect 466472 190454 466500 362918
rect 466472 190426 467144 190454
rect 467116 179466 467144 190426
rect 468496 181490 468524 368494
rect 471244 367192 471296 367198
rect 471244 367134 471296 367140
rect 469220 347064 469272 347070
rect 469220 347006 469272 347012
rect 469232 190454 469260 347006
rect 469232 190426 469536 190454
rect 468484 181484 468536 181490
rect 468484 181426 468536 181432
rect 469508 179466 469536 190426
rect 471256 184346 471284 367134
rect 471244 184340 471296 184346
rect 471244 184282 471296 184288
rect 471992 179466 472020 374002
rect 482284 327752 482336 327758
rect 482284 327694 482336 327700
rect 475384 307080 475436 307086
rect 475384 307022 475436 307028
rect 475396 218958 475424 307022
rect 478880 224256 478932 224262
rect 478880 224198 478932 224204
rect 475476 222896 475528 222902
rect 475476 222838 475528 222844
rect 475384 218952 475436 218958
rect 475384 218894 475436 218900
rect 475488 182170 475516 222838
rect 475476 182164 475528 182170
rect 475476 182106 475528 182112
rect 476580 182164 476632 182170
rect 476580 182106 476632 182112
rect 474188 181688 474240 181694
rect 474188 181630 474240 181636
rect 474200 179466 474228 181630
rect 476592 179466 476620 182106
rect 478892 179466 478920 224198
rect 480260 218952 480312 218958
rect 480260 218894 480312 218900
rect 480272 190454 480300 218894
rect 480272 190426 481128 190454
rect 481100 179466 481128 190426
rect 482296 181694 482324 327694
rect 483676 218754 483704 379510
rect 485044 361684 485096 361690
rect 485044 361626 485096 361632
rect 483664 218748 483716 218754
rect 483664 218690 483716 218696
rect 483020 210452 483072 210458
rect 483020 210394 483072 210400
rect 483032 190454 483060 210394
rect 483032 190426 483520 190454
rect 482284 181688 482336 181694
rect 482284 181630 482336 181636
rect 483492 179466 483520 190426
rect 485056 184414 485084 361626
rect 494058 356688 494114 356697
rect 494058 356623 494114 356632
rect 489184 349852 489236 349858
rect 489184 349794 489236 349800
rect 485136 225616 485188 225622
rect 485136 225558 485188 225564
rect 485044 184408 485096 184414
rect 485044 184350 485096 184356
rect 485148 182170 485176 225558
rect 486424 214668 486476 214674
rect 486424 214610 486476 214616
rect 485136 182164 485188 182170
rect 485136 182106 485188 182112
rect 485780 182164 485832 182170
rect 485780 182106 485832 182112
rect 485792 179466 485820 182106
rect 486436 181762 486464 214610
rect 488632 184340 488684 184346
rect 488632 184282 488684 184288
rect 486424 181756 486476 181762
rect 486424 181698 486476 181704
rect 488644 179466 488672 184282
rect 489196 182238 489224 349794
rect 493324 276684 493376 276690
rect 493324 276626 493376 276632
rect 490564 263628 490616 263634
rect 490564 263570 490616 263576
rect 490576 190454 490604 263570
rect 490576 190426 490696 190454
rect 489184 182232 489236 182238
rect 489184 182174 489236 182180
rect 490564 182232 490616 182238
rect 490564 182174 490616 182180
rect 453132 179438 453606 179466
rect 455616 179438 455998 179466
rect 458192 179438 458298 179466
rect 460216 179438 460598 179466
rect 462608 179438 462990 179466
rect 465092 179438 465290 179466
rect 467116 179438 467590 179466
rect 469508 179438 469890 179466
rect 471992 179438 472282 179466
rect 474200 179438 474582 179466
rect 476592 179438 476882 179466
rect 478892 179438 479274 179466
rect 481100 179438 481574 179466
rect 483492 179438 483874 179466
rect 485792 179438 486174 179466
rect 488566 179438 488672 179466
rect 490576 179466 490604 182174
rect 490668 179926 490696 190426
rect 492864 181756 492916 181762
rect 492864 181698 492916 181704
rect 490656 179920 490708 179926
rect 490656 179862 490708 179868
rect 492588 179512 492640 179518
rect 490576 179438 490866 179466
rect 492588 179454 492640 179460
rect 492876 179466 492904 181698
rect 493336 180198 493364 276626
rect 493324 180192 493376 180198
rect 493324 180134 493376 180140
rect 492600 179081 492628 179454
rect 492876 179438 493166 179466
rect 492586 179072 492642 179081
rect 492586 179007 492642 179016
rect 419632 133204 419684 133210
rect 419632 133146 419684 133152
rect 419644 129577 419672 133146
rect 419722 131336 419778 131345
rect 419722 131271 419778 131280
rect 419630 129568 419686 129577
rect 419630 129503 419686 129512
rect 419538 124536 419594 124545
rect 419538 124471 419594 124480
rect 419736 122834 419764 131271
rect 494072 129033 494100 356623
rect 497476 340202 497504 565082
rect 504376 563718 504404 565082
rect 504364 563712 504416 563718
rect 504364 563654 504416 563660
rect 512000 376780 512052 376786
rect 512000 376722 512052 376728
rect 510620 365764 510672 365770
rect 510620 365706 510672 365712
rect 508504 364336 508556 364342
rect 508504 364278 508556 364284
rect 499578 359544 499634 359553
rect 499578 359479 499634 359488
rect 497464 340196 497516 340202
rect 497464 340138 497516 340144
rect 494152 326392 494204 326398
rect 494152 326334 494204 326340
rect 494164 134745 494192 326334
rect 495440 288448 495492 288454
rect 495440 288390 495492 288396
rect 494336 188352 494388 188358
rect 494336 188294 494388 188300
rect 494242 171728 494298 171737
rect 494242 171663 494298 171672
rect 494150 134736 494206 134745
rect 494150 134671 494206 134680
rect 494058 129024 494114 129033
rect 494058 128959 494114 128968
rect 419644 122806 419764 122834
rect 419644 99346 419672 122806
rect 493966 101144 494022 101153
rect 493966 101079 494022 101088
rect 419632 99340 419684 99346
rect 419632 99282 419684 99288
rect 420184 97368 420236 97374
rect 420184 97310 420236 97316
rect 420196 93226 420224 97310
rect 420564 96830 420592 100028
rect 420932 100014 421774 100042
rect 422312 100014 422970 100042
rect 423692 100014 424166 100042
rect 425072 100014 425362 100042
rect 420552 96824 420604 96830
rect 420552 96766 420604 96772
rect 420932 93838 420960 100014
rect 421564 97300 421616 97306
rect 421564 97242 421616 97248
rect 420920 93832 420972 93838
rect 420920 93774 420972 93780
rect 420184 93220 420236 93226
rect 420184 93162 420236 93168
rect 421576 86970 421604 97242
rect 421564 86964 421616 86970
rect 421564 86906 421616 86912
rect 419356 73160 419408 73166
rect 419356 73102 419408 73108
rect 422312 45490 422340 100014
rect 422300 45484 422352 45490
rect 422300 45426 422352 45432
rect 417424 14544 417476 14550
rect 417424 14486 417476 14492
rect 423692 9654 423720 100014
rect 425072 33114 425100 100014
rect 426544 73098 426572 100028
rect 427740 97374 427768 100028
rect 427832 100014 428950 100042
rect 429212 100014 430146 100042
rect 430592 100014 431342 100042
rect 431972 100014 432538 100042
rect 433352 100014 433734 100042
rect 434732 100014 434930 100042
rect 436126 100014 436232 100042
rect 427728 97368 427780 97374
rect 427728 97310 427780 97316
rect 426532 73092 426584 73098
rect 426532 73034 426584 73040
rect 427832 43450 427860 100014
rect 427820 43444 427872 43450
rect 427820 43386 427872 43392
rect 429212 42090 429240 100014
rect 429200 42084 429252 42090
rect 429200 42026 429252 42032
rect 430592 40730 430620 100014
rect 430580 40724 430632 40730
rect 430580 40666 430632 40672
rect 425060 33108 425112 33114
rect 425060 33050 425112 33056
rect 423680 9648 423732 9654
rect 423680 9590 423732 9596
rect 431972 7614 432000 100014
rect 433352 39438 433380 100014
rect 433340 39432 433392 39438
rect 433340 39374 433392 39380
rect 434732 38622 434760 100014
rect 434720 38616 434772 38622
rect 434720 38558 434772 38564
rect 436204 36650 436232 100014
rect 436296 100014 437322 100042
rect 437492 100014 438518 100042
rect 438872 100014 439714 100042
rect 436192 36644 436244 36650
rect 436192 36586 436244 36592
rect 436296 35222 436324 100014
rect 436284 35216 436336 35222
rect 436284 35158 436336 35164
rect 437492 34474 437520 100014
rect 437480 34468 437532 34474
rect 437480 34410 437532 34416
rect 438872 31074 438900 100014
rect 440896 96966 440924 100028
rect 441632 100014 442106 100042
rect 443012 100014 443302 100042
rect 444392 100014 444498 100042
rect 445786 100014 445892 100042
rect 439504 96960 439556 96966
rect 439504 96902 439556 96908
rect 440884 96960 440936 96966
rect 440884 96902 440936 96908
rect 438860 31068 438912 31074
rect 438860 31010 438912 31016
rect 431960 7608 432012 7614
rect 431960 7550 432012 7556
rect 439516 6866 439544 96902
rect 441632 30326 441660 100014
rect 441620 30320 441672 30326
rect 441620 30262 441672 30268
rect 443012 28354 443040 100014
rect 443000 28348 443052 28354
rect 443000 28290 443052 28296
rect 444392 26994 444420 100014
rect 444380 26988 444432 26994
rect 444380 26930 444432 26936
rect 445864 25634 445892 100014
rect 445956 100014 446982 100042
rect 447152 100014 448178 100042
rect 448532 100014 449374 100042
rect 449912 100014 450570 100042
rect 451292 100014 451766 100042
rect 452672 100014 452962 100042
rect 445852 25628 445904 25634
rect 445852 25570 445904 25576
rect 445956 24206 445984 100014
rect 445944 24200 445996 24206
rect 445944 24142 445996 24148
rect 447152 22982 447180 100014
rect 447140 22976 447192 22982
rect 447140 22918 447192 22924
rect 439504 6860 439556 6866
rect 439504 6802 439556 6808
rect 363604 6792 363656 6798
rect 363604 6734 363656 6740
rect 448532 5506 448560 100014
rect 449912 22098 449940 100014
rect 449900 22092 449952 22098
rect 449900 22034 449952 22040
rect 451292 20058 451320 100014
rect 451280 20052 451332 20058
rect 451280 19994 451332 20000
rect 452672 18698 452700 100014
rect 454040 96960 454092 96966
rect 454040 96902 454092 96908
rect 452660 18692 452712 18698
rect 452660 18634 452712 18640
rect 454052 15910 454080 96902
rect 454144 17338 454172 100028
rect 455064 100014 455354 100042
rect 455432 100014 456550 100042
rect 456812 100014 457746 100042
rect 455064 96966 455092 100014
rect 455052 96960 455104 96966
rect 455052 96902 455104 96908
rect 455432 86290 455460 100014
rect 456812 87650 456840 100014
rect 458928 97306 458956 100028
rect 459572 100014 460138 100042
rect 460952 100014 461334 100042
rect 462332 100014 462530 100042
rect 458916 97300 458968 97306
rect 458916 97242 458968 97248
rect 456800 87644 456852 87650
rect 456800 87586 456852 87592
rect 455420 86284 455472 86290
rect 455420 86226 455472 86232
rect 459572 74526 459600 100014
rect 460952 84862 460980 100014
rect 461584 96960 461636 96966
rect 461584 96902 461636 96908
rect 460940 84856 460992 84862
rect 460940 84798 460992 84804
rect 461596 82142 461624 96902
rect 462332 89010 462360 100014
rect 462320 89004 462372 89010
rect 462320 88946 462372 88952
rect 463712 83502 463740 100028
rect 464908 96966 464936 100028
rect 465092 100014 466118 100042
rect 464896 96960 464948 96966
rect 464896 96902 464948 96908
rect 465092 90370 465120 100014
rect 467104 97300 467156 97306
rect 467104 97242 467156 97248
rect 465724 96960 465776 96966
rect 465724 96902 465776 96908
rect 465080 90364 465132 90370
rect 465080 90306 465132 90312
rect 463700 83496 463752 83502
rect 463700 83438 463752 83444
rect 461584 82136 461636 82142
rect 461584 82078 461636 82084
rect 465736 81394 465764 96902
rect 465724 81388 465776 81394
rect 465724 81330 465776 81336
rect 459560 74520 459612 74526
rect 459560 74462 459612 74468
rect 467116 52426 467144 97242
rect 467300 96966 467328 100028
rect 467852 100014 468510 100042
rect 469232 100014 469706 100042
rect 470612 100014 470994 100042
rect 471992 100014 472190 100042
rect 467288 96960 467340 96966
rect 467288 96902 467340 96908
rect 467104 52420 467156 52426
rect 467104 52362 467156 52368
rect 454132 17332 454184 17338
rect 454132 17274 454184 17280
rect 454040 15904 454092 15910
rect 454040 15846 454092 15852
rect 467852 13802 467880 100014
rect 469232 75206 469260 100014
rect 470612 79354 470640 100014
rect 470600 79348 470652 79354
rect 470600 79290 470652 79296
rect 471992 78674 472020 100014
rect 472624 96960 472676 96966
rect 472624 96902 472676 96908
rect 471980 78668 472032 78674
rect 471980 78610 472032 78616
rect 469220 75200 469272 75206
rect 469220 75142 469272 75148
rect 472636 69698 472664 96902
rect 473372 76537 473400 100028
rect 474568 96966 474596 100028
rect 474752 100014 475778 100042
rect 476132 100014 476974 100042
rect 477512 100014 478170 100042
rect 478892 100014 479366 100042
rect 480272 100014 480562 100042
rect 474556 96960 474608 96966
rect 474556 96902 474608 96908
rect 473358 76528 473414 76537
rect 473358 76463 473414 76472
rect 472624 69692 472676 69698
rect 472624 69634 472676 69640
rect 474752 68950 474780 100014
rect 474740 68944 474792 68950
rect 474740 68886 474792 68892
rect 476132 67590 476160 100014
rect 476120 67584 476172 67590
rect 476120 67526 476172 67532
rect 477512 66230 477540 100014
rect 477500 66224 477552 66230
rect 477500 66166 477552 66172
rect 467840 13796 467892 13802
rect 467840 13738 467892 13744
rect 478892 11762 478920 100014
rect 480272 64870 480300 100014
rect 481640 96960 481692 96966
rect 481640 96902 481692 96908
rect 480260 64864 480312 64870
rect 480260 64806 480312 64812
rect 481652 62082 481680 96902
rect 481744 62830 481772 100028
rect 482664 100014 482954 100042
rect 483032 100014 484150 100042
rect 484412 100014 485346 100042
rect 485792 100014 486542 100042
rect 482664 96966 482692 100014
rect 482652 96960 482704 96966
rect 482652 96902 482704 96908
rect 481732 62824 481784 62830
rect 481732 62766 481784 62772
rect 481640 62076 481692 62082
rect 481640 62018 481692 62024
rect 483032 60042 483060 100014
rect 483020 60036 483072 60042
rect 483020 59978 483072 59984
rect 484412 58818 484440 100014
rect 484400 58812 484452 58818
rect 484400 58754 484452 58760
rect 485792 57934 485820 100014
rect 487724 96966 487752 100028
rect 488552 100014 488934 100042
rect 489932 100014 490130 100042
rect 486424 96960 486476 96966
rect 486424 96902 486476 96908
rect 487712 96960 487764 96966
rect 487712 96902 487764 96908
rect 485780 57928 485832 57934
rect 485780 57870 485832 57876
rect 478880 11756 478932 11762
rect 478880 11698 478932 11704
rect 486436 10402 486464 96902
rect 488552 55894 488580 100014
rect 488540 55888 488592 55894
rect 488540 55830 488592 55836
rect 489932 54602 489960 100014
rect 489920 54596 489972 54602
rect 489920 54538 489972 54544
rect 491312 53174 491340 100028
rect 492508 97306 492536 100028
rect 492692 100014 493718 100042
rect 492496 97300 492548 97306
rect 492496 97242 492548 97248
rect 491300 53168 491352 53174
rect 491300 53110 491352 53116
rect 492692 51066 492720 100014
rect 493980 99278 494008 101079
rect 494060 100700 494112 100706
rect 494060 100642 494112 100648
rect 494072 100473 494100 100642
rect 494058 100464 494114 100473
rect 494058 100399 494114 100408
rect 493968 99272 494020 99278
rect 493968 99214 494020 99220
rect 494150 98696 494206 98705
rect 494150 98631 494206 98640
rect 492680 51060 492732 51066
rect 492680 51002 492732 51008
rect 494164 46238 494192 98631
rect 494256 94518 494284 171663
rect 494348 132161 494376 188294
rect 494334 132152 494390 132161
rect 494334 132087 494390 132096
rect 495452 113937 495480 288390
rect 498292 237448 498344 237454
rect 498292 237390 498344 237396
rect 496820 231124 496872 231130
rect 496820 231066 496872 231072
rect 495532 179920 495584 179926
rect 495532 179862 495584 179868
rect 495544 175982 495572 179862
rect 495532 175976 495584 175982
rect 495532 175918 495584 175924
rect 495530 169960 495586 169969
rect 495530 169895 495586 169904
rect 495438 113928 495494 113937
rect 495438 113863 495494 113872
rect 494334 103728 494390 103737
rect 494334 103663 494390 103672
rect 494348 97986 494376 103663
rect 494336 97980 494388 97986
rect 494336 97922 494388 97928
rect 494244 94512 494296 94518
rect 494244 94454 494296 94460
rect 495544 48278 495572 169895
rect 495622 168872 495678 168881
rect 495622 168807 495678 168816
rect 495636 49026 495664 168807
rect 496832 150929 496860 231066
rect 498106 175672 498162 175681
rect 498162 175630 498240 175658
rect 498106 175607 498162 175616
rect 496910 173360 496966 173369
rect 496910 173295 496966 173304
rect 496924 172582 496952 173295
rect 496912 172576 496964 172582
rect 496912 172518 496964 172524
rect 496912 168360 496964 168366
rect 496912 168302 496964 168308
rect 496924 167793 496952 168302
rect 496910 167784 496966 167793
rect 496910 167719 496966 167728
rect 496912 167000 496964 167006
rect 496912 166942 496964 166948
rect 496924 166705 496952 166942
rect 496910 166696 496966 166705
rect 496910 166631 496966 166640
rect 497004 165572 497056 165578
rect 497004 165514 497056 165520
rect 496910 165472 496966 165481
rect 496910 165407 496966 165416
rect 496924 164898 496952 165407
rect 496912 164892 496964 164898
rect 496912 164834 496964 164840
rect 497016 164393 497044 165514
rect 497002 164384 497058 164393
rect 497002 164319 497058 164328
rect 496912 164212 496964 164218
rect 496912 164154 496964 164160
rect 496924 163305 496952 164154
rect 496910 163296 496966 163305
rect 496910 163231 496966 163240
rect 496912 162852 496964 162858
rect 496912 162794 496964 162800
rect 496924 162217 496952 162794
rect 496910 162208 496966 162217
rect 496910 162143 496966 162152
rect 496912 161424 496964 161430
rect 496912 161366 496964 161372
rect 496924 160993 496952 161366
rect 496910 160984 496966 160993
rect 496910 160919 496966 160928
rect 496912 160064 496964 160070
rect 496912 160006 496964 160012
rect 496924 159905 496952 160006
rect 497004 159996 497056 160002
rect 497004 159938 497056 159944
rect 496910 159896 496966 159905
rect 496910 159831 496966 159840
rect 497016 158817 497044 159938
rect 497002 158808 497058 158817
rect 497002 158743 497058 158752
rect 496912 158704 496964 158710
rect 496912 158646 496964 158652
rect 496924 157729 496952 158646
rect 496910 157720 496966 157729
rect 496910 157655 496966 157664
rect 496912 157344 496964 157350
rect 496912 157286 496964 157292
rect 496924 156505 496952 157286
rect 496910 156496 496966 156505
rect 496910 156431 496966 156440
rect 496912 155916 496964 155922
rect 496912 155858 496964 155864
rect 496924 155417 496952 155858
rect 496910 155408 496966 155417
rect 496910 155343 496966 155352
rect 497004 154556 497056 154562
rect 497004 154498 497056 154504
rect 496912 154488 496964 154494
rect 496912 154430 496964 154436
rect 496924 153241 496952 154430
rect 497016 154329 497044 154498
rect 497002 154320 497058 154329
rect 497002 154255 497058 154264
rect 496910 153232 496966 153241
rect 496910 153167 496966 153176
rect 496912 152652 496964 152658
rect 496912 152594 496964 152600
rect 496924 152153 496952 152594
rect 496910 152144 496966 152153
rect 496910 152079 496966 152088
rect 496818 150920 496874 150929
rect 496818 150855 496874 150864
rect 496820 150408 496872 150414
rect 496820 150350 496872 150356
rect 496832 149841 496860 150350
rect 496818 149832 496874 149841
rect 496818 149767 496874 149776
rect 496820 149048 496872 149054
rect 496820 148990 496872 148996
rect 496832 148753 496860 148990
rect 496818 148744 496874 148753
rect 496818 148679 496874 148688
rect 496818 147656 496874 147665
rect 496818 147591 496820 147600
rect 496872 147591 496874 147600
rect 496820 147562 496872 147568
rect 495714 146432 495770 146441
rect 495714 146367 495770 146376
rect 495728 71738 495756 146367
rect 496820 145716 496872 145722
rect 496820 145658 496872 145664
rect 496832 145353 496860 145658
rect 496818 145344 496874 145353
rect 496818 145279 496874 145288
rect 496818 144256 496874 144265
rect 496818 144191 496874 144200
rect 496832 143614 496860 144191
rect 496820 143608 496872 143614
rect 496820 143550 496872 143556
rect 496910 143168 496966 143177
rect 496910 143103 496966 143112
rect 496924 142186 496952 143103
rect 496912 142180 496964 142186
rect 496912 142122 496964 142128
rect 496820 142112 496872 142118
rect 496820 142054 496872 142060
rect 496832 141953 496860 142054
rect 496818 141944 496874 141953
rect 496818 141879 496874 141888
rect 496820 141432 496872 141438
rect 496820 141374 496872 141380
rect 496832 140865 496860 141374
rect 496818 140856 496874 140865
rect 496818 140791 496874 140800
rect 496820 140752 496872 140758
rect 496820 140694 496872 140700
rect 496832 139777 496860 140694
rect 496818 139768 496874 139777
rect 496818 139703 496874 139712
rect 496820 139392 496872 139398
rect 496820 139334 496872 139340
rect 496832 138689 496860 139334
rect 496818 138680 496874 138689
rect 496818 138615 496874 138624
rect 496820 137964 496872 137970
rect 496820 137906 496872 137912
rect 496832 137465 496860 137906
rect 496818 137456 496874 137465
rect 496818 137391 496874 137400
rect 496912 136604 496964 136610
rect 496912 136546 496964 136552
rect 496820 136536 496872 136542
rect 496820 136478 496872 136484
rect 496832 136377 496860 136478
rect 496818 136368 496874 136377
rect 496818 136303 496874 136312
rect 496924 135289 496952 136546
rect 496910 135280 496966 135289
rect 496910 135215 496966 135224
rect 496820 133884 496872 133890
rect 496820 133826 496872 133832
rect 496832 132977 496860 133826
rect 496818 132968 496874 132977
rect 496818 132903 496874 132912
rect 496820 131096 496872 131102
rect 496820 131038 496872 131044
rect 496832 130801 496860 131038
rect 496818 130792 496874 130801
rect 496818 130727 496874 130736
rect 496820 129736 496872 129742
rect 496818 129704 496820 129713
rect 496872 129704 496874 129713
rect 496818 129639 496874 129648
rect 496820 128308 496872 128314
rect 496820 128250 496872 128256
rect 496832 127401 496860 128250
rect 496818 127392 496874 127401
rect 496818 127327 496874 127336
rect 496820 126540 496872 126546
rect 496820 126482 496872 126488
rect 496832 126313 496860 126482
rect 496818 126304 496874 126313
rect 496818 126239 496874 126248
rect 496820 125588 496872 125594
rect 496820 125530 496872 125536
rect 496832 125225 496860 125530
rect 496818 125216 496874 125225
rect 496818 125151 496874 125160
rect 496912 124160 496964 124166
rect 496818 124128 496874 124137
rect 496912 124102 496964 124108
rect 496818 124063 496820 124072
rect 496872 124063 496874 124072
rect 496820 124034 496872 124040
rect 496924 122913 496952 124102
rect 496910 122904 496966 122913
rect 496910 122839 496966 122848
rect 496820 122800 496872 122806
rect 496820 122742 496872 122748
rect 496832 121825 496860 122742
rect 496818 121816 496874 121825
rect 496818 121751 496874 121760
rect 496820 119672 496872 119678
rect 496818 119640 496820 119649
rect 496872 119640 496874 119649
rect 496818 119575 496874 119584
rect 496820 118448 496872 118454
rect 496818 118416 496820 118425
rect 496872 118416 496874 118425
rect 496818 118351 496874 118360
rect 496820 117700 496872 117706
rect 496820 117642 496872 117648
rect 496832 117337 496860 117642
rect 496818 117328 496874 117337
rect 496818 117263 496874 117272
rect 496912 117292 496964 117298
rect 496912 117234 496964 117240
rect 496924 116249 496952 117234
rect 496910 116240 496966 116249
rect 496910 116175 496966 116184
rect 496910 112840 496966 112849
rect 496910 112775 496966 112784
rect 496924 111858 496952 112775
rect 496912 111852 496964 111858
rect 496912 111794 496964 111800
rect 496820 111784 496872 111790
rect 496818 111752 496820 111761
rect 496872 111752 496874 111761
rect 496818 111687 496874 111696
rect 496820 110424 496872 110430
rect 496820 110366 496872 110372
rect 496832 109449 496860 110366
rect 496818 109440 496874 109449
rect 496818 109375 496874 109384
rect 497094 108352 497150 108361
rect 497094 108287 497150 108296
rect 497002 107264 497058 107273
rect 497002 107199 497058 107208
rect 496820 106276 496872 106282
rect 496820 106218 496872 106224
rect 496832 104961 496860 106218
rect 496910 106176 496966 106185
rect 496910 106111 496966 106120
rect 496818 104952 496874 104961
rect 496818 104887 496874 104896
rect 496924 104802 496952 106111
rect 496832 104774 496952 104802
rect 496832 100638 496860 104774
rect 497016 104666 497044 107199
rect 496924 104638 497044 104666
rect 496820 100632 496872 100638
rect 496820 100574 496872 100580
rect 496924 99210 496952 104638
rect 497108 103514 497136 108287
rect 497016 103486 497136 103514
rect 496912 99204 496964 99210
rect 496912 99146 496964 99152
rect 497016 97918 497044 103486
rect 497004 97912 497056 97918
rect 497004 97854 497056 97860
rect 495716 71732 495768 71738
rect 495716 71674 495768 71680
rect 495624 49020 495676 49026
rect 495624 48962 495676 48968
rect 495532 48272 495584 48278
rect 495532 48214 495584 48220
rect 494152 46232 494204 46238
rect 494152 46174 494204 46180
rect 498212 45558 498240 175630
rect 498304 115161 498332 237390
rect 498384 235272 498436 235278
rect 498384 235214 498436 235220
rect 498396 120737 498424 235214
rect 498476 185632 498528 185638
rect 498476 185574 498528 185580
rect 498488 152658 498516 185574
rect 498476 152652 498528 152658
rect 498476 152594 498528 152600
rect 498382 120728 498438 120737
rect 498382 120663 498438 120672
rect 499592 119678 499620 359479
rect 504364 351212 504416 351218
rect 504364 351154 504416 351160
rect 499672 320204 499724 320210
rect 499672 320146 499724 320152
rect 499684 145722 499712 320146
rect 500960 313948 501012 313954
rect 500960 313890 501012 313896
rect 499764 267028 499816 267034
rect 499764 266970 499816 266976
rect 499672 145716 499724 145722
rect 499672 145658 499724 145664
rect 499776 124098 499804 266970
rect 499854 224224 499910 224233
rect 499854 224159 499910 224168
rect 499868 126546 499896 224159
rect 499856 126540 499908 126546
rect 499856 126482 499908 126488
rect 499764 124092 499816 124098
rect 499764 124034 499816 124040
rect 499580 119672 499632 119678
rect 499580 119614 499632 119620
rect 500972 117706 501000 313890
rect 502340 240168 502392 240174
rect 502340 240110 502392 240116
rect 501144 184408 501196 184414
rect 501144 184350 501196 184356
rect 501052 172576 501104 172582
rect 501052 172518 501104 172524
rect 500960 117700 501012 117706
rect 500960 117642 501012 117648
rect 498290 115152 498346 115161
rect 498290 115087 498346 115096
rect 499580 111852 499632 111858
rect 499580 111794 499632 111800
rect 499592 95198 499620 111794
rect 501064 96626 501092 172518
rect 501156 118454 501184 184350
rect 501236 181484 501288 181490
rect 501236 181426 501288 181432
rect 501248 164898 501276 181426
rect 502352 168366 502380 240110
rect 504376 237046 504404 351154
rect 506480 287700 506532 287706
rect 506480 287642 506532 287648
rect 504364 237040 504416 237046
rect 504364 236982 504416 236988
rect 504376 236026 504404 236982
rect 503720 236020 503772 236026
rect 503720 235962 503772 235968
rect 504364 236020 504416 236026
rect 504364 235962 504416 235968
rect 502984 214600 503036 214606
rect 502984 214542 503036 214548
rect 502524 181688 502576 181694
rect 502524 181630 502576 181636
rect 502432 175976 502484 175982
rect 502432 175918 502484 175924
rect 502340 168360 502392 168366
rect 502340 168302 502392 168308
rect 501236 164892 501288 164898
rect 501236 164834 501288 164840
rect 502444 136542 502472 175918
rect 502536 154494 502564 181630
rect 502996 178702 503024 214542
rect 502984 178696 503036 178702
rect 502984 178638 503036 178644
rect 502524 154488 502576 154494
rect 502524 154430 502576 154436
rect 502996 140758 503024 178638
rect 503628 168360 503680 168366
rect 503628 168302 503680 168308
rect 503640 167686 503668 168302
rect 503628 167680 503680 167686
rect 503628 167622 503680 167628
rect 503732 160002 503760 235962
rect 505192 206372 505244 206378
rect 505192 206314 505244 206320
rect 503812 195288 503864 195294
rect 503812 195230 503864 195236
rect 503720 159996 503772 160002
rect 503720 159938 503772 159944
rect 502984 140752 503036 140758
rect 502984 140694 503036 140700
rect 502432 136536 502484 136542
rect 502432 136478 502484 136484
rect 503824 133890 503852 195230
rect 503904 191140 503956 191146
rect 503904 191082 503956 191088
rect 503916 167006 503944 191082
rect 505100 182912 505152 182918
rect 505100 182854 505152 182860
rect 503904 167000 503956 167006
rect 503904 166942 503956 166948
rect 504180 167000 504232 167006
rect 504180 166942 504232 166948
rect 504192 166326 504220 166942
rect 504180 166320 504232 166326
rect 504180 166262 504232 166268
rect 504364 164892 504416 164898
rect 504364 164834 504416 164840
rect 503812 133884 503864 133890
rect 503812 133826 503864 133832
rect 501144 118448 501196 118454
rect 501144 118390 501196 118396
rect 501052 96620 501104 96626
rect 501052 96562 501104 96568
rect 499580 95192 499632 95198
rect 499580 95134 499632 95140
rect 504376 86970 504404 164834
rect 505112 124166 505140 182854
rect 505204 149054 505232 206314
rect 505284 181620 505336 181626
rect 505284 181562 505336 181568
rect 505296 154562 505324 181562
rect 505284 154556 505336 154562
rect 505284 154498 505336 154504
rect 505192 149048 505244 149054
rect 505192 148990 505244 148996
rect 505100 124160 505152 124166
rect 505100 124102 505152 124108
rect 506492 111790 506520 287642
rect 507860 211812 507912 211818
rect 507860 211754 507912 211760
rect 506572 196648 506624 196654
rect 506572 196590 506624 196596
rect 506584 150414 506612 196590
rect 506664 184204 506716 184210
rect 506664 184146 506716 184152
rect 506676 164218 506704 184146
rect 506664 164212 506716 164218
rect 506664 164154 506716 164160
rect 506572 150408 506624 150414
rect 506572 150350 506624 150356
rect 507768 144220 507820 144226
rect 507768 144162 507820 144168
rect 507780 143614 507808 144162
rect 507768 143608 507820 143614
rect 507768 143550 507820 143556
rect 506480 111784 506532 111790
rect 506480 111726 506532 111732
rect 504364 86964 504416 86970
rect 504364 86906 504416 86912
rect 498200 45552 498252 45558
rect 498200 45494 498252 45500
rect 507780 20670 507808 143550
rect 507872 128314 507900 211754
rect 507952 181552 508004 181558
rect 507952 181494 508004 181500
rect 507860 128308 507912 128314
rect 507860 128250 507912 128256
rect 507964 106282 507992 181494
rect 508516 136610 508544 364278
rect 509332 199436 509384 199442
rect 509332 199378 509384 199384
rect 509240 180124 509292 180130
rect 509240 180066 509292 180072
rect 508504 136604 508556 136610
rect 508504 136546 508556 136552
rect 509252 131102 509280 180066
rect 509344 165578 509372 199378
rect 509332 165572 509384 165578
rect 509332 165514 509384 165520
rect 510528 165572 510580 165578
rect 510528 165514 510580 165520
rect 510540 164898 510568 165514
rect 510528 164892 510580 164898
rect 510528 164834 510580 164840
rect 509240 131096 509292 131102
rect 509240 131038 509292 131044
rect 510632 110430 510660 365706
rect 510712 221468 510764 221474
rect 510712 221410 510764 221416
rect 510724 117298 510752 221410
rect 510804 184272 510856 184278
rect 510804 184214 510856 184220
rect 510816 147626 510844 184214
rect 510804 147620 510856 147626
rect 510804 147562 510856 147568
rect 512012 144226 512040 376722
rect 517520 369912 517572 369918
rect 517520 369854 517572 369860
rect 514760 361956 514812 361962
rect 514760 361898 514812 361904
rect 513288 209092 513340 209098
rect 513288 209034 513340 209040
rect 513300 206310 513328 209034
rect 512644 206304 512696 206310
rect 512644 206246 512696 206252
rect 513288 206304 513340 206310
rect 513288 206246 513340 206252
rect 512092 180192 512144 180198
rect 512092 180134 512144 180140
rect 512000 144220 512052 144226
rect 512000 144162 512052 144168
rect 512104 142118 512132 180134
rect 512656 162858 512684 206246
rect 513380 200796 513432 200802
rect 513380 200738 513432 200744
rect 512644 162852 512696 162858
rect 512644 162794 512696 162800
rect 513288 142180 513340 142186
rect 513392 142154 513420 200738
rect 513340 142128 513420 142154
rect 513288 142126 513420 142128
rect 513288 142122 513340 142126
rect 512092 142112 512144 142118
rect 512092 142054 512144 142060
rect 510712 117292 510764 117298
rect 510712 117234 510764 117240
rect 510620 110424 510672 110430
rect 510620 110366 510672 110372
rect 507952 106276 508004 106282
rect 507952 106218 508004 106224
rect 513300 60722 513328 142122
rect 514772 129742 514800 361898
rect 514852 218748 514904 218754
rect 514852 218690 514904 218696
rect 514864 218074 514892 218690
rect 514852 218068 514904 218074
rect 514852 218010 514904 218016
rect 514864 139398 514892 218010
rect 516140 198008 516192 198014
rect 516140 197950 516192 197956
rect 516152 141438 516180 197950
rect 516140 141432 516192 141438
rect 516140 141374 516192 141380
rect 516152 140078 516180 141374
rect 516140 140072 516192 140078
rect 516140 140014 516192 140020
rect 514852 139392 514904 139398
rect 514852 139334 514904 139340
rect 514760 129736 514812 129742
rect 514760 129678 514812 129684
rect 517532 125594 517560 369854
rect 517612 207664 517664 207670
rect 517612 207606 517664 207612
rect 517624 158710 517652 207606
rect 517612 158704 517664 158710
rect 517612 158646 517664 158652
rect 519556 155922 519584 700946
rect 521580 700330 521608 700946
rect 550560 700330 550588 702510
rect 521568 700324 521620 700330
rect 521568 700266 521620 700272
rect 550548 700324 550600 700330
rect 550548 700266 550600 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580276 592686 580304 670647
rect 580264 592680 580316 592686
rect 580264 592622 580316 592628
rect 580276 592074 580304 592622
rect 580264 592068 580316 592074
rect 580264 592010 580316 592016
rect 582380 592068 582432 592074
rect 582380 592010 582432 592016
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580172 582412 580224 582418
rect 580172 582354 580224 582360
rect 580184 577697 580212 582354
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563718 580212 564295
rect 580172 563712 580224 563718
rect 580172 563654 580224 563660
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 431254 580212 431559
rect 580172 431248 580224 431254
rect 580172 431190 580224 431196
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 544384 404388 544436 404394
rect 544384 404330 544436 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 520924 260160 520976 260166
rect 520924 260102 520976 260108
rect 520936 258738 520964 260102
rect 520924 258732 520976 258738
rect 520924 258674 520976 258680
rect 519544 155916 519596 155922
rect 519544 155858 519596 155864
rect 519544 142112 519596 142118
rect 519544 142054 519596 142060
rect 517520 125588 517572 125594
rect 517520 125530 517572 125536
rect 519556 100706 519584 142054
rect 520936 137970 520964 258674
rect 529938 240816 529994 240825
rect 529938 240751 529994 240760
rect 521660 228404 521712 228410
rect 521660 228346 521712 228352
rect 520924 137964 520976 137970
rect 520924 137906 520976 137912
rect 521672 122806 521700 228346
rect 525064 164892 525116 164898
rect 525064 164834 525116 164840
rect 525076 127634 525104 164834
rect 529952 160070 529980 240751
rect 535460 239420 535512 239426
rect 535460 239362 535512 239368
rect 535472 238814 535500 239362
rect 535460 238808 535512 238814
rect 535460 238750 535512 238756
rect 535472 161430 535500 238750
rect 543004 167680 543056 167686
rect 543004 167622 543056 167628
rect 535460 161424 535512 161430
rect 535460 161366 535512 161372
rect 529940 160064 529992 160070
rect 529940 160006 529992 160012
rect 525064 127628 525116 127634
rect 525064 127570 525116 127576
rect 521660 122800 521712 122806
rect 521660 122742 521712 122748
rect 519544 100700 519596 100706
rect 519544 100642 519596 100648
rect 513288 60716 513340 60722
rect 513288 60658 513340 60664
rect 507768 20664 507820 20670
rect 507768 20606 507820 20612
rect 486424 10396 486476 10402
rect 486424 10338 486476 10344
rect 543016 6866 543044 167622
rect 544396 158710 544424 404330
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 579620 364336 579672 364342
rect 579620 364278 579672 364284
rect 579632 363662 579660 364278
rect 579620 363656 579672 363662
rect 579620 363598 579672 363604
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580184 351218 580212 351863
rect 580172 351212 580224 351218
rect 580172 351154 580224 351160
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580262 312080 580318 312089
rect 580262 312015 580318 312024
rect 580276 300150 580304 312015
rect 580264 300144 580316 300150
rect 580264 300086 580316 300092
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258738 580028 258839
rect 579988 258732 580040 258738
rect 579988 258674 580040 258680
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 239426 580212 245511
rect 580276 240825 580304 298687
rect 580262 240816 580318 240825
rect 580262 240751 580318 240760
rect 580172 239420 580224 239426
rect 580172 239362 580224 239368
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580262 192536 580318 192545
rect 580262 192471 580318 192480
rect 580276 182850 580304 192471
rect 580264 182844 580316 182850
rect 580264 182786 580316 182792
rect 580264 179444 580316 179450
rect 580264 179386 580316 179392
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 555424 166320 555476 166326
rect 555424 166262 555476 166268
rect 544384 158704 544436 158710
rect 544384 158646 544436 158652
rect 555436 46918 555464 166262
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 556160 165640 556212 165646
rect 556160 165582 556212 165588
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 556172 164218 556200 165582
rect 556160 164212 556212 164218
rect 556160 164154 556212 164160
rect 580276 152697 580304 179386
rect 582392 157350 582420 592010
rect 582380 157344 582432 157350
rect 582380 157286 582432 157292
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 140072 580224 140078
rect 580172 140014 580224 140020
rect 580184 139369 580212 140014
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 127628 580224 127634
rect 580172 127570 580224 127576
rect 580184 126041 580212 127570
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580276 99346 580304 112775
rect 580264 99340 580316 99346
rect 580264 99282 580316 99288
rect 580264 93152 580316 93158
rect 580264 93094 580316 93100
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 555424 46912 555476 46918
rect 555424 46854 555476 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 33153 580304 93094
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 543004 6860 543056 6866
rect 543004 6802 543056 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 448520 5500 448572 5506
rect 448520 5442 448572 5448
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3422 619112 3478 619168
rect 3514 606056 3570 606112
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3422 553832 3478 553888
rect 3146 527856 3202 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3514 501744 3570 501800
rect 3422 475632 3478 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3422 449520 3478 449576
rect 3422 435920 3478 435976
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3238 371320 3294 371376
rect 3422 358400 3478 358456
rect 2778 345344 2834 345400
rect 3422 319232 3478 319288
rect 3422 306176 3478 306232
rect 2778 293156 2780 293176
rect 2780 293156 2832 293176
rect 2832 293156 2834 293176
rect 2778 293120 2834 293156
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 1306 217232 1362 217288
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3330 6432 3386 6488
rect 17222 18536 17278 18592
rect 20166 10240 20222 10296
rect 33138 42064 33194 42120
rect 30838 11600 30894 11656
rect 27710 4800 27766 4856
rect 39118 14456 39174 14512
rect 40958 339360 41014 339416
rect 42522 403552 42578 403608
rect 46662 442312 46718 442368
rect 47858 404912 47914 404968
rect 42798 17176 42854 17232
rect 51722 395936 51778 395992
rect 52274 447752 52330 447808
rect 53654 487192 53710 487248
rect 53838 473184 53894 473240
rect 52274 390632 52330 390688
rect 52182 300056 52238 300112
rect 52182 206216 52238 206272
rect 56414 538056 56470 538112
rect 54206 355408 54262 355464
rect 56506 387640 56562 387696
rect 57886 389136 57942 389192
rect 58622 386416 58678 386472
rect 56506 297336 56562 297392
rect 59082 383152 59138 383208
rect 58622 353232 58678 353288
rect 60370 463528 60426 463584
rect 59174 368328 59230 368384
rect 59174 367648 59230 367704
rect 58990 335960 59046 336016
rect 61750 448588 61806 448624
rect 61750 448568 61752 448588
rect 61752 448568 61804 448588
rect 61804 448568 61806 448588
rect 61474 380976 61530 381032
rect 61934 445712 61990 445768
rect 63130 477400 63186 477456
rect 63130 382200 63186 382256
rect 67638 581204 67640 581224
rect 67640 581204 67692 581224
rect 67692 581204 67694 581224
rect 67638 581168 67694 581204
rect 66902 579128 66958 579184
rect 65890 557368 65946 557424
rect 65798 478916 65854 478952
rect 65798 478896 65800 478916
rect 65800 478896 65852 478916
rect 65852 478896 65854 478916
rect 64418 386280 64474 386336
rect 64418 349832 64474 349888
rect 64602 349696 64658 349752
rect 65982 474308 65984 474328
rect 65984 474308 66036 474328
rect 66036 474308 66038 474328
rect 65982 474272 66038 474308
rect 66074 467880 66130 467936
rect 67638 578448 67694 578504
rect 67454 577088 67510 577144
rect 67638 575728 67694 575784
rect 67638 574368 67694 574424
rect 68098 573416 68154 573472
rect 67638 572756 67694 572792
rect 67638 572736 67640 572756
rect 67640 572736 67692 572756
rect 67692 572736 67694 572756
rect 68742 576408 68798 576464
rect 67822 571648 67878 571704
rect 68466 571648 68522 571704
rect 67638 570016 67694 570072
rect 67730 568928 67786 568984
rect 67638 568656 67694 568712
rect 67638 567568 67694 567624
rect 67730 567160 67786 567216
rect 67638 565836 67640 565856
rect 67640 565836 67692 565856
rect 67692 565836 67694 565856
rect 67638 565800 67694 565836
rect 67638 564848 67694 564904
rect 67546 564440 67602 564496
rect 66994 485696 67050 485752
rect 67270 478488 67326 478544
rect 67454 481616 67510 481672
rect 67454 466792 67510 466848
rect 66166 379636 66222 379672
rect 66166 379616 66168 379636
rect 66168 379616 66220 379636
rect 66220 379616 66222 379636
rect 66166 369688 66222 369744
rect 66074 365644 66076 365664
rect 66076 365644 66128 365664
rect 66128 365644 66130 365664
rect 66074 365608 66130 365644
rect 66166 337864 66222 337920
rect 67638 563488 67694 563544
rect 67638 562300 67640 562320
rect 67640 562300 67692 562320
rect 67692 562300 67694 562320
rect 67638 562264 67694 562300
rect 67638 562128 67694 562184
rect 67730 560768 67786 560824
rect 67638 560360 67694 560416
rect 67638 559408 67694 559464
rect 67638 557540 67640 557560
rect 67640 557540 67692 557560
rect 67692 557540 67694 557560
rect 67638 557504 67694 557540
rect 67822 556688 67878 556744
rect 67638 556144 67694 556200
rect 67638 555328 67694 555384
rect 67730 554784 67786 554840
rect 67638 553444 67694 553480
rect 67638 553424 67640 553444
rect 67640 553424 67692 553444
rect 67692 553424 67694 553444
rect 67638 552084 67694 552120
rect 67638 552064 67640 552084
rect 67640 552064 67692 552084
rect 67692 552064 67694 552084
rect 67638 551248 67694 551304
rect 68650 550704 68706 550760
rect 67638 549888 67694 549944
rect 67730 548528 67786 548584
rect 67638 548004 67694 548040
rect 67638 547984 67640 548004
rect 67640 547984 67692 548004
rect 67692 547984 67694 548004
rect 67730 547168 67786 547224
rect 67638 546508 67694 546544
rect 67638 546488 67640 546508
rect 67640 546488 67692 546508
rect 67692 546488 67694 546508
rect 68558 545264 68614 545320
rect 68190 544448 68246 544504
rect 68006 543904 68062 543960
rect 67730 543088 67786 543144
rect 67638 542544 67694 542600
rect 67638 541184 67694 541240
rect 67638 540096 67694 540152
rect 67638 488008 67694 488064
rect 67638 487872 67694 487928
rect 68006 486648 68062 486704
rect 67638 485152 67694 485208
rect 67638 483676 67694 483712
rect 67638 483656 67640 483676
rect 67640 483656 67692 483676
rect 67692 483656 67694 483676
rect 68098 482432 68154 482488
rect 67638 479848 67694 479904
rect 67730 477400 67786 477456
rect 67638 476312 67694 476368
rect 67730 476176 67786 476232
rect 67638 475632 67694 475688
rect 67730 475088 67786 475144
rect 67638 474308 67640 474328
rect 67640 474308 67692 474328
rect 67692 474308 67694 474328
rect 67638 474272 67694 474308
rect 67638 472640 67694 472696
rect 67638 470872 67694 470928
rect 67730 470328 67786 470384
rect 67638 469548 67640 469568
rect 67640 469548 67692 469568
rect 67692 469548 67694 469568
rect 67638 469512 67694 469548
rect 67638 468152 67694 468208
rect 67638 465568 67694 465624
rect 67914 465432 67970 465488
rect 67638 464208 67694 464264
rect 67638 463392 67694 463448
rect 67638 461488 67694 461544
rect 67638 460164 67640 460184
rect 67640 460164 67692 460184
rect 67692 460164 67694 460184
rect 67638 460128 67694 460164
rect 67638 459992 67694 460048
rect 67730 459484 67732 459504
rect 67732 459484 67784 459504
rect 67784 459484 67786 459504
rect 67730 459448 67786 459484
rect 67638 458768 67694 458824
rect 67638 457952 67694 458008
rect 67730 457408 67786 457464
rect 67638 455912 67694 455968
rect 67638 454552 67694 454608
rect 67730 453192 67786 453248
rect 67638 452684 67640 452704
rect 67640 452684 67692 452704
rect 67692 452684 67694 452704
rect 67638 452648 67694 452684
rect 67638 451832 67694 451888
rect 67638 450744 67694 450800
rect 67822 448568 67878 448624
rect 67638 447228 67694 447264
rect 67638 447208 67640 447228
rect 67640 447208 67692 447228
rect 67692 447208 67694 447228
rect 67730 446392 67786 446448
rect 67638 445848 67694 445904
rect 67638 443692 67694 443728
rect 67638 443672 67640 443692
rect 67640 443672 67692 443692
rect 67692 443672 67694 443692
rect 67638 442468 67694 442504
rect 67638 442448 67640 442468
rect 67640 442448 67692 442468
rect 67692 442448 67694 442468
rect 67638 442312 67694 442368
rect 67638 441088 67694 441144
rect 67638 440972 67694 441008
rect 67638 440952 67640 440972
rect 67640 440952 67692 440972
rect 67692 440952 67694 440972
rect 69018 580624 69074 580680
rect 68926 572464 68982 572520
rect 68926 571784 68982 571840
rect 68834 558864 68890 558920
rect 69846 581304 69902 581360
rect 69110 545264 69166 545320
rect 68926 543904 68982 543960
rect 68742 476992 68798 477048
rect 68742 451288 68798 451344
rect 68190 444352 68246 444408
rect 68282 443808 68338 443864
rect 67730 400288 67786 400344
rect 67638 384648 67694 384704
rect 67638 382472 67694 382528
rect 67730 379752 67786 379808
rect 67638 379636 67694 379672
rect 67638 379616 67640 379636
rect 67640 379616 67692 379636
rect 67692 379616 67694 379636
rect 67546 377304 67602 377360
rect 67638 377168 67694 377224
rect 67638 375536 67694 375592
rect 67638 374620 67640 374640
rect 67640 374620 67692 374640
rect 67692 374620 67694 374640
rect 67638 374584 67694 374620
rect 67638 374176 67694 374232
rect 67638 372952 67694 373008
rect 67638 371728 67694 371784
rect 67638 368500 67640 368520
rect 67640 368500 67692 368520
rect 67692 368500 67694 368520
rect 67638 368464 67694 368500
rect 67638 367004 67640 367024
rect 67640 367004 67692 367024
rect 67692 367004 67694 367024
rect 67638 366968 67694 367004
rect 68834 444352 68890 444408
rect 68374 369452 68376 369472
rect 68376 369452 68428 369472
rect 68428 369452 68430 369472
rect 68374 369416 68430 369452
rect 68742 369416 68798 369472
rect 67638 363704 67694 363760
rect 67546 361936 67602 361992
rect 67638 360868 67694 360904
rect 67638 360848 67640 360868
rect 67640 360848 67692 360868
rect 67692 360848 67694 360868
rect 68006 360576 68062 360632
rect 67638 359508 67694 359544
rect 67638 359488 67640 359508
rect 67640 359488 67692 359508
rect 67692 359488 67694 359508
rect 67638 358708 67640 358728
rect 67640 358708 67692 358728
rect 67692 358708 67694 358728
rect 66166 189624 66222 189680
rect 66166 129240 66222 129296
rect 65154 126248 65210 126304
rect 66074 123528 66130 123584
rect 66074 102312 66130 102368
rect 66166 94832 66222 94888
rect 67638 358672 67694 358708
rect 67638 358028 67640 358048
rect 67640 358028 67692 358048
rect 67692 358028 67694 358048
rect 67638 357992 67694 358028
rect 67914 356904 67970 356960
rect 67730 355544 67786 355600
rect 67638 355136 67694 355192
rect 67638 352144 67694 352200
rect 67638 351056 67694 351112
rect 68006 350104 68062 350160
rect 67638 349052 67640 349072
rect 67640 349052 67692 349072
rect 67692 349052 67694 349072
rect 67638 349016 67694 349052
rect 68558 353096 68614 353152
rect 67638 346996 67694 347032
rect 67638 346976 67640 346996
rect 67640 346976 67692 346996
rect 67692 346976 67694 346996
rect 67638 343732 67694 343768
rect 67638 343712 67640 343732
rect 67640 343712 67692 343732
rect 67692 343712 67694 343732
rect 67638 343596 67694 343632
rect 67638 343576 67640 343596
rect 67640 343576 67692 343596
rect 67692 343576 67694 343596
rect 67638 340992 67694 341048
rect 67638 340176 67694 340232
rect 68650 344936 68706 344992
rect 68650 341944 68706 342000
rect 69018 541728 69074 541784
rect 69846 536832 69902 536888
rect 72238 582392 72294 582448
rect 81438 583888 81494 583944
rect 81806 583888 81862 583944
rect 88246 583888 88302 583944
rect 91558 583752 91614 583808
rect 91006 582528 91062 582584
rect 95146 585112 95202 585168
rect 101862 582392 101918 582448
rect 102598 581712 102654 581768
rect 105634 561856 105690 561912
rect 106922 583888 106978 583944
rect 108946 580760 109002 580816
rect 108946 579400 109002 579456
rect 108946 578040 109002 578096
rect 108854 577496 108910 577552
rect 108762 576680 108818 576736
rect 108946 576000 109002 576056
rect 108946 574640 109002 574696
rect 107658 573280 107714 573336
rect 108670 573316 108672 573336
rect 108672 573316 108724 573336
rect 108724 573316 108726 573336
rect 108670 573280 108726 573316
rect 107014 572736 107070 572792
rect 106278 560360 106334 560416
rect 73894 538056 73950 538112
rect 71042 489912 71098 489968
rect 74814 493312 74870 493368
rect 77758 526360 77814 526416
rect 80334 538056 80390 538112
rect 79322 492768 79378 492824
rect 86774 497392 86830 497448
rect 84842 496032 84898 496088
rect 89626 534656 89682 534712
rect 87050 490456 87106 490512
rect 92478 491428 92534 491464
rect 92478 491408 92480 491428
rect 92480 491408 92532 491428
rect 92532 491408 92534 491428
rect 92570 490592 92626 490648
rect 94134 490456 94190 490512
rect 94962 490456 95018 490512
rect 95790 491816 95846 491872
rect 98550 529080 98606 529136
rect 96986 491680 97042 491736
rect 97814 491680 97870 491736
rect 97446 491136 97502 491192
rect 99286 491272 99342 491328
rect 69018 488960 69074 489016
rect 68926 443808 68982 443864
rect 69846 485832 69902 485888
rect 69846 482568 69902 482624
rect 69202 482432 69258 482488
rect 69110 481480 69166 481536
rect 69662 442176 69718 442232
rect 69754 440680 69810 440736
rect 69662 440000 69718 440056
rect 70398 440000 70454 440056
rect 68926 401376 68982 401432
rect 69202 383424 69258 383480
rect 69110 380704 69166 380760
rect 74630 407496 74686 407552
rect 75274 436736 75330 436792
rect 76010 435784 76066 435840
rect 75274 407496 75330 407552
rect 75274 407088 75330 407144
rect 77482 438640 77538 438696
rect 77114 435784 77170 435840
rect 77390 435240 77446 435296
rect 78678 434560 78734 434616
rect 79690 434560 79746 434616
rect 80058 386008 80114 386064
rect 84566 437280 84622 437336
rect 85118 401648 85174 401704
rect 85486 401648 85542 401704
rect 87418 437416 87474 437472
rect 85670 403552 85726 403608
rect 85670 403008 85726 403064
rect 87418 436464 87474 436520
rect 88246 436464 88302 436520
rect 88246 405048 88302 405104
rect 89718 404912 89774 404968
rect 89718 404368 89774 404424
rect 92846 439184 92902 439240
rect 93214 439184 93270 439240
rect 92478 407768 92534 407824
rect 93674 399472 93730 399528
rect 96618 438912 96674 438968
rect 98090 439184 98146 439240
rect 97722 438912 97778 438968
rect 98090 438912 98146 438968
rect 99470 537376 99526 537432
rect 100942 536832 100998 536888
rect 101218 491408 101274 491464
rect 99470 486648 99526 486704
rect 99378 439728 99434 439784
rect 96618 397976 96674 398032
rect 77482 385328 77538 385384
rect 100114 484472 100170 484528
rect 100666 439728 100722 439784
rect 102230 489268 102232 489288
rect 102232 489268 102284 489288
rect 102284 489268 102286 489288
rect 102230 489232 102286 489268
rect 102322 488008 102378 488064
rect 102230 487872 102286 487928
rect 102230 486648 102286 486704
rect 103518 486376 103574 486432
rect 103426 485696 103482 485752
rect 103426 485152 103482 485208
rect 103426 483792 103482 483848
rect 103334 482568 103390 482624
rect 103426 482432 103482 482488
rect 103426 481480 103482 481536
rect 103334 481208 103390 481264
rect 103426 479848 103482 479904
rect 103334 479712 103390 479768
rect 103426 477672 103482 477728
rect 103242 476992 103298 477048
rect 103334 476448 103390 476504
rect 102230 475632 102286 475688
rect 102322 475088 102378 475144
rect 102230 474272 102286 474328
rect 103426 474680 103482 474736
rect 102230 472912 102286 472968
rect 102230 472232 102286 472288
rect 102230 470872 102286 470928
rect 102322 470600 102378 470656
rect 102230 470192 102286 470248
rect 102230 469512 102286 469568
rect 102230 466928 102286 466984
rect 102230 466112 102286 466168
rect 102322 465568 102378 465624
rect 102230 464752 102286 464808
rect 103334 464208 103390 464264
rect 102230 463392 102286 463448
rect 102322 462032 102378 462088
rect 102230 461488 102286 461544
rect 102414 460672 102470 460728
rect 102230 460128 102286 460184
rect 102230 459312 102286 459368
rect 102322 458768 102378 458824
rect 102322 456592 102378 456648
rect 102230 456048 102286 456104
rect 102230 455268 102232 455288
rect 102232 455268 102284 455288
rect 102284 455268 102286 455288
rect 102230 455232 102286 455268
rect 102322 454688 102378 454744
rect 102230 453872 102286 453928
rect 102322 453328 102378 453384
rect 102230 452548 102232 452568
rect 102232 452548 102284 452568
rect 102284 452548 102286 452568
rect 102230 452512 102286 452548
rect 102230 450608 102286 450664
rect 102782 450472 102838 450528
rect 102230 448568 102286 448624
rect 102230 448468 102232 448488
rect 102232 448468 102284 448488
rect 102284 448468 102286 448488
rect 102230 448432 102286 448468
rect 102322 447888 102378 447944
rect 102322 446528 102378 446584
rect 102230 445732 102286 445768
rect 102230 445712 102232 445732
rect 102232 445712 102284 445732
rect 102284 445712 102286 445732
rect 102414 445168 102470 445224
rect 102230 443808 102286 443864
rect 102230 442448 102286 442504
rect 102230 441088 102286 441144
rect 102138 391176 102194 391232
rect 101402 387776 101458 387832
rect 103426 392536 103482 392592
rect 103610 468968 103666 469024
rect 103610 466792 103666 466848
rect 103610 458088 103666 458144
rect 103610 441904 103666 441960
rect 105634 536832 105690 536888
rect 106922 548800 106978 548856
rect 105910 543768 105966 543824
rect 105174 476756 105176 476776
rect 105176 476756 105228 476776
rect 105228 476756 105230 476776
rect 105174 476720 105230 476756
rect 106278 540640 106334 540696
rect 108946 571920 109002 571976
rect 107658 571376 107714 571432
rect 107474 540096 107530 540152
rect 106278 451288 106334 451344
rect 106278 449928 106334 449984
rect 108854 570560 108910 570616
rect 108946 570036 109002 570072
rect 108946 570016 108948 570036
rect 108948 570016 109000 570036
rect 109000 570016 109002 570036
rect 108946 569200 109002 569256
rect 108854 567840 108910 567896
rect 108946 567316 109002 567352
rect 108946 567296 108948 567316
rect 108948 567296 109000 567316
rect 109000 567296 109002 567316
rect 108394 566480 108450 566536
rect 108946 565956 109002 565992
rect 108946 565936 108948 565956
rect 108948 565936 109000 565956
rect 109000 565936 109002 565956
rect 108854 565120 108910 565176
rect 108946 564476 108948 564496
rect 108948 564476 109000 564496
rect 109000 564476 109002 564496
rect 108946 564440 109002 564476
rect 108946 563896 109002 563952
rect 108946 561040 109002 561096
rect 108210 560360 108266 560416
rect 108854 559680 108910 559736
rect 108946 559020 109002 559056
rect 108946 559000 108948 559020
rect 108948 559000 109000 559020
rect 109000 559000 109002 559020
rect 108946 558320 109002 558376
rect 108302 557640 108358 557696
rect 107842 551540 107898 551576
rect 107842 551520 107844 551540
rect 107844 551520 107896 551540
rect 107896 551520 107898 551540
rect 108946 556960 109002 557016
rect 108946 555736 109002 555792
rect 108854 554240 108910 554296
rect 108946 553560 109002 553616
rect 108946 552880 109002 552936
rect 108394 552200 108450 552256
rect 108946 550840 109002 550896
rect 108854 550160 108910 550216
rect 108946 549480 109002 549536
rect 108946 547440 109002 547496
rect 108486 546760 108542 546816
rect 108946 546080 109002 546136
rect 108946 545400 109002 545456
rect 108854 544856 108910 544912
rect 108946 543360 109002 543416
rect 108946 542000 109002 542056
rect 109130 580080 109186 580136
rect 108946 399608 109002 399664
rect 111062 491272 111118 491328
rect 109038 389836 109094 389872
rect 109038 389816 109040 389836
rect 109040 389816 109092 389836
rect 109092 389816 109094 389836
rect 110326 389816 110382 389872
rect 109130 388864 109186 388920
rect 105542 385736 105598 385792
rect 111706 459584 111762 459640
rect 111982 485052 111984 485072
rect 111984 485052 112036 485072
rect 112036 485052 112038 485072
rect 111982 485016 112038 485052
rect 112442 491136 112498 491192
rect 114834 538056 114890 538112
rect 114558 482316 114614 482352
rect 114558 482296 114560 482316
rect 114560 482296 114612 482316
rect 114612 482296 114614 482316
rect 111798 386960 111854 387016
rect 112350 386552 112406 386608
rect 69294 370096 69350 370152
rect 69018 363568 69074 363624
rect 69110 360576 69166 360632
rect 68834 346332 68836 346352
rect 68836 346332 68888 346352
rect 68888 346332 68890 346352
rect 68834 346296 68890 346332
rect 69662 380704 69718 380760
rect 115754 387932 115810 387968
rect 115754 387912 115756 387932
rect 115756 387912 115808 387932
rect 115808 387912 115810 387932
rect 69478 378256 69534 378312
rect 69846 378256 69902 378312
rect 115478 376352 115534 376408
rect 115478 371864 115534 371920
rect 115570 367648 115626 367704
rect 115294 364792 115350 364848
rect 69754 340040 69810 340096
rect 67546 298152 67602 298208
rect 67638 290808 67694 290864
rect 67638 289876 67694 289912
rect 67638 289856 67640 289876
rect 67640 289856 67692 289876
rect 67692 289856 67694 289876
rect 67454 288496 67510 288552
rect 67362 246336 67418 246392
rect 67362 244296 67418 244352
rect 67638 287136 67694 287192
rect 67822 287000 67878 287056
rect 67730 286728 67786 286784
rect 68190 286048 68246 286104
rect 67638 285368 67694 285424
rect 67638 284416 67694 284472
rect 67730 283328 67786 283384
rect 67638 282104 67694 282160
rect 67638 280336 67694 280392
rect 67730 279928 67786 279984
rect 67638 279248 67694 279304
rect 67638 278568 67694 278624
rect 67638 277616 67694 277672
rect 67730 276392 67786 276448
rect 67638 275848 67694 275904
rect 67638 274896 67694 274952
rect 67730 274488 67786 274544
rect 67638 273536 67694 273592
rect 67638 272312 67694 272368
rect 68098 271496 68154 271552
rect 67730 271088 67786 271144
rect 67638 269592 67694 269648
rect 67638 268096 67694 268152
rect 67638 267028 67694 267064
rect 67638 267008 67640 267028
rect 67640 267008 67692 267028
rect 67692 267008 67694 267028
rect 67730 266872 67786 266928
rect 68834 288088 68890 288144
rect 68834 272176 68890 272232
rect 68742 266192 68798 266248
rect 67638 265648 67694 265704
rect 67730 264152 67786 264208
rect 67638 263644 67640 263664
rect 67640 263644 67692 263664
rect 67692 263644 67694 263664
rect 67638 263608 67694 263644
rect 67638 263508 67640 263528
rect 67640 263508 67692 263528
rect 67692 263508 67694 263528
rect 67638 263472 67694 263508
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67730 261432 67786 261488
rect 67822 261296 67878 261352
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 258576 67694 258632
rect 67730 258168 67786 258224
rect 67638 257896 67694 257952
rect 67638 256808 67694 256864
rect 68742 255856 68798 255912
rect 67638 255332 67694 255368
rect 67638 255312 67640 255332
rect 67640 255312 67692 255332
rect 67692 255312 67694 255332
rect 67638 255196 67694 255232
rect 67638 255176 67640 255196
rect 67640 255176 67692 255196
rect 67692 255176 67694 255196
rect 67730 254768 67786 254824
rect 67638 253852 67640 253872
rect 67640 253852 67692 253872
rect 67692 253852 67694 253872
rect 67638 253816 67694 253852
rect 67730 253408 67786 253464
rect 67638 251132 67640 251152
rect 67640 251132 67692 251152
rect 67692 251132 67694 251152
rect 67638 251096 67694 251132
rect 68558 249872 68614 249928
rect 67638 249056 67694 249112
rect 68374 248648 68430 248704
rect 67638 247696 67694 247752
rect 67546 245656 67602 245712
rect 67638 245248 67694 245304
rect 67638 243752 67694 243808
rect 67730 243616 67786 243672
rect 68926 251368 68982 251424
rect 68834 231104 68890 231160
rect 68926 198056 68982 198112
rect 69110 281288 69166 281344
rect 69110 268232 69166 268288
rect 71686 292304 71742 292360
rect 75826 339360 75882 339416
rect 77298 338680 77354 338736
rect 76562 295976 76618 296032
rect 77390 335960 77446 336016
rect 79322 337864 79378 337920
rect 89994 337728 90050 337784
rect 90914 337728 90970 337784
rect 86406 320728 86462 320784
rect 91282 297336 91338 297392
rect 91282 296792 91338 296848
rect 96526 331064 96582 331120
rect 95790 330656 95846 330712
rect 96526 330656 96582 330712
rect 97078 292576 97134 292632
rect 99286 338136 99342 338192
rect 102230 339224 102286 339280
rect 102230 338136 102286 338192
rect 104162 294480 104218 294536
rect 103150 291896 103206 291952
rect 107658 331744 107714 331800
rect 111246 337864 111302 337920
rect 111614 337864 111670 337920
rect 107382 295296 107438 295352
rect 107474 293120 107530 293176
rect 115110 339496 115166 339552
rect 114190 294616 114246 294672
rect 117502 496032 117558 496088
rect 116030 384648 116086 384704
rect 116030 360576 116086 360632
rect 115938 353948 115940 353968
rect 115940 353948 115992 353968
rect 115992 353948 115994 353968
rect 115938 353912 115994 353948
rect 117686 480800 117742 480856
rect 117410 384920 117466 384976
rect 117318 373360 117374 373416
rect 116582 369960 116638 370016
rect 117410 365200 117466 365256
rect 116122 355680 116178 355736
rect 119066 391176 119122 391232
rect 118514 384920 118570 384976
rect 118054 384240 118110 384296
rect 118146 383560 118202 383616
rect 118606 382220 118662 382256
rect 118606 382200 118608 382220
rect 118608 382200 118660 382220
rect 118660 382200 118662 382220
rect 118606 381540 118662 381576
rect 118606 381520 118608 381540
rect 118608 381520 118660 381540
rect 118660 381520 118662 381540
rect 118606 380840 118662 380896
rect 118330 379480 118386 379536
rect 118606 378800 118662 378856
rect 118054 378120 118110 378176
rect 117870 376780 117926 376816
rect 117870 376760 117872 376780
rect 117872 376760 117924 376780
rect 117924 376760 117926 376780
rect 118514 376080 118570 376136
rect 118606 375400 118662 375456
rect 118606 374040 118662 374096
rect 118054 372680 118110 372736
rect 117870 371320 117926 371376
rect 118606 370640 118662 370696
rect 118238 369980 118294 370016
rect 118238 369960 118240 369980
rect 118240 369960 118292 369980
rect 118292 369960 118294 369980
rect 118606 368600 118662 368656
rect 118606 367940 118662 367976
rect 118606 367920 118608 367940
rect 118608 367920 118660 367940
rect 118660 367920 118662 367940
rect 118606 365880 118662 365936
rect 117870 364520 117926 364576
rect 118146 363160 118202 363216
rect 118606 362480 118662 362536
rect 117594 361800 117650 361856
rect 118606 361820 118662 361856
rect 118606 361800 118608 361820
rect 118608 361800 118660 361820
rect 118660 361800 118662 361820
rect 118054 361120 118110 361176
rect 118606 359760 118662 359816
rect 118514 359080 118570 359136
rect 118606 358400 118662 358456
rect 118606 357040 118662 357096
rect 118606 356360 118662 356416
rect 118146 355680 118202 355736
rect 117778 354320 117834 354376
rect 118606 352960 118662 353016
rect 117502 351600 117558 351656
rect 118606 351600 118662 351656
rect 118054 350920 118110 350976
rect 118606 350276 118608 350296
rect 118608 350276 118660 350296
rect 118660 350276 118662 350296
rect 118606 350240 118662 350276
rect 120078 387640 120134 387696
rect 117686 348200 117742 348256
rect 117410 347520 117466 347576
rect 117502 343440 117558 343496
rect 117318 340756 117320 340776
rect 117320 340756 117372 340776
rect 117372 340756 117374 340776
rect 117318 340720 117374 340756
rect 117410 340040 117466 340096
rect 117870 342760 117926 342816
rect 118606 348880 118662 348936
rect 118514 346160 118570 346216
rect 118606 345480 118662 345536
rect 118606 344800 118662 344856
rect 118606 342080 118662 342136
rect 118974 295160 119030 295216
rect 69202 260208 69258 260264
rect 69202 251776 69258 251832
rect 119802 251096 119858 251152
rect 69846 247016 69902 247072
rect 121734 462848 121790 462904
rect 120262 358672 120318 358728
rect 122286 387912 122342 387968
rect 122194 386552 122250 386608
rect 122470 380160 122526 380216
rect 122194 376760 122250 376816
rect 122194 359216 122250 359272
rect 125690 583752 125746 583808
rect 123390 483112 123446 483168
rect 120170 295976 120226 296032
rect 121458 291760 121514 291816
rect 121550 291080 121606 291136
rect 121458 290400 121514 290456
rect 121458 289740 121514 289776
rect 121458 289720 121460 289740
rect 121460 289720 121512 289740
rect 121512 289720 121514 289740
rect 121550 289040 121606 289096
rect 121458 288380 121514 288416
rect 121458 288360 121460 288380
rect 121460 288360 121512 288380
rect 121512 288360 121514 288380
rect 121550 287680 121606 287736
rect 121458 287000 121514 287056
rect 121550 286320 121606 286376
rect 121642 285640 121698 285696
rect 121458 284960 121514 285016
rect 121550 284280 121606 284336
rect 121458 283600 121514 283656
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121550 280880 121606 280936
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121642 279520 121698 279576
rect 121458 278840 121514 278896
rect 121458 277480 121514 277536
rect 121458 276800 121514 276856
rect 121458 276120 121514 276176
rect 120170 275440 120226 275496
rect 120722 275440 120778 275496
rect 120170 250960 120226 251016
rect 120078 241440 120134 241496
rect 72422 239808 72478 239864
rect 75826 233008 75882 233064
rect 78678 200640 78734 200696
rect 86130 234504 86186 234560
rect 98366 235864 98422 235920
rect 107382 237088 107438 237144
rect 106738 235864 106794 235920
rect 69018 186904 69074 186960
rect 100666 183640 100722 183696
rect 97814 176976 97870 177032
rect 105726 180784 105782 180840
rect 117042 239672 117098 239728
rect 121458 274760 121514 274816
rect 124126 378700 124128 378720
rect 124128 378700 124180 378720
rect 124180 378700 124182 378720
rect 124126 378664 124182 378700
rect 125690 491816 125746 491872
rect 136822 581712 136878 581768
rect 125782 453872 125838 453928
rect 123666 295160 123722 295216
rect 123482 294616 123538 294672
rect 122194 282240 122250 282296
rect 121550 274080 121606 274136
rect 121458 273400 121514 273456
rect 121458 272720 121514 272776
rect 121458 271360 121514 271416
rect 121458 270000 121514 270056
rect 121458 269320 121514 269376
rect 121550 268640 121606 268696
rect 121458 267960 121514 268016
rect 121550 267280 121606 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121458 264560 121514 264616
rect 121458 263880 121514 263936
rect 121458 263200 121514 263256
rect 121550 262520 121606 262576
rect 121458 261840 121514 261896
rect 121550 261160 121606 261216
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 121642 259120 121698 259176
rect 121550 258440 121606 258496
rect 122746 278160 122802 278216
rect 122286 272040 122342 272096
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121458 255720 121514 255776
rect 121458 255040 121514 255096
rect 122102 254360 122158 254416
rect 121458 253000 121514 253056
rect 120722 239808 120778 239864
rect 121458 252320 121514 252376
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121550 249600 121606 249656
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 121550 247560 121606 247616
rect 121550 246880 121606 246936
rect 121458 246220 121514 246256
rect 121458 246200 121460 246220
rect 121460 246200 121512 246220
rect 121512 246200 121514 246220
rect 121550 245520 121606 245576
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121458 242120 121514 242176
rect 121458 240760 121514 240816
rect 121458 240080 121514 240136
rect 122194 253680 122250 253736
rect 122746 232464 122802 232520
rect 124402 293120 124458 293176
rect 123666 235864 123722 235920
rect 123482 195336 123538 195392
rect 125506 331744 125562 331800
rect 125782 309168 125838 309224
rect 125598 300056 125654 300112
rect 126334 363024 126390 363080
rect 126886 363024 126942 363080
rect 126794 343576 126850 343632
rect 126794 342932 126796 342952
rect 126796 342932 126848 342952
rect 126848 342932 126850 342952
rect 126794 342896 126850 342932
rect 126426 291896 126482 291952
rect 126334 237224 126390 237280
rect 126334 226208 126390 226264
rect 127622 442992 127678 443048
rect 131118 485016 131174 485072
rect 128634 318688 128690 318744
rect 129002 191120 129058 191176
rect 129738 288360 129794 288416
rect 129186 190984 129242 191040
rect 102046 177656 102102 177712
rect 105726 177656 105782 177712
rect 107566 177656 107622 177712
rect 98734 176704 98790 176760
rect 100666 176704 100722 176760
rect 103334 176704 103390 176760
rect 110694 177656 110750 177712
rect 112442 177656 112498 177712
rect 118422 177656 118478 177712
rect 119526 177656 119582 177712
rect 124034 177656 124090 177712
rect 125506 177656 125562 177712
rect 115846 176976 115902 177032
rect 126610 176976 126666 177032
rect 130566 251232 130622 251288
rect 134706 394848 134762 394904
rect 135166 374584 135222 374640
rect 137098 499568 137154 499624
rect 136546 389852 136548 389872
rect 136548 389852 136600 389872
rect 136600 389852 136602 389872
rect 136546 389816 136602 389852
rect 130382 178608 130438 178664
rect 133878 256708 133880 256728
rect 133880 256708 133932 256728
rect 133932 256708 133934 256728
rect 133878 256672 133934 256708
rect 137282 353948 137284 353968
rect 137284 353948 137336 353968
rect 137336 353948 137338 353968
rect 137282 353912 137338 353948
rect 140778 462324 140834 462360
rect 140778 462304 140780 462324
rect 140780 462304 140832 462324
rect 140832 462304 140834 462324
rect 140226 322088 140282 322144
rect 140686 242800 140742 242856
rect 140686 234368 140742 234424
rect 142066 462304 142122 462360
rect 142250 338020 142306 338056
rect 142250 338000 142252 338020
rect 142252 338000 142304 338020
rect 142304 338000 142306 338020
rect 143446 345616 143502 345672
rect 143906 389000 143962 389056
rect 144274 346296 144330 346352
rect 146206 356632 146262 356688
rect 146390 363568 146446 363624
rect 146482 360324 146538 360360
rect 146482 360304 146484 360324
rect 146484 360304 146536 360324
rect 146536 360304 146538 360324
rect 146298 238584 146354 238640
rect 147770 351056 147826 351112
rect 147126 298152 147182 298208
rect 148598 295296 148654 295352
rect 149702 359352 149758 359408
rect 150530 342896 150586 342952
rect 148414 197920 148470 197976
rect 151174 296792 151230 296848
rect 151174 227568 151230 227624
rect 153014 348336 153070 348392
rect 154578 375400 154634 375456
rect 155406 238720 155462 238776
rect 155314 235864 155370 235920
rect 133234 181328 133290 181384
rect 161018 230424 161074 230480
rect 129462 177656 129518 177712
rect 132406 177656 132462 177712
rect 134706 176976 134762 177032
rect 162122 177248 162178 177304
rect 104622 176740 104624 176760
rect 104624 176740 104676 176760
rect 104676 176740 104678 176760
rect 104622 176704 104678 176740
rect 108118 176704 108174 176760
rect 110326 176704 110382 176760
rect 113730 176704 113786 176760
rect 127070 176704 127126 176760
rect 133142 176704 133198 176760
rect 136086 176704 136142 176760
rect 148230 176704 148286 176760
rect 159914 176704 159970 176760
rect 128174 176432 128230 176488
rect 165434 307808 165490 307864
rect 164882 222808 164938 222864
rect 102046 175344 102102 175400
rect 116950 175344 117006 175400
rect 120814 175344 120870 175400
rect 121918 175344 121974 175400
rect 130750 175344 130806 175400
rect 167642 171536 167698 171592
rect 67362 128016 67418 128072
rect 67270 122576 67326 122632
rect 67454 125160 67510 125216
rect 67362 93744 67418 93800
rect 67638 120808 67694 120864
rect 67454 91024 67510 91080
rect 67730 100680 67786 100736
rect 67270 89664 67326 89720
rect 85578 94696 85634 94752
rect 112350 94696 112406 94752
rect 122838 94696 122894 94752
rect 124494 94696 124550 94752
rect 123206 93472 123262 93528
rect 100574 93200 100630 93256
rect 110142 93200 110198 93256
rect 74814 92384 74870 92440
rect 84842 92384 84898 92440
rect 86774 92384 86830 92440
rect 88062 92420 88064 92440
rect 88064 92420 88116 92440
rect 88116 92420 88118 92440
rect 88062 92384 88118 92420
rect 100114 92384 100170 92440
rect 101954 92384 102010 92440
rect 103426 92384 103482 92440
rect 104438 92384 104494 92440
rect 105726 92384 105782 92440
rect 107566 92384 107622 92440
rect 107934 92384 107990 92440
rect 108302 92384 108358 92440
rect 110050 92384 110106 92440
rect 88982 91704 89038 91760
rect 97446 91432 97502 91488
rect 99194 91432 99250 91488
rect 95054 91296 95110 91352
rect 90638 91160 90694 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97078 91160 97134 91216
rect 99102 91160 99158 91216
rect 99102 81368 99158 81424
rect 99286 91296 99342 91352
rect 99194 80008 99250 80064
rect 101862 92248 101918 92304
rect 103334 92248 103390 92304
rect 102046 92112 102102 92168
rect 104622 92248 104678 92304
rect 106186 92248 106242 92304
rect 107474 92248 107530 92304
rect 105726 88168 105782 88224
rect 101862 78512 101918 78568
rect 108302 86808 108358 86864
rect 110694 92384 110750 92440
rect 113822 92384 113878 92440
rect 119342 92404 119398 92440
rect 119342 92384 119344 92404
rect 119344 92384 119396 92404
rect 119396 92384 119398 92404
rect 111614 91704 111670 91760
rect 110326 91160 110382 91216
rect 107566 78376 107622 78432
rect 77298 51720 77354 51776
rect 113086 91160 113142 91216
rect 119894 92384 119950 92440
rect 129462 92384 129518 92440
rect 117134 92112 117190 92168
rect 115754 91296 115810 91352
rect 114374 91160 114430 91216
rect 115294 91160 115350 91216
rect 113086 84088 113142 84144
rect 115846 91160 115902 91216
rect 118054 91568 118110 91624
rect 118606 91160 118662 91216
rect 115846 82728 115902 82784
rect 151726 93608 151782 93664
rect 133142 92384 133198 92440
rect 136086 92384 136142 92440
rect 151542 92384 151598 92440
rect 152094 92384 152150 92440
rect 134890 91704 134946 91760
rect 120906 91568 120962 91624
rect 122102 91296 122158 91352
rect 126702 91296 126758 91352
rect 121366 91160 121422 91216
rect 122746 91160 122802 91216
rect 124126 91160 124182 91216
rect 125506 91160 125562 91216
rect 126058 91160 126114 91216
rect 126886 91160 126942 91216
rect 128266 91160 128322 91216
rect 131026 91160 131082 91216
rect 151634 91160 151690 91216
rect 169206 237224 169262 237280
rect 172426 333240 172482 333296
rect 172426 332560 172482 332616
rect 170402 182824 170458 182880
rect 167734 101360 167790 101416
rect 167918 111732 167920 111752
rect 167920 111732 167972 111752
rect 167972 111732 167974 111752
rect 167918 111696 167974 111732
rect 168010 110064 168066 110120
rect 169022 108704 169078 108760
rect 120078 37848 120134 37904
rect 125874 3304 125930 3360
rect 173162 204856 173218 204912
rect 176106 238448 176162 238504
rect 177394 335960 177450 336016
rect 179418 267008 179474 267064
rect 178682 84768 178738 84824
rect 180246 88168 180302 88224
rect 181626 288360 181682 288416
rect 186226 302232 186282 302288
rect 190366 237904 190422 237960
rect 188986 95104 189042 95160
rect 192850 251232 192906 251288
rect 193126 233824 193182 233880
rect 195334 294480 195390 294536
rect 195058 236544 195114 236600
rect 195150 235184 195206 235240
rect 197358 356244 197414 356280
rect 197358 356224 197360 356244
rect 197360 356224 197412 356244
rect 197412 356224 197414 356244
rect 198002 353640 198058 353696
rect 198646 356224 198702 356280
rect 198186 351464 198242 351520
rect 198094 349560 198150 349616
rect 197358 347384 197414 347440
rect 198094 344664 198150 344720
rect 198002 342624 198058 342680
rect 197358 340584 197414 340640
rect 197358 337864 197414 337920
rect 197726 335824 197782 335880
rect 197358 331744 197414 331800
rect 197358 329024 197414 329080
rect 197358 327140 197414 327176
rect 197358 327120 197360 327140
rect 197360 327120 197412 327140
rect 197412 327120 197414 327140
rect 197358 322360 197414 322416
rect 197358 320204 197414 320240
rect 197358 320184 197360 320204
rect 197360 320184 197412 320204
rect 197412 320184 197414 320204
rect 197358 318144 197414 318200
rect 197358 315424 197414 315480
rect 197358 313384 197414 313440
rect 197358 311344 197414 311400
rect 197358 309304 197414 309360
rect 197266 306584 197322 306640
rect 197358 302504 197414 302560
rect 197358 299920 197414 299976
rect 197358 297744 197414 297800
rect 197726 304544 197782 304600
rect 198922 333784 198978 333840
rect 198278 324944 198334 325000
rect 198646 324808 198702 324864
rect 198830 313384 198886 313440
rect 196714 293664 196770 293720
rect 195702 240216 195758 240272
rect 195886 239672 195942 239728
rect 195978 236680 196034 236736
rect 195886 236000 195942 236056
rect 197450 295704 197506 295760
rect 197450 290944 197506 291000
rect 197450 288904 197506 288960
rect 197450 286864 197506 286920
rect 197450 284144 197506 284200
rect 197450 282104 197506 282160
rect 197450 280220 197506 280256
rect 197450 280200 197452 280220
rect 197452 280200 197504 280220
rect 197504 280200 197506 280220
rect 197450 277480 197506 277536
rect 197450 275304 197506 275360
rect 197450 273284 197506 273320
rect 197450 273264 197452 273284
rect 197452 273264 197504 273284
rect 197504 273264 197506 273284
rect 197450 271224 197506 271280
rect 197450 268504 197506 268560
rect 197358 266464 197414 266520
rect 197358 264424 197414 264480
rect 197358 261704 197414 261760
rect 197358 259664 197414 259720
rect 197358 257624 197414 257680
rect 197358 255584 197414 255640
rect 197358 252864 197414 252920
rect 197450 252456 197506 252512
rect 197358 250824 197414 250880
rect 197358 248956 197360 248976
rect 197360 248956 197412 248976
rect 197412 248956 197414 248976
rect 197358 248920 197414 248956
rect 196806 242120 196862 242176
rect 198554 271224 198610 271280
rect 198094 246064 198150 246120
rect 198278 244024 198334 244080
rect 199474 361800 199530 361856
rect 206466 364384 206522 364440
rect 219346 361800 219402 361856
rect 244922 376760 244978 376816
rect 248970 361664 249026 361720
rect 249706 361700 249708 361720
rect 249708 361700 249760 361720
rect 249760 361700 249762 361720
rect 249706 361664 249762 361700
rect 300122 396208 300178 396264
rect 286322 396072 286378 396128
rect 282918 369824 282974 369880
rect 293406 363160 293462 363216
rect 292486 361936 292542 361992
rect 286598 360304 286654 360360
rect 291474 360168 291530 360224
rect 292486 360168 292542 360224
rect 300122 361800 300178 361856
rect 304354 360168 304410 360224
rect 271970 359488 272026 359544
rect 314842 359488 314898 359544
rect 319258 361664 319314 361720
rect 316866 359624 316922 359680
rect 319350 359624 319406 359680
rect 319350 359352 319406 359408
rect 319350 356632 319406 356688
rect 319350 244296 319406 244352
rect 200946 239672 201002 239728
rect 201590 238448 201646 238504
rect 198186 92248 198242 92304
rect 200762 93608 200818 93664
rect 203522 237904 203578 237960
rect 206282 233824 206338 233880
rect 204902 177248 204958 177304
rect 210238 238720 210294 238776
rect 207662 181464 207718 181520
rect 207754 91568 207810 91624
rect 207846 89664 207902 89720
rect 211894 236680 211950 236736
rect 211894 224168 211950 224224
rect 216126 228248 216182 228304
rect 209226 181464 209282 181520
rect 213918 176160 213974 176216
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214102 173304 214158 173360
rect 213918 172352 213974 172408
rect 214194 171944 214250 172000
rect 214562 170856 214618 170912
rect 213918 170720 213974 170776
rect 214654 169632 214710 169688
rect 213918 169360 213974 169416
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 168000 214066 168056
rect 213918 166912 213974 166968
rect 214010 166640 214066 166696
rect 214102 166096 214158 166152
rect 213918 165280 213974 165336
rect 213918 164092 213920 164112
rect 213920 164092 213972 164112
rect 213972 164092 213974 164112
rect 213918 164056 213974 164092
rect 214010 163376 214066 163432
rect 213918 162560 213974 162616
rect 214010 162016 214066 162072
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 214010 160792 214066 160848
rect 214470 158752 214526 158808
rect 214010 158616 214066 158672
rect 213918 158072 213974 158128
rect 213918 157292 213920 157312
rect 213920 157292 213972 157312
rect 213972 157292 213974 157312
rect 213918 157256 213974 157292
rect 213918 155896 213974 155952
rect 214010 155488 214066 155544
rect 214010 153856 214066 153912
rect 213918 153448 213974 153504
rect 213366 152632 213422 152688
rect 213918 151952 213974 152008
rect 214010 150864 214066 150920
rect 213918 150592 213974 150648
rect 214010 150048 214066 150104
rect 214654 151816 214710 151872
rect 214562 149504 214618 149560
rect 213918 148688 213974 148744
rect 214562 148008 214618 148064
rect 214010 146648 214066 146704
rect 213918 146376 213974 146432
rect 213918 144916 213920 144936
rect 213920 144916 213972 144936
rect 213972 144916 213974 144936
rect 213918 144880 213974 144916
rect 213918 143556 213920 143576
rect 213920 143556 213972 143576
rect 213972 143556 213974 143576
rect 213918 143520 213974 143556
rect 213918 142704 213974 142760
rect 214470 142316 214526 142352
rect 214470 142296 214472 142316
rect 214472 142296 214524 142316
rect 214524 142296 214526 142316
rect 214010 141344 214066 141400
rect 213918 140820 213974 140856
rect 213918 140800 213920 140820
rect 213920 140800 213972 140820
rect 213972 140800 213974 140820
rect 214010 139984 214066 140040
rect 213918 139460 213974 139496
rect 213918 139440 213920 139460
rect 213920 139440 213972 139460
rect 213972 139440 213974 139460
rect 214010 138760 214066 138816
rect 213918 138080 213974 138136
rect 213918 137400 213974 137456
rect 214010 136040 214066 136096
rect 213918 135632 213974 135688
rect 213918 134000 213974 134056
rect 214010 131416 214066 131472
rect 213918 131164 213974 131200
rect 213918 131144 213920 131164
rect 213920 131144 213972 131164
rect 213972 131144 213974 131164
rect 214010 130056 214066 130112
rect 213918 129804 213974 129840
rect 213918 129784 213920 129804
rect 213920 129784 213972 129804
rect 213972 129784 213974 129804
rect 213458 128832 213514 128888
rect 213458 128424 213514 128480
rect 213918 127064 213974 127120
rect 214010 126112 214066 126168
rect 213918 125724 213974 125760
rect 213918 125704 213920 125724
rect 213920 125704 213972 125724
rect 213972 125704 213974 125724
rect 214010 124752 214066 124808
rect 213918 124228 213974 124264
rect 213918 124208 213920 124228
rect 213920 124208 213972 124228
rect 213972 124208 213974 124228
rect 214010 123528 214066 123584
rect 213918 122868 213974 122904
rect 213918 122848 213920 122868
rect 213920 122848 213972 122868
rect 213972 122848 213974 122868
rect 214010 122168 214066 122224
rect 213918 121760 213974 121816
rect 214010 120808 214066 120864
rect 213918 120400 213974 120456
rect 214010 119584 214066 119640
rect 213458 119040 213514 119096
rect 213918 118904 213974 118960
rect 214010 117544 214066 117600
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 214010 116184 214066 116240
rect 213918 115948 213920 115968
rect 213920 115948 213972 115968
rect 213972 115948 213974 115968
rect 213918 115912 213974 115948
rect 214010 114960 214066 115016
rect 213918 114572 213974 114608
rect 213918 114552 213920 114572
rect 213920 114552 213972 114572
rect 213972 114552 213974 114572
rect 214010 113600 214066 113656
rect 213918 113228 213920 113248
rect 213920 113228 213972 113248
rect 213972 113228 213974 113248
rect 213918 113192 213974 113228
rect 214010 112240 214066 112296
rect 213918 111868 213920 111888
rect 213920 111868 213972 111888
rect 213972 111868 213974 111888
rect 213918 111832 213974 111868
rect 214010 110880 214066 110936
rect 213918 110508 213920 110528
rect 213920 110508 213972 110528
rect 213972 110508 213974 110528
rect 213918 110472 213974 110508
rect 214010 109656 214066 109712
rect 213918 109132 213974 109168
rect 213918 109112 213920 109132
rect 213920 109112 213972 109132
rect 213972 109112 213974 109132
rect 214010 108296 214066 108352
rect 213918 107772 213974 107808
rect 213918 107752 213920 107772
rect 213920 107752 213972 107772
rect 213972 107752 213974 107772
rect 214010 106936 214066 106992
rect 213918 106412 213974 106448
rect 213918 106392 213920 106412
rect 213920 106392 213972 106412
rect 213972 106392 213974 106412
rect 213918 105712 213974 105768
rect 213918 103672 213974 103728
rect 214010 102448 214066 102504
rect 213918 102312 213974 102368
rect 214010 101224 214066 101280
rect 213918 101088 213974 101144
rect 214654 143928 214710 143984
rect 213918 99728 213974 99784
rect 214010 99456 214066 99512
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 213918 95784 213974 95840
rect 214746 134136 214802 134192
rect 214562 97008 214618 97064
rect 214838 96600 214894 96656
rect 227074 235864 227130 235920
rect 226982 184320 227038 184376
rect 232594 187040 232650 187096
rect 232502 182960 232558 183016
rect 233882 180104 233938 180160
rect 239402 180240 239458 180296
rect 240874 192480 240930 192536
rect 244462 234368 244518 234424
rect 245014 178744 245070 178800
rect 235262 175888 235318 175944
rect 247958 175752 248014 175808
rect 249154 175208 249210 175264
rect 249338 173712 249394 173768
rect 249246 172760 249302 172816
rect 249154 149232 249210 149288
rect 255962 228928 256018 228984
rect 249982 169496 250038 169552
rect 251178 159568 251234 159624
rect 252466 173304 252522 173360
rect 252466 172352 252522 172408
rect 252466 171808 252522 171864
rect 252098 171400 252154 171456
rect 252466 170448 252522 170504
rect 252374 170040 252430 170096
rect 252466 169124 252468 169144
rect 252468 169124 252520 169144
rect 252520 169124 252522 169144
rect 252466 169088 252522 169124
rect 252374 168544 252430 168600
rect 252466 168136 252522 168192
rect 252466 167612 252522 167648
rect 252466 167592 252468 167612
rect 252468 167592 252520 167612
rect 252520 167592 252522 167612
rect 252466 166640 252522 166696
rect 252374 166232 252430 166288
rect 252282 165688 252338 165744
rect 252466 165280 252522 165336
rect 252374 164736 252430 164792
rect 252282 164328 252338 164384
rect 252466 163920 252522 163976
rect 252374 162968 252430 163024
rect 252466 162424 252522 162480
rect 252374 162016 252430 162072
rect 252742 167184 252798 167240
rect 252834 161472 252890 161528
rect 252466 160520 252522 160576
rect 251454 160112 251510 160168
rect 251362 159160 251418 159216
rect 251270 158752 251326 158808
rect 252190 158208 252246 158264
rect 251362 157800 251418 157856
rect 250258 155352 250314 155408
rect 251546 153448 251602 153504
rect 249798 139440 249854 139496
rect 249890 136992 249946 137048
rect 217322 135496 217378 135552
rect 216126 105304 216182 105360
rect 216126 94832 216182 94888
rect 242162 84904 242218 84960
rect 217322 80688 217378 80744
rect 243542 62872 243598 62928
rect 249154 96600 249210 96656
rect 249062 19896 249118 19952
rect 252466 157292 252468 157312
rect 252468 157292 252520 157312
rect 252520 157292 252522 157312
rect 252466 157256 252522 157292
rect 252374 156848 252430 156904
rect 252558 155896 252614 155952
rect 252466 154436 252468 154456
rect 252468 154436 252520 154456
rect 252520 154436 252522 154456
rect 252466 154400 252522 154436
rect 252374 153992 252430 154048
rect 252374 153040 252430 153096
rect 252466 152632 252522 152688
rect 252282 152088 252338 152144
rect 252466 151680 252522 151736
rect 252282 151136 252338 151192
rect 252374 150728 252430 150784
rect 252466 150184 252522 150240
rect 252282 149776 252338 149832
rect 252374 148824 252430 148880
rect 252466 148280 252522 148336
rect 252466 147464 252522 147520
rect 252098 146920 252154 146976
rect 252466 145968 252522 146024
rect 252374 145560 252430 145616
rect 252466 144064 252522 144120
rect 252374 143656 252430 143712
rect 252466 143112 252522 143168
rect 252374 142704 252430 142760
rect 252466 140392 252522 140448
rect 252374 139848 252430 139904
rect 251914 129512 251970 129568
rect 251914 125704 251970 125760
rect 252466 138488 252522 138544
rect 252466 137944 252522 138000
rect 252374 137536 252430 137592
rect 252466 136584 252522 136640
rect 252190 135632 252246 135688
rect 252374 136176 252430 136232
rect 252282 135224 252338 135280
rect 252466 134680 252522 134736
rect 252374 134272 252430 134328
rect 252466 133764 252468 133784
rect 252468 133764 252520 133784
rect 252520 133764 252522 133784
rect 252466 133728 252522 133764
rect 252374 133320 252430 133376
rect 252098 132776 252154 132832
rect 252466 132404 252468 132424
rect 252468 132404 252520 132424
rect 252520 132404 252522 132424
rect 252466 132368 252522 132404
rect 252374 131824 252430 131880
rect 252466 131416 252522 131472
rect 252466 130872 252522 130928
rect 252466 130484 252522 130520
rect 252466 130464 252468 130484
rect 252468 130464 252520 130484
rect 252520 130464 252522 130484
rect 252374 130056 252430 130112
rect 252374 129104 252430 129160
rect 252466 128560 252522 128616
rect 252466 128172 252522 128208
rect 252466 128152 252468 128172
rect 252468 128152 252520 128172
rect 252520 128152 252522 128172
rect 252374 127608 252430 127664
rect 252282 127200 252338 127256
rect 252466 126656 252522 126712
rect 252190 126248 252246 126304
rect 252374 125296 252430 125352
rect 252282 124344 252338 124400
rect 252466 124752 252522 124808
rect 252374 123936 252430 123992
rect 252466 123392 252522 123448
rect 252006 118768 252062 118824
rect 251822 117272 251878 117328
rect 251822 105576 251878 105632
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252282 121488 252338 121544
rect 252282 121080 252338 121136
rect 252466 120536 252522 120592
rect 252374 120128 252430 120184
rect 252466 119584 252522 119640
rect 252374 119176 252430 119232
rect 252466 118224 252522 118280
rect 252374 117816 252430 117872
rect 252282 116320 252338 116376
rect 252466 116864 252522 116920
rect 252374 115912 252430 115968
rect 252466 115368 252522 115424
rect 252374 114960 252430 115016
rect 252466 114436 252522 114472
rect 252466 114416 252468 114436
rect 252468 114416 252520 114436
rect 252520 114416 252522 114436
rect 252374 114008 252430 114064
rect 252282 113464 252338 113520
rect 252466 113092 252468 113112
rect 252468 113092 252520 113112
rect 252520 113092 252522 113112
rect 252466 113056 252522 113092
rect 252466 112648 252522 112704
rect 252374 112104 252430 112160
rect 252466 111732 252468 111752
rect 252468 111732 252520 111752
rect 252520 111732 252522 111752
rect 252466 111696 252522 111732
rect 252374 111152 252430 111208
rect 252466 110744 252522 110800
rect 252466 110200 252522 110256
rect 252374 109792 252430 109848
rect 252282 109248 252338 109304
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 252282 108296 252338 108352
rect 252374 107888 252430 107944
rect 252466 107480 252522 107536
rect 252374 106936 252430 106992
rect 252098 106528 252154 106584
rect 252466 105984 252522 106040
rect 252006 105032 252062 105088
rect 252466 104624 252522 104680
rect 252374 104080 252430 104136
rect 252282 103672 252338 103728
rect 251178 102176 251234 102232
rect 251914 98504 251970 98560
rect 251822 97960 251878 98016
rect 251362 97008 251418 97064
rect 251270 96192 251326 96248
rect 251178 80688 251234 80744
rect 252466 103128 252522 103184
rect 252374 102720 252430 102776
rect 252466 101768 252522 101824
rect 253294 141072 253350 141128
rect 253294 140800 253350 140856
rect 253202 101360 253258 101416
rect 252282 100816 252338 100872
rect 252466 100408 252522 100464
rect 252374 99864 252430 99920
rect 252282 99456 252338 99512
rect 252466 98912 252522 98968
rect 252190 97552 252246 97608
rect 252006 96600 252062 96656
rect 256882 175888 256938 175944
rect 253570 141752 253626 141808
rect 253570 140800 253626 140856
rect 254950 119312 255006 119368
rect 255318 87488 255374 87544
rect 260286 79328 260342 79384
rect 260286 26152 260342 26208
rect 259458 24928 259514 24984
rect 260286 24928 260342 24984
rect 261666 83408 261722 83464
rect 262218 67496 262274 67552
rect 267002 175888 267058 175944
rect 271142 195200 271198 195256
rect 270590 184184 270646 184240
rect 268566 6840 268622 6896
rect 274086 83408 274142 83464
rect 278042 46144 278098 46200
rect 276846 28192 276902 28248
rect 278226 28192 278282 28248
rect 289450 233144 289506 233200
rect 292026 226208 292082 226264
rect 280894 62736 280950 62792
rect 280894 45464 280950 45520
rect 280158 44240 280214 44296
rect 280894 44240 280950 44296
rect 286414 149640 286470 149696
rect 289174 42200 289230 42256
rect 299202 238448 299258 238504
rect 305642 238584 305698 238640
rect 304906 236544 304962 236600
rect 292026 189624 292082 189680
rect 295430 35164 295432 35184
rect 295432 35164 295484 35184
rect 295484 35164 295486 35184
rect 295430 35128 295486 35164
rect 300674 39500 300730 39536
rect 300674 39480 300676 39500
rect 300676 39480 300728 39500
rect 300728 39480 300730 39500
rect 307022 178608 307078 178664
rect 307022 175616 307078 175672
rect 306930 172216 306986 172272
rect 306746 171400 306802 171456
rect 306562 170176 306618 170232
rect 306562 168408 306618 168464
rect 307298 175208 307354 175264
rect 307114 173984 307170 174040
rect 307114 173168 307170 173224
rect 307574 174800 307630 174856
rect 307666 174392 307722 174448
rect 307574 173576 307630 173632
rect 307666 172624 307722 172680
rect 307666 171808 307722 171864
rect 307298 170992 307354 171048
rect 307666 170584 307722 170640
rect 307482 169788 307538 169824
rect 307482 169768 307484 169788
rect 307484 169768 307536 169788
rect 307536 169768 307538 169788
rect 307114 169224 307170 169280
rect 307666 168816 307722 168872
rect 307482 168000 307538 168056
rect 307390 167592 307446 167648
rect 307298 167184 307354 167240
rect 306746 165824 306802 165880
rect 307206 165416 307262 165472
rect 307022 165008 307078 165064
rect 306746 163376 306802 163432
rect 305642 162832 305698 162888
rect 306562 159976 306618 160032
rect 306562 158616 306618 158672
rect 306562 156168 306618 156224
rect 306562 154400 306618 154456
rect 306654 153584 306710 153640
rect 306930 151000 306986 151056
rect 306562 150184 306618 150240
rect 306930 149776 306986 149832
rect 306930 147600 306986 147656
rect 306930 145424 306986 145480
rect 306562 144608 306618 144664
rect 306838 141616 306894 141672
rect 307114 164192 307170 164248
rect 307114 152224 307170 152280
rect 307666 166776 307722 166832
rect 307482 166368 307538 166424
rect 307666 164600 307722 164656
rect 307574 163784 307630 163840
rect 307666 162968 307722 163024
rect 307574 162832 307630 162888
rect 307482 162424 307538 162480
rect 307574 162016 307630 162072
rect 307666 161608 307722 161664
rect 307482 161200 307538 161256
rect 307574 160792 307630 160848
rect 307666 160384 307722 160440
rect 307574 159568 307630 159624
rect 307666 159024 307722 159080
rect 307666 158208 307722 158264
rect 307482 157800 307538 157856
rect 307390 157392 307446 157448
rect 307666 156984 307722 157040
rect 307574 156576 307630 156632
rect 307574 155624 307630 155680
rect 307482 155216 307538 155272
rect 307666 154808 307722 154864
rect 307666 153992 307722 154048
rect 307666 153176 307722 153232
rect 307666 151836 307722 151872
rect 307666 151816 307668 151836
rect 307668 151816 307720 151836
rect 307720 151816 307722 151836
rect 307298 151408 307354 151464
rect 307666 150612 307722 150648
rect 307666 150592 307668 150612
rect 307668 150592 307720 150612
rect 307720 150592 307722 150612
rect 307298 149232 307354 149288
rect 307482 148824 307538 148880
rect 307574 148416 307630 148472
rect 307666 148008 307722 148064
rect 307482 147192 307538 147248
rect 307574 146784 307630 146840
rect 307666 146396 307722 146432
rect 307666 146376 307668 146396
rect 307668 146376 307720 146396
rect 307720 146376 307722 146396
rect 307482 145832 307538 145888
rect 307390 145016 307446 145072
rect 307298 143792 307354 143848
rect 307206 142432 307262 142488
rect 307114 137400 307170 137456
rect 307022 136992 307078 137048
rect 306930 133184 306986 133240
rect 307114 136176 307170 136232
rect 306562 132232 306618 132288
rect 306562 128016 306618 128072
rect 306562 126792 306618 126848
rect 305826 123256 305882 123312
rect 305734 107752 305790 107808
rect 305642 99592 305698 99648
rect 299570 3576 299626 3632
rect 300766 3576 300822 3632
rect 307022 122032 307078 122088
rect 306746 117816 306802 117872
rect 306746 113228 306748 113248
rect 306748 113228 306800 113248
rect 306800 113228 306802 113248
rect 306746 113192 306802 113228
rect 305918 111968 305974 112024
rect 306746 109792 306802 109848
rect 306930 108840 306986 108896
rect 306746 104216 306802 104272
rect 306746 102992 306802 103048
rect 306930 100816 306986 100872
rect 306746 98640 306802 98696
rect 306930 97824 306986 97880
rect 307666 144200 307722 144256
rect 307574 143384 307630 143440
rect 307666 142976 307722 143032
rect 307574 142024 307630 142080
rect 307666 140820 307722 140856
rect 307666 140800 307668 140820
rect 307668 140800 307720 140820
rect 307720 140800 307722 140820
rect 307482 140392 307538 140448
rect 307574 139984 307630 140040
rect 307666 139576 307722 139632
rect 307666 138216 307722 138272
rect 307574 138080 307630 138136
rect 307666 137808 307722 137864
rect 307482 136584 307538 136640
rect 307574 135632 307630 135688
rect 307666 135224 307722 135280
rect 307574 134816 307630 134872
rect 307666 134408 307722 134464
rect 307574 133592 307630 133648
rect 307666 132640 307722 132696
rect 307666 131824 307722 131880
rect 307574 131416 307630 131472
rect 307298 131008 307354 131064
rect 307574 130600 307630 130656
rect 307666 130192 307722 130248
rect 307574 128560 307630 128616
rect 307666 128424 307722 128480
rect 307666 127200 307722 127256
rect 307574 126384 307630 126440
rect 307666 125840 307722 125896
rect 307298 125432 307354 125488
rect 307206 124208 307262 124264
rect 307574 125024 307630 125080
rect 307666 124616 307722 124672
rect 307574 123800 307630 123856
rect 308494 152632 308550 152688
rect 308402 123392 308458 123448
rect 307666 122984 307722 123040
rect 307574 122440 307630 122496
rect 307666 121624 307722 121680
rect 307482 121216 307538 121272
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307574 119992 307630 120048
rect 307298 119040 307354 119096
rect 307666 119584 307722 119640
rect 307482 118632 307538 118688
rect 307574 118224 307630 118280
rect 307666 117408 307722 117464
rect 307482 117000 307538 117056
rect 307574 116592 307630 116648
rect 307666 116184 307722 116240
rect 307574 115640 307630 115696
rect 307666 115232 307722 115288
rect 307574 114008 307630 114064
rect 307666 113600 307722 113656
rect 307574 112648 307630 112704
rect 307666 111852 307722 111888
rect 307666 111832 307668 111852
rect 307668 111832 307720 111852
rect 307720 111832 307722 111852
rect 309690 138624 309746 138680
rect 309690 138080 309746 138136
rect 307482 111424 307538 111480
rect 307574 111016 307630 111072
rect 307666 110608 307722 110664
rect 307574 110200 307630 110256
rect 307666 109248 307722 109304
rect 307574 108432 307630 108488
rect 307666 108024 307722 108080
rect 307574 107752 307630 107808
rect 307482 107616 307538 107672
rect 307574 107208 307630 107264
rect 307482 106800 307538 106856
rect 307666 106392 307722 106448
rect 307482 105848 307538 105904
rect 307574 105440 307630 105496
rect 307666 105032 307722 105088
rect 307574 104624 307630 104680
rect 307666 103808 307722 103864
rect 307574 103400 307630 103456
rect 307666 102448 307722 102504
rect 307574 102040 307630 102096
rect 307666 100952 307722 101008
rect 307574 100408 307630 100464
rect 307666 99476 307722 99512
rect 307666 99456 307668 99476
rect 307668 99456 307720 99476
rect 307720 99456 307722 99476
rect 307666 99048 307722 99104
rect 307574 97416 307630 97472
rect 307666 96600 307722 96656
rect 307666 96192 307722 96248
rect 316774 177248 316830 177304
rect 320086 361664 320142 361720
rect 319534 307672 319590 307728
rect 319534 298152 319590 298208
rect 320086 239944 320142 240000
rect 320270 356904 320326 356960
rect 321742 358944 321798 359000
rect 322202 358944 322258 359000
rect 322202 357992 322258 358048
rect 322110 352144 322166 352200
rect 321650 347520 321706 347576
rect 322754 350104 322810 350160
rect 322478 345480 322534 345536
rect 322478 343304 322534 343360
rect 322570 341400 322626 341456
rect 322386 338680 322442 338736
rect 322478 336504 322534 336560
rect 322478 334620 322534 334656
rect 322478 334600 322480 334620
rect 322480 334600 322532 334620
rect 322532 334600 322534 334620
rect 321558 331744 321614 331800
rect 322202 331764 322258 331800
rect 322202 331744 322204 331764
rect 322204 331744 322256 331764
rect 322256 331744 322258 331764
rect 322754 329840 322810 329896
rect 322754 327700 322756 327720
rect 322756 327700 322808 327720
rect 322808 327700 322810 327720
rect 322754 327664 322810 327700
rect 320362 324944 320418 325000
rect 322478 322940 322480 322960
rect 322480 322940 322532 322960
rect 322532 322940 322534 322960
rect 322478 322904 322534 322940
rect 322846 320864 322902 320920
rect 322478 316240 322534 316296
rect 322478 314200 322534 314256
rect 322846 312160 322902 312216
rect 322478 309440 322534 309496
rect 321742 307672 321798 307728
rect 322478 305224 322534 305280
rect 322478 303184 322534 303240
rect 322570 300464 322626 300520
rect 322478 296384 322534 296440
rect 322846 293664 322902 293720
rect 322478 291624 322534 291680
rect 321558 289584 321614 289640
rect 320362 242800 320418 242856
rect 321466 242800 321522 242856
rect 320822 239808 320878 239864
rect 322478 286864 322534 286920
rect 322754 284960 322810 285016
rect 322478 282940 322534 282976
rect 322478 282920 322480 282940
rect 322480 282920 322532 282940
rect 322532 282920 322534 282940
rect 322478 280744 322534 280800
rect 321834 278024 321890 278080
rect 322202 275984 322258 276040
rect 321650 271224 321706 271280
rect 320362 230424 320418 230480
rect 321834 255584 321890 255640
rect 321742 244704 321798 244760
rect 321650 224440 321706 224496
rect 319442 177384 319498 177440
rect 313922 175616 313978 175672
rect 321374 175752 321430 175808
rect 321374 173712 321430 173768
rect 321282 172624 321338 172680
rect 321558 132640 321614 132696
rect 322386 274080 322442 274136
rect 322846 269184 322902 269240
rect 322478 267280 322534 267336
rect 322478 265104 322534 265160
rect 322478 262384 322534 262440
rect 322478 260344 322534 260400
rect 322846 258304 322902 258360
rect 322846 253544 322902 253600
rect 322478 248784 322534 248840
rect 322478 246744 322534 246800
rect 321742 162152 321798 162208
rect 322938 174664 322994 174720
rect 323122 354320 323178 354376
rect 323122 163104 323178 163160
rect 323030 160792 323086 160848
rect 322202 158616 322258 158672
rect 324318 331084 324374 331120
rect 324318 331064 324320 331084
rect 324320 331064 324372 331084
rect 324372 331064 324374 331084
rect 323582 251504 323638 251560
rect 325698 363024 325754 363080
rect 324594 331064 324650 331120
rect 328550 386416 328606 386472
rect 324318 235184 324374 235240
rect 324502 237224 324558 237280
rect 324594 234504 324650 234560
rect 324410 227568 324466 227624
rect 324318 171672 324374 171728
rect 324318 170856 324374 170912
rect 324318 169360 324374 169416
rect 324318 167728 324374 167784
rect 324318 166232 324374 166288
rect 324318 165416 324374 165472
rect 324318 163920 324374 163976
rect 324318 162424 324374 162480
rect 324318 160112 324374 160168
rect 324318 159296 324374 159352
rect 324318 157800 324374 157856
rect 324318 156984 324374 157040
rect 324502 173984 324558 174040
rect 324502 168544 324558 168600
rect 324502 167048 324558 167104
rect 324502 164736 324558 164792
rect 324410 156304 324466 156360
rect 324318 155488 324374 155544
rect 324318 153992 324374 154048
rect 324410 153176 324466 153232
rect 324318 152360 324374 152416
rect 324318 150864 324374 150920
rect 324318 150048 324374 150104
rect 324502 149640 324558 149696
rect 324410 149368 324466 149424
rect 324318 148552 324374 148608
rect 324410 147736 324466 147792
rect 324318 147056 324374 147112
rect 324318 146240 324374 146296
rect 324410 145424 324466 145480
rect 324318 143112 324374 143168
rect 324502 142432 324558 142488
rect 324318 141616 324374 141672
rect 324410 140800 324466 140856
rect 324318 138488 324374 138544
rect 324318 137844 324320 137864
rect 324320 137844 324372 137864
rect 324372 137844 324374 137864
rect 324318 137808 324374 137844
rect 324410 136992 324466 137048
rect 324318 136312 324374 136368
rect 323306 135496 323362 135552
rect 324318 134680 324374 134736
rect 324410 134000 324466 134056
rect 324318 133184 324374 133240
rect 324318 130056 324374 130112
rect 321650 129648 321706 129704
rect 324318 128560 324374 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324318 125432 324374 125488
rect 324410 124752 324466 124808
rect 324318 123936 324374 123992
rect 324410 123120 324466 123176
rect 324318 122440 324374 122496
rect 324410 121624 324466 121680
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 324318 117000 324374 117056
rect 324410 116320 324466 116376
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 321834 110472 321890 110528
rect 321650 102720 321706 102776
rect 321558 99592 321614 99648
rect 321374 98776 321430 98832
rect 321466 96620 321522 96656
rect 321466 96600 321468 96620
rect 321468 96600 321520 96620
rect 321520 96600 321522 96620
rect 321742 102176 321798 102232
rect 308402 59880 308458 59936
rect 308494 40568 308550 40624
rect 316682 43424 316738 43480
rect 317326 43444 317382 43480
rect 317326 43424 317328 43444
rect 317328 43424 317380 43444
rect 317380 43424 317382 43444
rect 324318 112376 324374 112432
rect 323030 111696 323086 111752
rect 324318 109384 324374 109440
rect 324318 107752 324374 107808
rect 324318 107072 324374 107128
rect 323122 106256 323178 106312
rect 323214 105440 323270 105496
rect 324962 151680 325018 151736
rect 324686 108568 324742 108624
rect 324410 104760 324466 104816
rect 325606 103944 325662 104000
rect 325790 143928 325846 143984
rect 325882 119312 325938 119368
rect 335450 390632 335506 390688
rect 324502 101632 324558 101688
rect 324410 97824 324466 97880
rect 324318 97008 324374 97064
rect 324594 100816 324650 100872
rect 324318 82084 324320 82104
rect 324320 82084 324372 82104
rect 324372 82084 324374 82104
rect 324318 82048 324374 82084
rect 332690 185544 332746 185600
rect 331954 86128 332010 86184
rect 336830 177248 336886 177304
rect 336922 175208 336978 175264
rect 338302 177384 338358 177440
rect 339406 78512 339462 78568
rect 337014 15136 337070 15192
rect 342350 144744 342406 144800
rect 340878 46180 340880 46200
rect 340880 46180 340932 46200
rect 340932 46180 340934 46200
rect 340878 46144 340934 46180
rect 343730 182960 343786 183016
rect 347042 182824 347098 182880
rect 346582 179968 346638 180024
rect 342166 11736 342222 11792
rect 340970 7520 341026 7576
rect 348422 3984 348478 4040
rect 353390 222808 353446 222864
rect 362958 221448 363014 221504
rect 354770 8200 354826 8256
rect 354770 7520 354826 7576
rect 369858 148280 369914 148336
rect 403714 192480 403770 192536
rect 410522 359352 410578 359408
rect 414662 360168 414718 360224
rect 396722 96464 396778 96520
rect 416778 176976 416834 177032
rect 416778 175208 416834 175264
rect 416778 168428 416834 168464
rect 416778 168408 416780 168428
rect 416780 168408 416832 168428
rect 416832 168408 416834 168428
rect 416778 166776 416834 166832
rect 416778 165008 416834 165064
rect 416778 161744 416834 161800
rect 416778 158344 416834 158400
rect 416778 156576 416834 156632
rect 416778 154944 416834 155000
rect 416778 153212 416780 153232
rect 416780 153212 416832 153232
rect 416832 153212 416834 153232
rect 416778 153176 416834 153212
rect 416778 151544 416834 151600
rect 416778 149776 416834 149832
rect 416778 148144 416834 148200
rect 416778 146512 416834 146568
rect 416870 144744 416926 144800
rect 416778 143112 416834 143168
rect 416778 141344 416834 141400
rect 416778 139712 416834 139768
rect 416778 137944 416834 138000
rect 416778 136312 416834 136368
rect 417330 134544 417386 134600
rect 417330 131280 417386 131336
rect 416778 122748 416780 122768
rect 416780 122748 416832 122768
rect 416832 122748 416834 122768
rect 416778 122712 416834 122748
rect 416778 121080 416834 121136
rect 417422 119312 417478 119368
rect 416778 116048 416834 116104
rect 416778 112648 416834 112704
rect 416778 110880 416834 110936
rect 416778 109248 416834 109304
rect 416778 107480 416834 107536
rect 416778 105848 416834 105904
rect 416778 104080 416834 104136
rect 416778 102448 416834 102504
rect 419170 134544 419226 134600
rect 417606 127880 417662 127936
rect 417514 100816 417570 100872
rect 419354 132912 419410 132968
rect 419262 127880 419318 127936
rect 419446 126112 419502 126168
rect 458178 355272 458234 355328
rect 494058 356632 494114 356688
rect 492586 179016 492642 179072
rect 419722 131280 419778 131336
rect 419630 129512 419686 129568
rect 419538 124480 419594 124536
rect 499578 359488 499634 359544
rect 494242 171672 494298 171728
rect 494150 134680 494206 134736
rect 494058 128968 494114 129024
rect 493966 101088 494022 101144
rect 473358 76472 473414 76528
rect 494058 100408 494114 100464
rect 494150 98640 494206 98696
rect 494334 132096 494390 132152
rect 495530 169904 495586 169960
rect 495438 113872 495494 113928
rect 494334 103672 494390 103728
rect 495622 168816 495678 168872
rect 498106 175616 498162 175672
rect 496910 173304 496966 173360
rect 496910 167728 496966 167784
rect 496910 166640 496966 166696
rect 496910 165416 496966 165472
rect 497002 164328 497058 164384
rect 496910 163240 496966 163296
rect 496910 162152 496966 162208
rect 496910 160928 496966 160984
rect 496910 159840 496966 159896
rect 497002 158752 497058 158808
rect 496910 157664 496966 157720
rect 496910 156440 496966 156496
rect 496910 155352 496966 155408
rect 497002 154264 497058 154320
rect 496910 153176 496966 153232
rect 496910 152088 496966 152144
rect 496818 150864 496874 150920
rect 496818 149776 496874 149832
rect 496818 148688 496874 148744
rect 496818 147620 496874 147656
rect 496818 147600 496820 147620
rect 496820 147600 496872 147620
rect 496872 147600 496874 147620
rect 495714 146376 495770 146432
rect 496818 145288 496874 145344
rect 496818 144200 496874 144256
rect 496910 143112 496966 143168
rect 496818 141888 496874 141944
rect 496818 140800 496874 140856
rect 496818 139712 496874 139768
rect 496818 138624 496874 138680
rect 496818 137400 496874 137456
rect 496818 136312 496874 136368
rect 496910 135224 496966 135280
rect 496818 132912 496874 132968
rect 496818 130736 496874 130792
rect 496818 129684 496820 129704
rect 496820 129684 496872 129704
rect 496872 129684 496874 129704
rect 496818 129648 496874 129684
rect 496818 127336 496874 127392
rect 496818 126248 496874 126304
rect 496818 125160 496874 125216
rect 496818 124092 496874 124128
rect 496818 124072 496820 124092
rect 496820 124072 496872 124092
rect 496872 124072 496874 124092
rect 496910 122848 496966 122904
rect 496818 121760 496874 121816
rect 496818 119620 496820 119640
rect 496820 119620 496872 119640
rect 496872 119620 496874 119640
rect 496818 119584 496874 119620
rect 496818 118396 496820 118416
rect 496820 118396 496872 118416
rect 496872 118396 496874 118416
rect 496818 118360 496874 118396
rect 496818 117272 496874 117328
rect 496910 116184 496966 116240
rect 496910 112784 496966 112840
rect 496818 111732 496820 111752
rect 496820 111732 496872 111752
rect 496872 111732 496874 111752
rect 496818 111696 496874 111732
rect 496818 109384 496874 109440
rect 497094 108296 497150 108352
rect 497002 107208 497058 107264
rect 496910 106120 496966 106176
rect 496818 104896 496874 104952
rect 498382 120672 498438 120728
rect 499854 224168 499910 224224
rect 498290 115096 498346 115152
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 524456 579858 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 529938 240760 529994 240816
rect 580170 378392 580226 378448
rect 579802 365064 579858 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580262 312024 580318 312080
rect 580262 298696 580318 298752
rect 580170 272176 580226 272232
rect 579986 258848 580042 258904
rect 580170 245520 580226 245576
rect 580262 240760 580318 240816
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580262 192480 580318 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580262 152632 580318 152688
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 580262 112784 580318 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580262 33088 580318 33144
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 95141 585170 95207 585173
rect 115974 585170 115980 585172
rect 95141 585168 115980 585170
rect 95141 585112 95146 585168
rect 95202 585112 115980 585168
rect 95141 585110 115980 585112
rect 95141 585107 95207 585110
rect 115974 585108 115980 585110
rect 116044 585108 116050 585172
rect 52310 583884 52316 583948
rect 52380 583946 52386 583948
rect 81433 583946 81499 583949
rect 81801 583946 81867 583949
rect 52380 583944 81867 583946
rect 52380 583888 81438 583944
rect 81494 583888 81806 583944
rect 81862 583888 81867 583944
rect 52380 583886 81867 583888
rect 52380 583884 52386 583886
rect 81433 583883 81499 583886
rect 81801 583883 81867 583886
rect 88241 583946 88307 583949
rect 106917 583946 106983 583949
rect 88241 583944 106983 583946
rect 88241 583888 88246 583944
rect 88302 583888 106922 583944
rect 106978 583888 106983 583944
rect 88241 583886 106983 583888
rect 88241 583883 88307 583886
rect 106917 583883 106983 583886
rect 91553 583810 91619 583813
rect 125685 583810 125751 583813
rect 91553 583808 125751 583810
rect 91553 583752 91558 583808
rect 91614 583752 125690 583808
rect 125746 583752 125751 583808
rect 91553 583750 125751 583752
rect 91553 583747 91619 583750
rect 125685 583747 125751 583750
rect 91001 582586 91067 582589
rect 111742 582586 111748 582588
rect 91001 582584 111748 582586
rect 91001 582528 91006 582584
rect 91062 582528 111748 582584
rect 91001 582526 111748 582528
rect 91001 582523 91067 582526
rect 111742 582524 111748 582526
rect 111812 582524 111818 582588
rect 39798 582388 39804 582452
rect 39868 582450 39874 582452
rect 72233 582450 72299 582453
rect 39868 582448 72299 582450
rect 39868 582392 72238 582448
rect 72294 582392 72299 582448
rect 39868 582390 72299 582392
rect 39868 582388 39874 582390
rect 72233 582387 72299 582390
rect 101857 582450 101923 582453
rect 124254 582450 124260 582452
rect 101857 582448 124260 582450
rect 101857 582392 101862 582448
rect 101918 582392 124260 582448
rect 101857 582390 124260 582392
rect 101857 582387 101923 582390
rect 124254 582388 124260 582390
rect 124324 582388 124330 582452
rect 102593 581770 102659 581773
rect 136817 581770 136883 581773
rect 102593 581768 136883 581770
rect 102593 581712 102598 581768
rect 102654 581712 136822 581768
rect 136878 581712 136883 581768
rect 102593 581710 136883 581712
rect 102593 581707 102659 581710
rect 136817 581707 136883 581710
rect 69841 581364 69907 581365
rect 69790 581362 69796 581364
rect 69750 581302 69796 581362
rect 69860 581360 69907 581364
rect 69902 581304 69907 581360
rect 69790 581300 69796 581302
rect 69860 581300 69907 581304
rect 69841 581299 69907 581300
rect 67633 581226 67699 581229
rect 70166 581226 70226 581468
rect 67633 581224 70226 581226
rect 67633 581168 67638 581224
rect 67694 581168 70226 581224
rect 67633 581166 70226 581168
rect 67633 581163 67699 581166
rect 108941 580818 109007 580821
rect 105892 580816 109007 580818
rect 69013 580682 69079 580685
rect 70166 580682 70226 580788
rect 105892 580760 108946 580816
rect 109002 580760 109007 580816
rect 105892 580758 109007 580760
rect 108941 580755 109007 580758
rect 69013 580680 70226 580682
rect 69013 580624 69018 580680
rect 69074 580624 70226 580680
rect 69013 580622 70226 580624
rect 69013 580619 69079 580622
rect 109125 580138 109191 580141
rect 105892 580136 109191 580138
rect -960 580002 480 580092
rect 105892 580080 109130 580136
rect 109186 580080 109191 580136
rect 105892 580078 109191 580080
rect 109125 580075 109191 580078
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 108941 579458 109007 579461
rect 105892 579456 109007 579458
rect 66897 579186 66963 579189
rect 70166 579186 70226 579428
rect 105892 579400 108946 579456
rect 109002 579400 109007 579456
rect 105892 579398 109007 579400
rect 108941 579395 109007 579398
rect 66897 579184 70226 579186
rect 66897 579128 66902 579184
rect 66958 579128 70226 579184
rect 66897 579126 70226 579128
rect 66897 579123 66963 579126
rect 107694 578778 107700 578780
rect 67633 578506 67699 578509
rect 70166 578506 70226 578748
rect 105892 578718 107700 578778
rect 107694 578716 107700 578718
rect 107764 578716 107770 578780
rect 67633 578504 70226 578506
rect 67633 578448 67638 578504
rect 67694 578448 70226 578504
rect 67633 578446 70226 578448
rect 67633 578443 67699 578446
rect 108941 578098 109007 578101
rect 105892 578096 109007 578098
rect 66110 577764 66116 577828
rect 66180 577826 66186 577828
rect 70166 577826 70226 578068
rect 105892 578040 108946 578096
rect 109002 578040 109007 578096
rect 105892 578038 109007 578040
rect 108941 578035 109007 578038
rect 66180 577766 70226 577826
rect 66180 577764 66186 577766
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 108849 577554 108915 577557
rect 110638 577554 110644 577556
rect 105892 577552 110644 577554
rect 105892 577496 108854 577552
rect 108910 577496 110644 577552
rect 105892 577494 110644 577496
rect 108849 577491 108915 577494
rect 110638 577492 110644 577494
rect 110708 577492 110714 577556
rect 583520 577540 584960 577630
rect 67449 577146 67515 577149
rect 70166 577146 70226 577388
rect 67449 577144 70226 577146
rect 67449 577088 67454 577144
rect 67510 577088 70226 577144
rect 67449 577086 70226 577088
rect 67449 577083 67515 577086
rect 108757 576738 108823 576741
rect 105892 576736 108823 576738
rect 68737 576466 68803 576469
rect 70166 576466 70226 576708
rect 105892 576680 108762 576736
rect 108818 576680 108823 576736
rect 105892 576678 108823 576680
rect 108757 576675 108823 576678
rect 68737 576464 70226 576466
rect 68737 576408 68742 576464
rect 68798 576408 70226 576464
rect 68737 576406 70226 576408
rect 68737 576403 68803 576406
rect 108941 576058 109007 576061
rect 105892 576056 109007 576058
rect 67633 575786 67699 575789
rect 70166 575786 70226 576028
rect 105892 576000 108946 576056
rect 109002 576000 109007 576056
rect 105892 575998 109007 576000
rect 108941 575995 109007 575998
rect 67633 575784 70226 575786
rect 67633 575728 67638 575784
rect 67694 575728 70226 575784
rect 67633 575726 70226 575728
rect 67633 575723 67699 575726
rect 64638 575044 64644 575108
rect 64708 575106 64714 575108
rect 70166 575106 70226 575348
rect 64708 575046 70226 575106
rect 64708 575044 64714 575046
rect 108941 574698 109007 574701
rect 105892 574696 109007 574698
rect 67633 574426 67699 574429
rect 70166 574426 70226 574668
rect 105892 574640 108946 574696
rect 109002 574640 109007 574696
rect 105892 574638 109007 574640
rect 108941 574635 109007 574638
rect 67633 574424 70226 574426
rect 67633 574368 67638 574424
rect 67694 574368 70226 574424
rect 67633 574366 70226 574368
rect 67633 574363 67699 574366
rect 68093 573474 68159 573477
rect 70166 573474 70226 573988
rect 105862 573746 105922 573988
rect 105862 573686 113190 573746
rect 68093 573472 70226 573474
rect 68093 573416 68098 573472
rect 68154 573416 70226 573472
rect 68093 573414 70226 573416
rect 68093 573411 68159 573414
rect 107653 573338 107719 573341
rect 108665 573338 108731 573341
rect 105892 573336 108731 573338
rect 105892 573280 107658 573336
rect 107714 573280 108670 573336
rect 108726 573280 108731 573336
rect 105892 573278 108731 573280
rect 107653 573275 107719 573278
rect 108665 573275 108731 573278
rect 113130 573202 113190 573686
rect 114502 573202 114508 573204
rect 113130 573142 114508 573202
rect 114502 573140 114508 573142
rect 114572 573140 114578 573204
rect 67633 572794 67699 572797
rect 107009 572794 107075 572797
rect 67633 572792 70042 572794
rect 67633 572736 67638 572792
rect 67694 572736 70042 572792
rect 105892 572792 107075 572794
rect 67633 572734 70042 572736
rect 67633 572731 67699 572734
rect 69982 572730 70042 572734
rect 70166 572730 70226 572764
rect 105892 572736 107014 572792
rect 107070 572736 107075 572792
rect 105892 572734 107075 572736
rect 107009 572731 107075 572734
rect 69982 572670 70226 572730
rect 68921 572522 68987 572525
rect 68921 572520 70226 572522
rect 68921 572464 68926 572520
rect 68982 572464 70226 572520
rect 68921 572462 70226 572464
rect 68921 572459 68987 572462
rect 70166 572084 70226 572462
rect 55070 571916 55076 571980
rect 55140 571978 55146 571980
rect 108941 571978 109007 571981
rect 55140 571918 64890 571978
rect 105892 571976 109007 571978
rect 105892 571920 108946 571976
rect 109002 571920 109007 571976
rect 105892 571918 109007 571920
rect 55140 571916 55146 571918
rect 64830 571842 64890 571918
rect 108941 571915 109007 571918
rect 68921 571842 68987 571845
rect 64830 571840 68987 571842
rect 64830 571784 68926 571840
rect 68982 571784 68987 571840
rect 64830 571782 68987 571784
rect 68921 571779 68987 571782
rect 67817 571706 67883 571709
rect 68461 571706 68527 571709
rect 67817 571704 70226 571706
rect 67817 571648 67822 571704
rect 67878 571648 68466 571704
rect 68522 571648 70226 571704
rect 67817 571646 70226 571648
rect 67817 571643 67883 571646
rect 68461 571643 68527 571646
rect 70166 571404 70226 571646
rect 107653 571434 107719 571437
rect 105892 571432 107719 571434
rect 105892 571376 107658 571432
rect 107714 571376 107719 571432
rect 105892 571374 107719 571376
rect 107653 571371 107719 571374
rect 108849 570618 108915 570621
rect 105892 570616 108915 570618
rect 70166 570346 70226 570588
rect 105892 570560 108854 570616
rect 108910 570560 108915 570616
rect 105892 570558 108915 570560
rect 108849 570555 108915 570558
rect 64830 570286 70226 570346
rect 62982 570148 62988 570212
rect 63052 570210 63058 570212
rect 64830 570210 64890 570286
rect 63052 570150 64890 570210
rect 63052 570148 63058 570150
rect 67633 570074 67699 570077
rect 108941 570074 109007 570077
rect 67633 570072 70042 570074
rect 67633 570016 67638 570072
rect 67694 570016 70042 570072
rect 67633 570014 70042 570016
rect 105892 570072 109007 570074
rect 105892 570016 108946 570072
rect 109002 570016 109007 570072
rect 105892 570014 109007 570016
rect 67633 570011 67699 570014
rect 69982 569802 70042 570014
rect 108941 570011 109007 570014
rect 70166 569802 70226 569908
rect 69982 569742 70226 569802
rect 108941 569258 109007 569261
rect 105892 569256 109007 569258
rect 67725 568986 67791 568989
rect 70166 568986 70226 569228
rect 105892 569200 108946 569256
rect 109002 569200 109007 569256
rect 105892 569198 109007 569200
rect 108941 569195 109007 569198
rect 67725 568984 70226 568986
rect 67725 568928 67730 568984
rect 67786 568928 70226 568984
rect 67725 568926 70226 568928
rect 67725 568923 67791 568926
rect 67633 568714 67699 568717
rect 67633 568712 70042 568714
rect 67633 568656 67638 568712
rect 67694 568680 70042 568712
rect 70166 568680 70226 568684
rect 67694 568656 70226 568680
rect 67633 568654 70226 568656
rect 67633 568651 67699 568654
rect 69982 568620 70226 568654
rect 108849 567898 108915 567901
rect 105892 567896 108915 567898
rect 67633 567626 67699 567629
rect 70166 567626 70226 567868
rect 105892 567840 108854 567896
rect 108910 567840 108915 567896
rect 105892 567838 108915 567840
rect 108849 567835 108915 567838
rect 67633 567624 70226 567626
rect 67633 567568 67638 567624
rect 67694 567568 70226 567624
rect 67633 567566 70226 567568
rect 67633 567563 67699 567566
rect 108941 567354 109007 567357
rect 105892 567352 109007 567354
rect 105892 567296 108946 567352
rect 109002 567296 109007 567352
rect 105892 567294 109007 567296
rect 108941 567291 109007 567294
rect 67725 567218 67791 567221
rect 67725 567216 70042 567218
rect 67725 567160 67730 567216
rect 67786 567210 70042 567216
rect 67786 567160 70226 567210
rect 67725 567158 70226 567160
rect 67725 567155 67791 567158
rect 69982 567150 70226 567158
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 108389 566538 108455 566541
rect 105892 566536 108455 566538
rect 105892 566480 108394 566536
rect 108450 566480 108455 566536
rect 105892 566478 108455 566480
rect 108389 566475 108455 566478
rect 108941 565994 109007 565997
rect 105892 565992 109007 565994
rect 70166 565892 70226 565964
rect 105892 565936 108946 565992
rect 109002 565936 109007 565992
rect 105892 565934 109007 565936
rect 108941 565931 109007 565934
rect 67633 565858 67699 565861
rect 69982 565858 70226 565892
rect 67633 565856 70226 565858
rect 67633 565800 67638 565856
rect 67694 565832 70226 565856
rect 67694 565800 70042 565832
rect 67633 565798 70042 565800
rect 67633 565795 67699 565798
rect 108849 565178 108915 565181
rect 105892 565176 108915 565178
rect 67633 564906 67699 564909
rect 70166 564906 70226 565148
rect 105892 565120 108854 565176
rect 108910 565120 108915 565176
rect 105892 565118 108915 565120
rect 108849 565115 108915 565118
rect 67633 564904 70226 564906
rect 67633 564848 67638 564904
rect 67694 564848 70226 564904
rect 67633 564846 70226 564848
rect 67633 564843 67699 564846
rect 67541 564498 67607 564501
rect 108941 564498 109007 564501
rect 67541 564496 70042 564498
rect 67541 564440 67546 564496
rect 67602 564440 70042 564496
rect 105892 564496 109007 564498
rect 67541 564438 70042 564440
rect 67541 564435 67607 564438
rect 69982 564362 70042 564438
rect 70166 564362 70226 564468
rect 105892 564440 108946 564496
rect 109002 564440 109007 564496
rect 105892 564438 109007 564440
rect 108941 564435 109007 564438
rect 69982 564302 70226 564362
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 108941 563954 109007 563957
rect 105892 563952 109007 563954
rect 105892 563896 108946 563952
rect 109002 563896 109007 563952
rect 105892 563894 109007 563896
rect 108941 563891 109007 563894
rect 67633 563546 67699 563549
rect 70166 563546 70226 563788
rect 67633 563544 70226 563546
rect 67633 563488 67638 563544
rect 67694 563488 70226 563544
rect 67633 563486 70226 563488
rect 67633 563483 67699 563486
rect 59118 563212 59124 563276
rect 59188 563274 59194 563276
rect 59188 563214 70042 563274
rect 59188 563212 59194 563214
rect 69982 563002 70042 563214
rect 70166 563002 70226 563108
rect 105494 563004 105554 563108
rect 69982 562942 70226 563002
rect 105486 562940 105492 563004
rect 105556 562940 105562 563004
rect 67633 562322 67699 562325
rect 70166 562322 70226 562428
rect 67633 562320 70226 562322
rect 67633 562264 67638 562320
rect 67694 562264 70226 562320
rect 67633 562262 70226 562264
rect 67633 562259 67699 562262
rect 67633 562186 67699 562189
rect 67633 562184 70410 562186
rect 67633 562128 67638 562184
rect 67694 562128 70410 562184
rect 67633 562126 70410 562128
rect 67633 562123 67699 562126
rect 70350 561884 70410 562126
rect 105678 561917 105738 562428
rect 105629 561912 105738 561917
rect 105629 561856 105634 561912
rect 105690 561856 105738 561912
rect 105629 561854 105738 561856
rect 105629 561851 105695 561854
rect 108941 561098 109007 561101
rect 105892 561096 109007 561098
rect 67725 560826 67791 560829
rect 70166 560826 70226 561068
rect 105892 561040 108946 561096
rect 109002 561040 109007 561096
rect 105892 561038 109007 561040
rect 108941 561035 109007 561038
rect 67725 560824 70226 560826
rect 67725 560768 67730 560824
rect 67786 560768 70226 560824
rect 67725 560766 70226 560768
rect 67725 560763 67791 560766
rect 67633 560418 67699 560421
rect 106273 560418 106339 560421
rect 108205 560418 108271 560421
rect 67633 560416 70042 560418
rect 67633 560360 67638 560416
rect 67694 560360 70042 560416
rect 105892 560416 108271 560418
rect 67633 560358 70042 560360
rect 67633 560355 67699 560358
rect 69982 560282 70042 560358
rect 70166 560282 70226 560388
rect 105892 560360 106278 560416
rect 106334 560360 108210 560416
rect 108266 560360 108271 560416
rect 105892 560358 108271 560360
rect 106273 560355 106339 560358
rect 108205 560355 108271 560358
rect 69982 560222 70226 560282
rect 108849 559738 108915 559741
rect 105892 559736 108915 559738
rect 105892 559680 108854 559736
rect 108910 559680 108915 559736
rect 105892 559678 108915 559680
rect 108849 559675 108915 559678
rect 67633 559466 67699 559469
rect 67633 559464 70410 559466
rect 67633 559408 67638 559464
rect 67694 559408 70410 559464
rect 67633 559406 70410 559408
rect 67633 559403 67699 559406
rect 70350 559164 70410 559406
rect 108941 559058 109007 559061
rect 105892 559056 109007 559058
rect 105892 559000 108946 559056
rect 109002 559000 109007 559056
rect 105892 558998 109007 559000
rect 108941 558995 109007 558998
rect 68829 558922 68895 558925
rect 68829 558920 70226 558922
rect 68829 558864 68834 558920
rect 68890 558864 70226 558920
rect 68829 558862 70226 558864
rect 68829 558859 68895 558862
rect 70166 558484 70226 558862
rect 108941 558378 109007 558381
rect 105892 558376 109007 558378
rect 105892 558320 108946 558376
rect 109002 558320 109007 558376
rect 105892 558318 109007 558320
rect 108941 558315 109007 558318
rect 108297 557698 108363 557701
rect 105892 557696 108363 557698
rect 67633 557562 67699 557565
rect 70166 557562 70226 557668
rect 105892 557640 108302 557696
rect 108358 557640 108363 557696
rect 105892 557638 108363 557640
rect 108297 557635 108363 557638
rect 67633 557560 70226 557562
rect 67633 557504 67638 557560
rect 67694 557504 70226 557560
rect 67633 557502 70226 557504
rect 67633 557499 67699 557502
rect 65885 557426 65951 557429
rect 69974 557426 69980 557428
rect 65885 557424 69980 557426
rect 65885 557368 65890 557424
rect 65946 557368 69980 557424
rect 65885 557366 69980 557368
rect 65885 557363 65951 557366
rect 69974 557364 69980 557366
rect 70044 557364 70050 557428
rect 108941 557018 109007 557021
rect 105892 557016 109007 557018
rect 67817 556746 67883 556749
rect 70166 556746 70226 556988
rect 105892 556960 108946 557016
rect 109002 556960 109007 557016
rect 105892 556958 109007 556960
rect 108941 556955 109007 556958
rect 67817 556744 70226 556746
rect 67817 556688 67822 556744
rect 67878 556688 70226 556744
rect 67817 556686 70226 556688
rect 67817 556683 67883 556686
rect 106406 556338 106412 556340
rect 67633 556202 67699 556205
rect 70166 556202 70226 556308
rect 105892 556278 106412 556338
rect 106406 556276 106412 556278
rect 106476 556276 106482 556340
rect 67633 556200 70226 556202
rect 67633 556144 67638 556200
rect 67694 556144 70226 556200
rect 67633 556142 70226 556144
rect 67633 556139 67699 556142
rect 108941 555794 109007 555797
rect 105892 555792 109007 555794
rect 105892 555736 108946 555792
rect 109002 555736 109007 555792
rect 105892 555734 109007 555736
rect 108941 555731 109007 555734
rect 67633 555386 67699 555389
rect 70166 555386 70226 555628
rect 67633 555384 70226 555386
rect 67633 555328 67638 555384
rect 67694 555328 70226 555384
rect 67633 555326 70226 555328
rect 67633 555323 67699 555326
rect 67725 554842 67791 554845
rect 70166 554842 70226 554948
rect 67725 554840 70226 554842
rect 67725 554784 67730 554840
rect 67786 554784 70226 554840
rect 67725 554782 70226 554784
rect 67725 554779 67791 554782
rect 108849 554298 108915 554301
rect 105892 554296 108915 554298
rect -960 553890 480 553980
rect 68870 553964 68876 554028
rect 68940 554026 68946 554028
rect 70166 554026 70226 554268
rect 105892 554240 108854 554296
rect 108910 554240 108915 554296
rect 105892 554238 108915 554240
rect 108849 554235 108915 554238
rect 68940 553966 70226 554026
rect 68940 553964 68946 553966
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 108941 553618 109007 553621
rect 105892 553616 109007 553618
rect 67633 553482 67699 553485
rect 70166 553482 70226 553588
rect 105892 553560 108946 553616
rect 109002 553560 109007 553616
rect 105892 553558 109007 553560
rect 108941 553555 109007 553558
rect 67633 553480 70226 553482
rect 67633 553424 67638 553480
rect 67694 553424 70226 553480
rect 67633 553422 70226 553424
rect 67633 553419 67699 553422
rect 108941 552938 109007 552941
rect 105892 552936 109007 552938
rect 105892 552880 108946 552936
rect 109002 552880 109007 552936
rect 105892 552878 109007 552880
rect 108941 552875 109007 552878
rect 108389 552258 108455 552261
rect 105892 552256 108455 552258
rect 67633 552122 67699 552125
rect 70166 552122 70226 552228
rect 105892 552200 108394 552256
rect 108450 552200 108455 552256
rect 105892 552198 108455 552200
rect 108389 552195 108455 552198
rect 67633 552120 70226 552122
rect 67633 552064 67638 552120
rect 67694 552064 70226 552120
rect 67633 552062 70226 552064
rect 67633 552059 67699 552062
rect 107837 551578 107903 551581
rect 105892 551576 107903 551578
rect 67633 551306 67699 551309
rect 70166 551306 70226 551548
rect 105892 551520 107842 551576
rect 107898 551520 107903 551576
rect 105892 551518 107903 551520
rect 107837 551515 107903 551518
rect 67633 551304 70226 551306
rect 67633 551248 67638 551304
rect 67694 551248 70226 551304
rect 67633 551246 70226 551248
rect 67633 551243 67699 551246
rect 583520 551020 584960 551260
rect 108941 550898 109007 550901
rect 105892 550896 109007 550898
rect 68645 550762 68711 550765
rect 70166 550762 70226 550868
rect 105892 550840 108946 550896
rect 109002 550840 109007 550896
rect 105892 550838 109007 550840
rect 108941 550835 109007 550838
rect 68645 550760 70226 550762
rect 68645 550704 68650 550760
rect 68706 550704 70226 550760
rect 68645 550702 70226 550704
rect 68645 550699 68711 550702
rect 108849 550218 108915 550221
rect 105892 550216 108915 550218
rect 67633 549946 67699 549949
rect 70166 549946 70226 550188
rect 105892 550160 108854 550216
rect 108910 550160 108915 550216
rect 105892 550158 108915 550160
rect 108849 550155 108915 550158
rect 67633 549944 70226 549946
rect 67633 549888 67638 549944
rect 67694 549888 70226 549944
rect 67633 549886 70226 549888
rect 67633 549883 67699 549886
rect 61878 549476 61884 549540
rect 61948 549538 61954 549540
rect 108941 549538 109007 549541
rect 61948 549478 64890 549538
rect 105892 549536 109007 549538
rect 61948 549476 61954 549478
rect 64830 549402 64890 549478
rect 70166 549402 70226 549508
rect 105892 549480 108946 549536
rect 109002 549480 109007 549536
rect 105892 549478 109007 549480
rect 108941 549475 109007 549478
rect 64830 549342 70226 549402
rect 106917 548858 106983 548861
rect 105892 548856 106983 548858
rect 67725 548586 67791 548589
rect 70166 548586 70226 548828
rect 105892 548800 106922 548856
rect 106978 548800 106983 548856
rect 105892 548798 106983 548800
rect 106917 548795 106983 548798
rect 67725 548584 70226 548586
rect 67725 548528 67730 548584
rect 67786 548528 70226 548584
rect 67725 548526 70226 548528
rect 67725 548523 67791 548526
rect 67633 548042 67699 548045
rect 70166 548042 70226 548148
rect 67633 548040 70226 548042
rect 67633 547984 67638 548040
rect 67694 547984 70226 548040
rect 67633 547982 70226 547984
rect 67633 547979 67699 547982
rect 108941 547498 109007 547501
rect 105892 547496 109007 547498
rect 67725 547226 67791 547229
rect 70166 547226 70226 547468
rect 105892 547440 108946 547496
rect 109002 547440 109007 547496
rect 105892 547438 109007 547440
rect 108941 547435 109007 547438
rect 67725 547224 70226 547226
rect 67725 547168 67730 547224
rect 67786 547168 70226 547224
rect 67725 547166 70226 547168
rect 67725 547163 67791 547166
rect 108481 546818 108547 546821
rect 105892 546816 108547 546818
rect 67633 546546 67699 546549
rect 70166 546546 70226 546788
rect 105892 546760 108486 546816
rect 108542 546760 108547 546816
rect 105892 546758 108547 546760
rect 108481 546755 108547 546758
rect 67633 546544 70226 546546
rect 67633 546488 67638 546544
rect 67694 546488 70226 546544
rect 67633 546486 70226 546488
rect 67633 546483 67699 546486
rect 108941 546138 109007 546141
rect 105892 546136 109007 546138
rect 105892 546080 108946 546136
rect 109002 546080 109007 546136
rect 105892 546078 109007 546080
rect 108941 546075 109007 546078
rect 108941 545458 109007 545461
rect 105892 545456 109007 545458
rect 68553 545322 68619 545325
rect 69105 545322 69171 545325
rect 70166 545322 70226 545428
rect 105892 545400 108946 545456
rect 109002 545400 109007 545456
rect 105892 545398 109007 545400
rect 108941 545395 109007 545398
rect 68553 545320 70226 545322
rect 68553 545264 68558 545320
rect 68614 545264 69110 545320
rect 69166 545264 70226 545320
rect 68553 545262 70226 545264
rect 68553 545259 68619 545262
rect 69105 545259 69171 545262
rect 108849 544914 108915 544917
rect 105892 544912 108915 544914
rect 105892 544856 108854 544912
rect 108910 544856 108915 544912
rect 105892 544854 108915 544856
rect 108849 544851 108915 544854
rect 68185 544506 68251 544509
rect 70166 544506 70226 544748
rect 68185 544504 70226 544506
rect 68185 544448 68190 544504
rect 68246 544448 70226 544504
rect 68185 544446 70226 544448
rect 68185 544443 68251 544446
rect 68001 543962 68067 543965
rect 68921 543962 68987 543965
rect 70166 543962 70226 544068
rect 68001 543960 70226 543962
rect 68001 543904 68006 543960
rect 68062 543904 68926 543960
rect 68982 543904 70226 543960
rect 68001 543902 70226 543904
rect 68001 543899 68067 543902
rect 68921 543899 68987 543902
rect 105862 543829 105922 544068
rect 105862 543824 105971 543829
rect 105862 543768 105910 543824
rect 105966 543768 105971 543824
rect 105862 543766 105971 543768
rect 105905 543763 105971 543766
rect 108941 543418 109007 543421
rect 105892 543416 109007 543418
rect 67725 543146 67791 543149
rect 70166 543146 70226 543388
rect 105892 543360 108946 543416
rect 109002 543360 109007 543416
rect 105892 543358 109007 543360
rect 108941 543355 109007 543358
rect 67725 543144 70226 543146
rect 67725 543088 67730 543144
rect 67786 543088 70226 543144
rect 67725 543086 70226 543088
rect 67725 543083 67791 543086
rect 107878 542738 107884 542740
rect 67633 542602 67699 542605
rect 70166 542602 70226 542708
rect 105892 542678 107884 542738
rect 107878 542676 107884 542678
rect 107948 542676 107954 542740
rect 67633 542600 70226 542602
rect 67633 542544 67638 542600
rect 67694 542544 70226 542600
rect 67633 542542 70226 542544
rect 67633 542539 67699 542542
rect 108941 542058 109007 542061
rect 105892 542056 109007 542058
rect 69013 541786 69079 541789
rect 70166 541786 70226 542028
rect 105892 542000 108946 542056
rect 109002 542000 109007 542056
rect 105892 541998 109007 542000
rect 108941 541995 109007 541998
rect 69013 541784 70226 541786
rect 69013 541728 69018 541784
rect 69074 541728 70226 541784
rect 69013 541726 70226 541728
rect 69013 541723 69079 541726
rect 67633 541242 67699 541245
rect 70166 541242 70226 541348
rect 67633 541240 70226 541242
rect 67633 541184 67638 541240
rect 67694 541184 70226 541240
rect 67633 541182 70226 541184
rect 67633 541179 67699 541182
rect -960 540684 480 540924
rect 106273 540698 106339 540701
rect 105892 540696 106339 540698
rect 67633 540154 67699 540157
rect 70166 540154 70226 540668
rect 105892 540640 106278 540696
rect 106334 540640 106339 540696
rect 105892 540638 106339 540640
rect 106273 540635 106339 540638
rect 107469 540154 107535 540157
rect 67633 540152 70226 540154
rect 67633 540096 67638 540152
rect 67694 540096 70226 540152
rect 67633 540094 70226 540096
rect 105892 540152 107535 540154
rect 105892 540096 107474 540152
rect 107530 540096 107535 540152
rect 105892 540094 107535 540096
rect 67633 540091 67699 540094
rect 107469 540091 107535 540094
rect 56409 538114 56475 538117
rect 73889 538114 73955 538117
rect 56409 538112 73955 538114
rect 56409 538056 56414 538112
rect 56470 538056 73894 538112
rect 73950 538056 73955 538112
rect 56409 538054 73955 538056
rect 56409 538051 56475 538054
rect 73889 538051 73955 538054
rect 80329 538114 80395 538117
rect 114829 538114 114895 538117
rect 80329 538112 114895 538114
rect 80329 538056 80334 538112
rect 80390 538056 114834 538112
rect 114890 538056 114895 538112
rect 80329 538054 114895 538056
rect 80329 538051 80395 538054
rect 114829 538051 114895 538054
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 99465 537434 99531 537437
rect 107694 537434 107700 537436
rect 99465 537432 107700 537434
rect 99465 537376 99470 537432
rect 99526 537376 107700 537432
rect 99465 537374 107700 537376
rect 99465 537371 99531 537374
rect 107694 537372 107700 537374
rect 107764 537372 107770 537436
rect 69606 536828 69612 536892
rect 69676 536890 69682 536892
rect 69841 536890 69907 536893
rect 69676 536888 69907 536890
rect 69676 536832 69846 536888
rect 69902 536832 69907 536888
rect 69676 536830 69907 536832
rect 69676 536828 69682 536830
rect 69841 536827 69907 536830
rect 100937 536890 101003 536893
rect 101254 536890 101260 536892
rect 100937 536888 101260 536890
rect 100937 536832 100942 536888
rect 100998 536832 101260 536888
rect 100937 536830 101260 536832
rect 100937 536827 101003 536830
rect 101254 536828 101260 536830
rect 101324 536828 101330 536892
rect 101990 536828 101996 536892
rect 102060 536890 102066 536892
rect 105629 536890 105695 536893
rect 102060 536888 105695 536890
rect 102060 536832 105634 536888
rect 105690 536832 105695 536888
rect 102060 536830 105695 536832
rect 102060 536828 102066 536830
rect 105629 536827 105695 536830
rect 89621 534714 89687 534717
rect 115974 534714 115980 534716
rect 89621 534712 115980 534714
rect 89621 534656 89626 534712
rect 89682 534656 115980 534712
rect 89621 534654 115980 534656
rect 89621 534651 89687 534654
rect 115974 534652 115980 534654
rect 116044 534652 116050 534716
rect 98545 529138 98611 529141
rect 110822 529138 110828 529140
rect 98545 529136 110828 529138
rect 98545 529080 98550 529136
rect 98606 529080 110828 529136
rect 98545 529078 110828 529080
rect 98545 529075 98611 529078
rect 110822 529076 110828 529078
rect 110892 529076 110898 529140
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 44030 526356 44036 526420
rect 44100 526418 44106 526420
rect 77753 526418 77819 526421
rect 44100 526416 77819 526418
rect 44100 526360 77758 526416
rect 77814 526360 77819 526416
rect 44100 526358 77819 526360
rect 44100 526356 44106 526358
rect 77753 526355 77819 526358
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 137093 499626 137159 499629
rect 143574 499626 143580 499628
rect 137093 499624 143580 499626
rect 137093 499568 137098 499624
rect 137154 499568 143580 499624
rect 137093 499566 143580 499568
rect 137093 499563 137159 499566
rect 143574 499564 143580 499566
rect 143644 499564 143650 499628
rect 583520 497844 584960 498084
rect 86769 497450 86835 497453
rect 115974 497450 115980 497452
rect 86769 497448 115980 497450
rect 86769 497392 86774 497448
rect 86830 497392 115980 497448
rect 86769 497390 115980 497392
rect 86769 497387 86835 497390
rect 115974 497388 115980 497390
rect 116044 497388 116050 497452
rect 84837 496090 84903 496093
rect 111742 496090 111748 496092
rect 84837 496088 111748 496090
rect 84837 496032 84842 496088
rect 84898 496032 111748 496088
rect 84837 496030 111748 496032
rect 84837 496027 84903 496030
rect 111742 496028 111748 496030
rect 111812 496090 111818 496092
rect 117497 496090 117563 496093
rect 111812 496088 117563 496090
rect 111812 496032 117502 496088
rect 117558 496032 117563 496088
rect 111812 496030 117563 496032
rect 111812 496028 111818 496030
rect 117497 496027 117563 496030
rect 50838 493308 50844 493372
rect 50908 493370 50914 493372
rect 52310 493370 52316 493372
rect 50908 493310 52316 493370
rect 50908 493308 50914 493310
rect 52310 493308 52316 493310
rect 52380 493370 52386 493372
rect 74809 493370 74875 493373
rect 52380 493368 74875 493370
rect 52380 493312 74814 493368
rect 74870 493312 74875 493368
rect 52380 493310 74875 493312
rect 52380 493308 52386 493310
rect 74809 493307 74875 493310
rect 79317 492826 79383 492829
rect 111742 492826 111748 492828
rect 79317 492824 111748 492826
rect 79317 492768 79322 492824
rect 79378 492768 111748 492824
rect 79317 492766 111748 492768
rect 79317 492763 79383 492766
rect 111742 492764 111748 492766
rect 111812 492764 111818 492828
rect 95785 491874 95851 491877
rect 124254 491874 124260 491876
rect 95785 491872 124260 491874
rect 95785 491816 95790 491872
rect 95846 491816 124260 491872
rect 95785 491814 124260 491816
rect 95785 491811 95851 491814
rect 124254 491812 124260 491814
rect 124324 491874 124330 491876
rect 125685 491874 125751 491877
rect 124324 491872 125751 491874
rect 124324 491816 125690 491872
rect 125746 491816 125751 491872
rect 124324 491814 125751 491816
rect 124324 491812 124330 491814
rect 125685 491811 125751 491814
rect 96981 491738 97047 491741
rect 97809 491738 97875 491741
rect 99230 491738 99236 491740
rect 96981 491736 99236 491738
rect 96981 491680 96986 491736
rect 97042 491680 97814 491736
rect 97870 491680 99236 491736
rect 96981 491678 99236 491680
rect 96981 491675 97047 491678
rect 97809 491675 97875 491678
rect 99230 491676 99236 491678
rect 99300 491676 99306 491740
rect 92473 491466 92539 491469
rect 101213 491466 101279 491469
rect 92473 491464 101279 491466
rect 92473 491408 92478 491464
rect 92534 491408 101218 491464
rect 101274 491408 101279 491464
rect 92473 491406 101279 491408
rect 92473 491403 92539 491406
rect 101213 491403 101279 491406
rect 99281 491330 99347 491333
rect 111057 491330 111123 491333
rect 99281 491328 111123 491330
rect 99281 491272 99286 491328
rect 99342 491272 111062 491328
rect 111118 491272 111123 491328
rect 99281 491270 111123 491272
rect 99281 491267 99347 491270
rect 111057 491267 111123 491270
rect 97441 491194 97507 491197
rect 112437 491194 112503 491197
rect 97441 491192 112503 491194
rect 97441 491136 97446 491192
rect 97502 491136 112442 491192
rect 112498 491136 112503 491192
rect 97441 491134 112503 491136
rect 97441 491131 97507 491134
rect 112437 491131 112503 491134
rect 92565 490650 92631 490653
rect 103830 490650 103836 490652
rect 92565 490648 103836 490650
rect 92565 490592 92570 490648
rect 92626 490592 103836 490648
rect 92565 490590 103836 490592
rect 92565 490587 92631 490590
rect 103830 490588 103836 490590
rect 103900 490588 103906 490652
rect 57830 490452 57836 490516
rect 57900 490514 57906 490516
rect 87045 490514 87111 490517
rect 57900 490512 87111 490514
rect 57900 490456 87050 490512
rect 87106 490456 87111 490512
rect 57900 490454 87111 490456
rect 57900 490452 57906 490454
rect 87045 490451 87111 490454
rect 94129 490514 94195 490517
rect 94957 490514 95023 490517
rect 108982 490514 108988 490516
rect 94129 490512 108988 490514
rect 94129 490456 94134 490512
rect 94190 490456 94962 490512
rect 95018 490456 108988 490512
rect 94129 490454 108988 490456
rect 94129 490451 94195 490454
rect 94957 490451 95023 490454
rect 108982 490452 108988 490454
rect 109052 490452 109058 490516
rect 71037 489970 71103 489973
rect 69798 489968 71103 489970
rect 69798 489912 71042 489968
rect 71098 489912 71103 489968
rect 69798 489910 71103 489912
rect 53598 489092 53604 489156
rect 53668 489154 53674 489156
rect 69798 489154 69858 489910
rect 71037 489907 71103 489910
rect 53668 489094 69858 489154
rect 53668 489092 53674 489094
rect 69013 489018 69079 489021
rect 70166 489018 70226 489668
rect 102225 489290 102291 489293
rect 99790 489288 102291 489290
rect 99790 489232 102230 489288
rect 102286 489232 102291 489288
rect 99790 489230 102291 489232
rect 99790 489124 99850 489230
rect 102225 489227 102291 489230
rect 69013 489016 70226 489018
rect 69013 488960 69018 489016
rect 69074 488960 70226 489016
rect 69013 488958 70226 488960
rect 69013 488955 69079 488958
rect -960 488596 480 488836
rect 67633 488066 67699 488069
rect 70350 488066 70410 488308
rect 67633 488064 70410 488066
rect 67633 488008 67638 488064
rect 67694 488008 70410 488064
rect 67633 488006 70410 488008
rect 99606 488066 99666 488308
rect 102317 488066 102383 488069
rect 99606 488064 102383 488066
rect 99606 488008 102322 488064
rect 102378 488008 102383 488064
rect 99606 488006 102383 488008
rect 67633 488003 67699 488006
rect 102317 488003 102383 488006
rect 67633 487930 67699 487933
rect 102225 487930 102291 487933
rect 67633 487928 70226 487930
rect 67633 487872 67638 487928
rect 67694 487872 70226 487928
rect 67633 487870 70226 487872
rect 67633 487867 67699 487870
rect 70166 487764 70226 487870
rect 99790 487928 102291 487930
rect 99790 487872 102230 487928
rect 102286 487872 102291 487928
rect 99790 487870 102291 487872
rect 99790 487764 99850 487870
rect 102225 487867 102291 487870
rect 52310 487188 52316 487252
rect 52380 487250 52386 487252
rect 53649 487250 53715 487253
rect 52380 487248 53715 487250
rect 52380 487192 53654 487248
rect 53710 487192 53715 487248
rect 52380 487190 53715 487192
rect 52380 487188 52386 487190
rect 53649 487187 53715 487190
rect 68001 486706 68067 486709
rect 69054 486706 69060 486708
rect 68001 486704 69060 486706
rect 68001 486648 68006 486704
rect 68062 486648 69060 486704
rect 68001 486646 69060 486648
rect 68001 486643 68067 486646
rect 69054 486644 69060 486646
rect 69124 486706 69130 486708
rect 70350 486706 70410 486948
rect 69124 486646 70410 486706
rect 99422 486709 99482 486948
rect 99422 486704 99531 486709
rect 102225 486706 102291 486709
rect 99422 486648 99470 486704
rect 99526 486648 99531 486704
rect 99422 486646 99531 486648
rect 69124 486644 69130 486646
rect 99465 486643 99531 486646
rect 99790 486704 102291 486706
rect 99790 486648 102230 486704
rect 102286 486648 102291 486704
rect 99790 486646 102291 486648
rect 99790 486404 99850 486646
rect 102225 486643 102291 486646
rect 103513 486434 103579 486437
rect 110638 486434 110644 486436
rect 103513 486432 110644 486434
rect 103513 486376 103518 486432
rect 103574 486376 110644 486432
rect 103513 486374 110644 486376
rect 103513 486371 103579 486374
rect 110638 486372 110644 486374
rect 110708 486434 110714 486436
rect 122046 486434 122052 486436
rect 110708 486374 122052 486434
rect 110708 486372 110714 486374
rect 122046 486372 122052 486374
rect 122116 486372 122122 486436
rect 70166 486026 70226 486268
rect 67774 485966 70226 486026
rect 67774 485890 67834 485966
rect 69841 485892 69907 485893
rect 67590 485830 67834 485890
rect 39798 485692 39804 485756
rect 39868 485754 39874 485756
rect 66989 485754 67055 485757
rect 67590 485754 67650 485830
rect 69790 485828 69796 485892
rect 69860 485890 69907 485892
rect 69860 485888 69952 485890
rect 69902 485832 69952 485888
rect 69860 485830 69952 485832
rect 69860 485828 69907 485830
rect 69841 485827 69907 485828
rect 39868 485752 67650 485754
rect 39868 485696 66994 485752
rect 67050 485696 67650 485752
rect 99790 485754 100034 485790
rect 103421 485754 103487 485757
rect 99790 485752 103487 485754
rect 99790 485730 103426 485752
rect 99790 485724 99850 485730
rect 39868 485694 67650 485696
rect 99974 485696 103426 485730
rect 103482 485696 103487 485752
rect 99974 485694 103487 485696
rect 39868 485692 39874 485694
rect 66989 485691 67055 485694
rect 103421 485691 103487 485694
rect 67633 485210 67699 485213
rect 70166 485210 70226 485588
rect 103421 485210 103487 485213
rect 67633 485208 70226 485210
rect 67633 485152 67638 485208
rect 67694 485152 70226 485208
rect 67633 485150 70226 485152
rect 99790 485208 103487 485210
rect 99790 485152 103426 485208
rect 103482 485152 103487 485208
rect 99790 485150 103487 485152
rect 67633 485147 67699 485150
rect 99790 485044 99850 485150
rect 103421 485147 103487 485150
rect 111977 485074 112043 485077
rect 113030 485074 113036 485076
rect 111977 485072 113036 485074
rect 111977 485016 111982 485072
rect 112038 485016 113036 485072
rect 111977 485014 113036 485016
rect 111977 485011 112043 485014
rect 113030 485012 113036 485014
rect 113100 485074 113106 485076
rect 131113 485074 131179 485077
rect 113100 485072 131179 485074
rect 113100 485016 131118 485072
rect 131174 485016 131179 485072
rect 113100 485014 131179 485016
rect 113100 485012 113106 485014
rect 131113 485011 131179 485014
rect 65926 484604 65932 484668
rect 65996 484666 66002 484668
rect 70166 484666 70226 484908
rect 70342 484666 70348 484668
rect 65996 484606 70348 484666
rect 65996 484604 66002 484606
rect 70342 484604 70348 484606
rect 70412 484604 70418 484668
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 99414 484468 99420 484532
rect 99484 484530 99490 484532
rect 100109 484530 100175 484533
rect 99484 484528 100175 484530
rect 99484 484472 100114 484528
rect 100170 484472 100175 484528
rect 583520 484516 584960 484606
rect 99484 484470 100175 484472
rect 99484 484468 99490 484470
rect 100109 484467 100175 484470
rect 67633 483714 67699 483717
rect 70166 483714 70226 484228
rect 103421 483850 103487 483853
rect 67633 483712 70226 483714
rect 67633 483656 67638 483712
rect 67694 483656 70226 483712
rect 99790 483848 103487 483850
rect 99790 483792 103426 483848
rect 103482 483792 103487 483848
rect 99790 483790 103487 483792
rect 99790 483684 99850 483790
rect 103421 483787 103487 483790
rect 67633 483654 70226 483656
rect 67633 483651 67699 483654
rect 123385 483170 123451 483173
rect 124070 483170 124076 483172
rect 123385 483168 124076 483170
rect 123385 483112 123390 483168
rect 123446 483112 124076 483168
rect 123385 483110 124076 483112
rect 123385 483107 123451 483110
rect 124070 483108 124076 483110
rect 124140 483108 124146 483172
rect 69841 482626 69907 482629
rect 70350 482626 70410 482868
rect 69841 482624 70410 482626
rect 69841 482568 69846 482624
rect 69902 482568 70410 482624
rect 69841 482566 70410 482568
rect 99790 482626 99850 482868
rect 103329 482626 103395 482629
rect 99790 482624 103395 482626
rect 99790 482568 103334 482624
rect 103390 482568 103395 482624
rect 99790 482566 103395 482568
rect 69841 482563 69907 482566
rect 103329 482563 103395 482566
rect 68093 482490 68159 482493
rect 69197 482490 69263 482493
rect 103421 482490 103487 482493
rect 68093 482488 70226 482490
rect 68093 482432 68098 482488
rect 68154 482432 69202 482488
rect 69258 482432 70226 482488
rect 68093 482430 70226 482432
rect 68093 482427 68159 482430
rect 69197 482427 69263 482430
rect 70166 482324 70226 482430
rect 99790 482488 103487 482490
rect 99790 482432 103426 482488
rect 103482 482432 103487 482488
rect 99790 482430 103487 482432
rect 99790 482324 99850 482430
rect 103421 482427 103487 482430
rect 114553 482356 114619 482357
rect 114502 482292 114508 482356
rect 114572 482354 114619 482356
rect 114572 482352 114664 482354
rect 114614 482296 114664 482352
rect 114572 482294 114664 482296
rect 114572 482292 114619 482294
rect 114553 482291 114619 482292
rect 69982 481750 70226 481810
rect 67449 481672 67515 481677
rect 67449 481616 67454 481672
rect 67510 481616 67515 481672
rect 67449 481611 67515 481616
rect 67452 481266 67512 481611
rect 69105 481538 69171 481541
rect 69982 481538 70042 481750
rect 70166 481644 70226 481750
rect 99790 481750 100034 481810
rect 99790 481644 99850 481750
rect 69105 481536 70042 481538
rect 69105 481480 69110 481536
rect 69166 481480 70042 481536
rect 69105 481478 70042 481480
rect 99974 481538 100034 481750
rect 103421 481538 103487 481541
rect 99974 481536 103487 481538
rect 99974 481480 103426 481536
rect 103482 481480 103487 481536
rect 99974 481478 103487 481480
rect 69105 481475 69171 481478
rect 103421 481475 103487 481478
rect 103329 481266 103395 481269
rect 67452 481206 70226 481266
rect 70166 480964 70226 481206
rect 99790 481264 103395 481266
rect 99790 481208 103334 481264
rect 103390 481208 103395 481264
rect 99790 481206 103395 481208
rect 99790 480964 99850 481206
rect 103329 481203 103395 481206
rect 113030 480796 113036 480860
rect 113100 480858 113106 480860
rect 117681 480858 117747 480861
rect 113100 480856 117747 480858
rect 113100 480800 117686 480856
rect 117742 480800 117747 480856
rect 113100 480798 117747 480800
rect 113100 480796 113106 480798
rect 117681 480795 117747 480798
rect 67633 479906 67699 479909
rect 70350 479906 70410 480148
rect 67633 479904 70410 479906
rect 67633 479848 67638 479904
rect 67694 479848 70410 479904
rect 67633 479846 70410 479848
rect 99790 479906 99850 480148
rect 103421 479906 103487 479909
rect 99790 479904 103487 479906
rect 99790 479848 103426 479904
rect 103482 479848 103487 479904
rect 99790 479846 103487 479848
rect 67633 479843 67699 479846
rect 103421 479843 103487 479846
rect 103329 479770 103395 479773
rect 99790 479768 103395 479770
rect 99790 479712 103334 479768
rect 103390 479712 103395 479768
rect 99790 479710 103395 479712
rect 99790 479604 99850 479710
rect 103329 479707 103395 479710
rect 70166 479090 70226 479468
rect 66118 479030 70226 479090
rect 65793 478954 65859 478957
rect 66118 478956 66178 479030
rect 66110 478954 66116 478956
rect 65793 478952 66116 478954
rect 65793 478896 65798 478952
rect 65854 478896 66116 478952
rect 65793 478894 66116 478896
rect 65793 478891 65859 478894
rect 66110 478892 66116 478894
rect 66180 478892 66186 478956
rect 67265 478546 67331 478549
rect 70350 478546 70410 478788
rect 67265 478544 70410 478546
rect 67265 478488 67270 478544
rect 67326 478488 70410 478544
rect 67265 478486 70410 478488
rect 67265 478483 67331 478486
rect 99790 477730 99850 478108
rect 103421 477730 103487 477733
rect 99790 477728 103487 477730
rect 99790 477672 103426 477728
rect 103482 477672 103487 477728
rect 99790 477670 103487 477672
rect 103421 477667 103487 477670
rect 63125 477458 63191 477461
rect 64638 477458 64644 477460
rect 63125 477456 64644 477458
rect 63125 477400 63130 477456
rect 63186 477400 64644 477456
rect 63125 477398 64644 477400
rect 63125 477395 63191 477398
rect 64638 477396 64644 477398
rect 64708 477458 64714 477460
rect 67725 477458 67791 477461
rect 64708 477456 67791 477458
rect 64708 477400 67730 477456
rect 67786 477400 67791 477456
rect 64708 477398 67791 477400
rect 64708 477396 64714 477398
rect 67725 477395 67791 477398
rect 68737 477052 68803 477053
rect 68686 477050 68692 477052
rect 68610 476990 68692 477050
rect 68756 477050 68803 477052
rect 70166 477050 70226 477428
rect 68756 477048 70226 477050
rect 68798 476992 70226 477048
rect 68686 476988 68692 476990
rect 68756 476990 70226 476992
rect 99790 477050 99850 477428
rect 103237 477050 103303 477053
rect 99790 477048 103303 477050
rect 99790 476992 103242 477048
rect 103298 476992 103303 477048
rect 99790 476990 103303 476992
rect 68756 476988 68803 476990
rect 68737 476987 68803 476988
rect 103237 476987 103303 476990
rect 99790 476778 100034 476812
rect 105169 476778 105235 476781
rect 99790 476776 105235 476778
rect 99790 476752 105174 476776
rect 99790 476748 99850 476752
rect 67633 476370 67699 476373
rect 70534 476370 70594 476748
rect 99974 476720 105174 476752
rect 105230 476720 105235 476776
rect 99974 476718 105235 476720
rect 105169 476715 105235 476718
rect 103329 476506 103395 476509
rect 67633 476368 70594 476370
rect 67633 476312 67638 476368
rect 67694 476312 70594 476368
rect 67633 476310 70594 476312
rect 99790 476504 103395 476506
rect 99790 476448 103334 476504
rect 103390 476448 103395 476504
rect 99790 476446 103395 476448
rect 67633 476307 67699 476310
rect 67725 476234 67791 476237
rect 67725 476232 70042 476234
rect 67725 476176 67730 476232
rect 67786 476176 70042 476232
rect 99790 476204 99850 476446
rect 103329 476443 103395 476446
rect 67725 476174 70042 476176
rect 67725 476171 67791 476174
rect 69982 476130 70042 476174
rect 69982 476070 70226 476130
rect 70166 476068 70226 476070
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 67633 475690 67699 475693
rect 102225 475690 102291 475693
rect 67633 475688 70226 475690
rect 67633 475632 67638 475688
rect 67694 475632 70226 475688
rect 67633 475630 70226 475632
rect 67633 475627 67699 475630
rect 70166 475524 70226 475630
rect 99790 475688 102291 475690
rect 99790 475632 102230 475688
rect 102286 475632 102291 475688
rect 99790 475630 102291 475632
rect 99790 475524 99850 475630
rect 102225 475627 102291 475630
rect 67725 475146 67791 475149
rect 102317 475146 102383 475149
rect 67725 475144 70226 475146
rect 67725 475088 67730 475144
rect 67786 475088 70226 475144
rect 67725 475086 70226 475088
rect 67725 475083 67791 475086
rect 70166 474844 70226 475086
rect 99790 475144 102383 475146
rect 99790 475088 102322 475144
rect 102378 475088 102383 475144
rect 99790 475086 102383 475088
rect 99790 474844 99850 475086
rect 102317 475083 102383 475086
rect 103421 474738 103487 474741
rect 104934 474738 104940 474740
rect 103421 474736 104940 474738
rect 103421 474680 103426 474736
rect 103482 474680 104940 474736
rect 103421 474678 104940 474680
rect 103421 474675 103487 474678
rect 104934 474676 104940 474678
rect 105004 474676 105010 474740
rect 105486 474676 105492 474740
rect 105556 474738 105562 474740
rect 110822 474738 110828 474740
rect 105556 474678 110828 474738
rect 105556 474676 105562 474678
rect 110822 474676 110828 474678
rect 110892 474676 110898 474740
rect 65977 474330 66043 474333
rect 66110 474330 66116 474332
rect 65977 474328 66116 474330
rect 65977 474272 65982 474328
rect 66038 474272 66116 474328
rect 65977 474270 66116 474272
rect 65977 474267 66043 474270
rect 66110 474268 66116 474270
rect 66180 474268 66186 474332
rect 67633 474330 67699 474333
rect 102225 474330 102291 474333
rect 67633 474328 70226 474330
rect 67633 474272 67638 474328
rect 67694 474272 70226 474328
rect 67633 474270 70226 474272
rect 67633 474267 67699 474270
rect 70166 474164 70226 474270
rect 99790 474328 102291 474330
rect 99790 474272 102230 474328
rect 102286 474272 102291 474328
rect 99790 474270 102291 474272
rect 99790 474164 99850 474270
rect 102225 474267 102291 474270
rect 64830 473590 70226 473650
rect 53833 473242 53899 473245
rect 55070 473242 55076 473244
rect 53833 473240 55076 473242
rect 53833 473184 53838 473240
rect 53894 473184 55076 473240
rect 53833 473182 55076 473184
rect 53833 473179 53899 473182
rect 55070 473180 55076 473182
rect 55140 473242 55146 473244
rect 64830 473242 64890 473590
rect 70166 473484 70226 473590
rect 55140 473182 64890 473242
rect 55140 473180 55146 473182
rect 102225 472970 102291 472973
rect 99790 472968 102291 472970
rect 99790 472912 102230 472968
rect 102286 472912 102291 472968
rect 99790 472910 102291 472912
rect 99790 472804 99850 472910
rect 102225 472907 102291 472910
rect 67633 472698 67699 472701
rect 67633 472696 70226 472698
rect 67633 472640 67638 472696
rect 67694 472640 70226 472696
rect 67633 472638 70226 472640
rect 67633 472635 67699 472638
rect 70166 472124 70226 472638
rect 102225 472290 102291 472293
rect 99790 472288 102291 472290
rect 99790 472232 102230 472288
rect 102286 472232 102291 472288
rect 99790 472230 102291 472232
rect 99790 472124 99850 472230
rect 102225 472227 102291 472230
rect 62982 471548 62988 471612
rect 63052 471610 63058 471612
rect 63052 471550 70226 471610
rect 63052 471548 63058 471550
rect 70166 471444 70226 471550
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 61694 471276 61700 471340
rect 61764 471338 61770 471340
rect 62982 471338 62988 471340
rect 61764 471278 62988 471338
rect 61764 471276 61770 471278
rect 62982 471276 62988 471278
rect 63052 471276 63058 471340
rect 583520 471324 584960 471414
rect 67633 470930 67699 470933
rect 99790 470930 99850 471308
rect 102225 470930 102291 470933
rect 67633 470928 70226 470930
rect 67633 470872 67638 470928
rect 67694 470872 70226 470928
rect 67633 470870 70226 470872
rect 99790 470928 102291 470930
rect 99790 470872 102230 470928
rect 102286 470872 102291 470928
rect 99790 470870 102291 470872
rect 67633 470867 67699 470870
rect 70166 470764 70226 470870
rect 102225 470867 102291 470870
rect 102317 470658 102383 470661
rect 99974 470656 102383 470658
rect 99790 470610 99850 470628
rect 99974 470610 102322 470656
rect 99790 470600 102322 470610
rect 102378 470600 102383 470656
rect 99790 470598 102383 470600
rect 99790 470550 100034 470598
rect 102317 470595 102383 470598
rect 67725 470386 67791 470389
rect 67725 470384 70226 470386
rect 67725 470328 67730 470384
rect 67786 470328 70226 470384
rect 67725 470326 70226 470328
rect 67725 470323 67791 470326
rect 70166 470084 70226 470326
rect 102225 470250 102291 470253
rect 99790 470248 102291 470250
rect 99790 470192 102230 470248
rect 102286 470192 102291 470248
rect 99790 470190 102291 470192
rect 99790 470084 99850 470190
rect 102225 470187 102291 470190
rect 67633 469570 67699 469573
rect 102225 469570 102291 469573
rect 67633 469568 70226 469570
rect 67633 469512 67638 469568
rect 67694 469512 70226 469568
rect 67633 469510 70226 469512
rect 67633 469507 67699 469510
rect 70166 469404 70226 469510
rect 99790 469568 102291 469570
rect 99790 469512 102230 469568
rect 102286 469512 102291 469568
rect 99790 469510 102291 469512
rect 99790 469404 99850 469510
rect 102225 469507 102291 469510
rect 103605 469026 103671 469029
rect 99790 469024 103671 469026
rect 99790 468968 103610 469024
rect 103666 468968 103671 469024
rect 99790 468966 103671 468968
rect 99790 468724 99850 468966
rect 103605 468963 103671 468966
rect 67633 468210 67699 468213
rect 70166 468210 70226 468588
rect 67633 468208 70226 468210
rect 67633 468152 67638 468208
rect 67694 468152 70226 468208
rect 67633 468150 70226 468152
rect 67633 468147 67699 468150
rect 62982 467876 62988 467940
rect 63052 467938 63058 467940
rect 66069 467938 66135 467941
rect 63052 467936 69858 467938
rect 63052 467880 66074 467936
rect 66130 467880 69858 467936
rect 63052 467878 69858 467880
rect 63052 467876 63058 467878
rect 66069 467875 66135 467878
rect 69798 467666 69858 467878
rect 70350 467666 70410 467908
rect 69798 467606 70410 467666
rect 99790 466986 99850 467228
rect 102225 466986 102291 466989
rect 99790 466984 102291 466986
rect 99790 466928 102230 466984
rect 102286 466928 102291 466984
rect 99790 466926 102291 466928
rect 102225 466923 102291 466926
rect 67449 466850 67515 466853
rect 103605 466850 103671 466853
rect 67449 466848 70226 466850
rect 67449 466792 67454 466848
rect 67510 466792 70226 466848
rect 67449 466790 70226 466792
rect 67449 466787 67515 466790
rect 70166 466684 70226 466790
rect 99790 466848 103671 466850
rect 99790 466792 103610 466848
rect 103666 466792 103671 466848
rect 99790 466790 103671 466792
rect 99790 466684 99850 466790
rect 103605 466787 103671 466790
rect 102225 466170 102291 466173
rect 99790 466168 102291 466170
rect 99790 466112 102230 466168
rect 102286 466112 102291 466168
rect 99790 466110 102291 466112
rect 99790 466004 99850 466110
rect 102225 466107 102291 466110
rect 67633 465626 67699 465629
rect 70350 465626 70410 465868
rect 102317 465626 102383 465629
rect 67633 465624 70410 465626
rect 67633 465568 67638 465624
rect 67694 465568 70410 465624
rect 67633 465566 70410 465568
rect 99790 465624 102383 465626
rect 99790 465568 102322 465624
rect 102378 465568 102383 465624
rect 99790 465566 102383 465568
rect 67633 465563 67699 465566
rect 67909 465490 67975 465493
rect 67909 465488 70226 465490
rect 67909 465432 67914 465488
rect 67970 465432 70226 465488
rect 67909 465430 70226 465432
rect 67909 465427 67975 465430
rect 70166 465324 70226 465430
rect 99790 465324 99850 465566
rect 102317 465563 102383 465566
rect 102225 464810 102291 464813
rect 99790 464808 102291 464810
rect 99790 464752 102230 464808
rect 102286 464752 102291 464808
rect 99790 464750 102291 464752
rect 99790 464644 99850 464750
rect 102225 464747 102291 464750
rect 67633 464266 67699 464269
rect 70350 464266 70410 464508
rect 103329 464266 103395 464269
rect 106406 464266 106412 464268
rect 67633 464264 70410 464266
rect 67633 464208 67638 464264
rect 67694 464208 70410 464264
rect 67633 464206 70410 464208
rect 99790 464264 106412 464266
rect 99790 464208 103334 464264
rect 103390 464208 106412 464264
rect 99790 464206 106412 464208
rect 67633 464203 67699 464206
rect 64830 464070 70226 464130
rect 59118 463796 59124 463860
rect 59188 463858 59194 463860
rect 64830 463858 64890 464070
rect 70166 463964 70226 464070
rect 99790 463964 99850 464206
rect 103329 464203 103395 464206
rect 106406 464204 106412 464206
rect 106476 464204 106482 464268
rect 59188 463798 64890 463858
rect 59188 463796 59194 463798
rect 60365 463586 60431 463589
rect 60590 463586 60596 463588
rect 60365 463584 60596 463586
rect 60365 463528 60370 463584
rect 60426 463528 60596 463584
rect 60365 463526 60596 463528
rect 60365 463523 60431 463526
rect 60590 463524 60596 463526
rect 60660 463524 60666 463588
rect 67633 463450 67699 463453
rect 102225 463450 102291 463453
rect 67633 463448 70226 463450
rect 67633 463392 67638 463448
rect 67694 463392 70226 463448
rect 67633 463390 70226 463392
rect 67633 463387 67699 463390
rect 70166 463284 70226 463390
rect 99790 463448 102291 463450
rect 99790 463392 102230 463448
rect 102286 463392 102291 463448
rect 99790 463390 102291 463392
rect 99790 463284 99850 463390
rect 102225 463387 102291 463390
rect 60590 462844 60596 462908
rect 60660 462906 60666 462908
rect 60660 462846 70226 462906
rect 60660 462844 60666 462846
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect 70166 462604 70226 462846
rect 106774 462844 106780 462908
rect 106844 462906 106850 462908
rect 121729 462906 121795 462909
rect 106844 462904 121795 462906
rect 106844 462848 121734 462904
rect 121790 462848 121795 462904
rect 106844 462846 121795 462848
rect 106844 462844 106850 462846
rect 121729 462843 121795 462846
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 140773 462362 140839 462365
rect 142061 462362 142127 462365
rect 146518 462362 146524 462364
rect 140773 462360 146524 462362
rect 140773 462304 140778 462360
rect 140834 462304 142066 462360
rect 142122 462304 146524 462360
rect 140773 462302 146524 462304
rect 140773 462299 140839 462302
rect 142061 462299 142127 462302
rect 146518 462300 146524 462302
rect 146588 462300 146594 462364
rect 102317 462090 102383 462093
rect 99790 462088 102383 462090
rect 99790 462032 102322 462088
rect 102378 462032 102383 462088
rect 99790 462030 102383 462032
rect 99790 461924 99850 462030
rect 102317 462027 102383 462030
rect 67633 461546 67699 461549
rect 102225 461546 102291 461549
rect 67633 461544 70226 461546
rect 67633 461488 67638 461544
rect 67694 461488 70226 461544
rect 67633 461486 70226 461488
rect 67633 461483 67699 461486
rect 70166 461244 70226 461486
rect 99606 461544 102291 461546
rect 99606 461488 102230 461544
rect 102286 461488 102291 461544
rect 99606 461486 102291 461488
rect 99606 461244 99666 461486
rect 102225 461483 102291 461486
rect 102409 460730 102475 460733
rect 99790 460728 102475 460730
rect 99790 460672 102414 460728
rect 102470 460672 102475 460728
rect 99790 460670 102475 460672
rect 99790 460564 99850 460670
rect 102409 460667 102475 460670
rect 67633 460186 67699 460189
rect 70350 460186 70410 460428
rect 102225 460186 102291 460189
rect 67633 460184 70410 460186
rect 67633 460128 67638 460184
rect 67694 460128 70410 460184
rect 67633 460126 70410 460128
rect 99606 460184 102291 460186
rect 99606 460128 102230 460184
rect 102286 460128 102291 460184
rect 99606 460126 102291 460128
rect 67633 460123 67699 460126
rect 67633 460050 67699 460053
rect 67633 460048 70226 460050
rect 67633 459992 67638 460048
rect 67694 459992 70226 460048
rect 67633 459990 70226 459992
rect 67633 459987 67699 459990
rect 70166 459884 70226 459990
rect 99606 459884 99666 460126
rect 102225 460123 102291 460126
rect 111701 459644 111767 459645
rect 111701 459642 111748 459644
rect 111656 459640 111748 459642
rect 111656 459584 111706 459640
rect 111656 459582 111748 459584
rect 111701 459580 111748 459582
rect 111812 459580 111818 459644
rect 111701 459579 111767 459580
rect 67725 459506 67791 459509
rect 67725 459504 70226 459506
rect 67725 459448 67730 459504
rect 67786 459448 70226 459504
rect 67725 459446 70226 459448
rect 67725 459443 67791 459446
rect 70166 459204 70226 459446
rect 102225 459370 102291 459373
rect 99790 459368 102291 459370
rect 99790 459312 102230 459368
rect 102286 459312 102291 459368
rect 99790 459310 102291 459312
rect 99790 459204 99850 459310
rect 102225 459307 102291 459310
rect 67633 458826 67699 458829
rect 102317 458826 102383 458829
rect 67633 458824 70226 458826
rect 67633 458768 67638 458824
rect 67694 458768 70226 458824
rect 67633 458766 70226 458768
rect 67633 458763 67699 458766
rect 70166 458524 70226 458766
rect 99790 458824 102383 458826
rect 99790 458768 102322 458824
rect 102378 458768 102383 458824
rect 99790 458766 102383 458768
rect 99790 458524 99850 458766
rect 102317 458763 102383 458766
rect 103605 458146 103671 458149
rect 99790 458144 103671 458146
rect 99790 458088 103610 458144
rect 103666 458088 103671 458144
rect 99790 458086 103671 458088
rect 67633 458010 67699 458013
rect 67633 458008 70226 458010
rect 67633 457952 67638 458008
rect 67694 457952 70226 458008
rect 67633 457950 70226 457952
rect 67633 457947 67699 457950
rect 70166 457844 70226 457950
rect 99790 457844 99850 458086
rect 103605 458083 103671 458086
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 67725 457466 67791 457469
rect 67725 457464 70226 457466
rect 67725 457408 67730 457464
rect 67786 457408 70226 457464
rect 67725 457406 70226 457408
rect 67725 457403 67791 457406
rect 70166 457164 70226 457406
rect 102317 456650 102383 456653
rect 99790 456648 102383 456650
rect 99790 456592 102322 456648
rect 102378 456592 102383 456648
rect 99790 456590 102383 456592
rect 99790 456484 99850 456590
rect 102317 456587 102383 456590
rect 102225 456106 102291 456109
rect 99790 456104 102291 456106
rect 99790 456048 102230 456104
rect 102286 456048 102291 456104
rect 99790 456046 102291 456048
rect 67633 455970 67699 455973
rect 67633 455968 70226 455970
rect 67633 455912 67638 455968
rect 67694 455912 70226 455968
rect 67633 455910 70226 455912
rect 67633 455907 67699 455910
rect 70166 455804 70226 455910
rect 99790 455804 99850 456046
rect 102225 456043 102291 456046
rect 102225 455290 102291 455293
rect 99790 455288 102291 455290
rect 99790 455232 102230 455288
rect 102286 455232 102291 455288
rect 99790 455230 102291 455232
rect 99790 455124 99850 455230
rect 102225 455227 102291 455230
rect 67633 454610 67699 454613
rect 70166 454610 70226 454988
rect 102317 454746 102383 454749
rect 67633 454608 70226 454610
rect 67633 454552 67638 454608
rect 67694 454552 70226 454608
rect 67633 454550 70226 454552
rect 99790 454744 102383 454746
rect 99790 454688 102322 454744
rect 102378 454688 102383 454744
rect 99790 454686 102383 454688
rect 67633 454547 67699 454550
rect 99790 454444 99850 454686
rect 102317 454683 102383 454686
rect 68502 454004 68508 454068
rect 68572 454066 68578 454068
rect 68870 454066 68876 454068
rect 68572 454006 68876 454066
rect 68572 454004 68578 454006
rect 68870 454004 68876 454006
rect 68940 454066 68946 454068
rect 70166 454066 70226 454308
rect 68940 454006 70226 454066
rect 68940 454004 68946 454006
rect 102225 453930 102291 453933
rect 99790 453928 102291 453930
rect 99790 453872 102230 453928
rect 102286 453872 102291 453928
rect 99790 453870 102291 453872
rect 99790 453764 99850 453870
rect 102225 453867 102291 453870
rect 125777 453930 125843 453933
rect 126830 453930 126836 453932
rect 125777 453928 126836 453930
rect 125777 453872 125782 453928
rect 125838 453872 126836 453928
rect 125777 453870 126836 453872
rect 125777 453867 125843 453870
rect 126830 453868 126836 453870
rect 126900 453868 126906 453932
rect 67725 453250 67791 453253
rect 70166 453250 70226 453628
rect 102317 453386 102383 453389
rect 67725 453248 70226 453250
rect 67725 453192 67730 453248
rect 67786 453192 70226 453248
rect 67725 453190 70226 453192
rect 99790 453384 102383 453386
rect 99790 453328 102322 453384
rect 102378 453328 102383 453384
rect 99790 453326 102383 453328
rect 67725 453187 67791 453190
rect 99790 453084 99850 453326
rect 102317 453323 102383 453326
rect 67633 452706 67699 452709
rect 70350 452706 70410 452948
rect 67633 452704 70410 452706
rect 67633 452648 67638 452704
rect 67694 452648 70410 452704
rect 67633 452646 70410 452648
rect 67633 452643 67699 452646
rect 102225 452570 102291 452573
rect 99790 452568 102291 452570
rect 99790 452512 102230 452568
rect 102286 452512 102291 452568
rect 99790 452510 102291 452512
rect 99790 452404 99850 452510
rect 102225 452507 102291 452510
rect 67633 451890 67699 451893
rect 70166 451890 70226 452268
rect 67633 451888 70226 451890
rect 67633 451832 67638 451888
rect 67694 451832 70226 451888
rect 67633 451830 70226 451832
rect 67633 451827 67699 451830
rect 68737 451346 68803 451349
rect 70350 451346 70410 451588
rect 68737 451344 70410 451346
rect 68737 451288 68742 451344
rect 68798 451288 70410 451344
rect 68737 451286 70410 451288
rect 106273 451346 106339 451349
rect 107878 451346 107884 451348
rect 106273 451344 107884 451346
rect 106273 451288 106278 451344
rect 106334 451288 107884 451344
rect 106273 451286 107884 451288
rect 68737 451283 68803 451286
rect 106273 451283 106339 451286
rect 107878 451284 107884 451286
rect 107948 451284 107954 451348
rect 67633 450802 67699 450805
rect 67633 450800 70226 450802
rect 67633 450744 67638 450800
rect 67694 450744 70226 450800
rect 67633 450742 70226 450744
rect 67633 450739 67699 450742
rect 70166 450364 70226 450742
rect 99790 450666 99850 450908
rect 102225 450666 102291 450669
rect 99790 450664 102291 450666
rect 99790 450608 102230 450664
rect 102286 450608 102291 450664
rect 99790 450606 102291 450608
rect 102225 450603 102291 450606
rect 102777 450530 102843 450533
rect 99790 450528 102843 450530
rect 99790 450472 102782 450528
rect 102838 450472 102843 450528
rect 99790 450470 102843 450472
rect 99790 450364 99850 450470
rect 102777 450467 102843 450470
rect 106273 449986 106339 449989
rect 141918 449986 141924 449988
rect 103470 449984 141924 449986
rect 103470 449928 106278 449984
rect 106334 449928 141924 449984
rect 103470 449926 141924 449928
rect 61878 449788 61884 449852
rect 61948 449850 61954 449852
rect 103470 449850 103530 449926
rect 106273 449923 106339 449926
rect 141918 449924 141924 449926
rect 141988 449924 141994 449988
rect 61948 449790 70226 449850
rect 61948 449788 61954 449790
rect 70166 449684 70226 449790
rect 99790 449790 103530 449850
rect 99790 449684 99850 449790
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 61745 448626 61811 448629
rect 61878 448626 61884 448628
rect 61745 448624 61884 448626
rect 61745 448568 61750 448624
rect 61806 448568 61884 448624
rect 61745 448566 61884 448568
rect 61745 448563 61811 448566
rect 61878 448564 61884 448566
rect 61948 448564 61954 448628
rect 67817 448626 67883 448629
rect 70166 448626 70226 448868
rect 67817 448624 70226 448626
rect 67817 448568 67822 448624
rect 67878 448568 70226 448624
rect 67817 448566 70226 448568
rect 99606 448626 99666 448868
rect 102225 448626 102291 448629
rect 99606 448624 102291 448626
rect 99606 448568 102230 448624
rect 102286 448568 102291 448624
rect 99606 448566 102291 448568
rect 67817 448563 67883 448566
rect 102225 448563 102291 448566
rect 102225 448490 102291 448493
rect 99790 448488 102291 448490
rect 99790 448432 102230 448488
rect 102286 448432 102291 448488
rect 99790 448430 102291 448432
rect 99790 448324 99850 448430
rect 102225 448427 102291 448430
rect 52269 447810 52335 447813
rect 64638 447810 64644 447812
rect 52269 447808 64644 447810
rect 52269 447752 52274 447808
rect 52330 447752 64644 447808
rect 52269 447750 64644 447752
rect 52269 447747 52335 447750
rect 64638 447748 64644 447750
rect 64708 447810 64714 447812
rect 70166 447810 70226 448188
rect 102317 447946 102383 447949
rect 64708 447750 70226 447810
rect 99790 447944 102383 447946
rect 99790 447888 102322 447944
rect 102378 447888 102383 447944
rect 99790 447886 102383 447888
rect 64708 447748 64714 447750
rect 99790 447644 99850 447886
rect 102317 447883 102383 447886
rect 67633 447266 67699 447269
rect 70350 447266 70410 447508
rect 67633 447264 70410 447266
rect 67633 447208 67638 447264
rect 67694 447208 70410 447264
rect 67633 447206 70410 447208
rect 67633 447203 67699 447206
rect 67725 446450 67791 446453
rect 70166 446450 70226 446828
rect 99606 446586 99666 446828
rect 101990 446586 101996 446588
rect 99606 446526 101996 446586
rect 101990 446524 101996 446526
rect 102060 446586 102066 446588
rect 102317 446586 102383 446589
rect 102060 446584 102383 446586
rect 102060 446528 102322 446584
rect 102378 446528 102383 446584
rect 102060 446526 102383 446528
rect 102060 446524 102066 446526
rect 102317 446523 102383 446526
rect 67725 446448 70226 446450
rect 67725 446392 67730 446448
rect 67786 446392 70226 446448
rect 67725 446390 70226 446392
rect 67725 446387 67791 446390
rect 67633 445906 67699 445909
rect 70166 445906 70226 446148
rect 67633 445904 70226 445906
rect 67633 445848 67638 445904
rect 67694 445848 70226 445904
rect 67633 445846 70226 445848
rect 67633 445843 67699 445846
rect 61929 445772 61995 445773
rect 61878 445770 61884 445772
rect 61838 445710 61884 445770
rect 61948 445768 61995 445772
rect 102225 445770 102291 445773
rect 61990 445712 61995 445768
rect 61878 445708 61884 445710
rect 61948 445708 61995 445712
rect 61929 445707 61995 445708
rect 99790 445768 102291 445770
rect 99790 445712 102230 445768
rect 102286 445712 102291 445768
rect 99790 445710 102291 445712
rect 99790 445604 99850 445710
rect 102225 445707 102291 445710
rect 102409 445226 102475 445229
rect 99790 445224 102475 445226
rect 99790 445168 102414 445224
rect 102470 445168 102475 445224
rect 99790 445166 102475 445168
rect 99790 444924 99850 445166
rect 102409 445163 102475 445166
rect 68185 444410 68251 444413
rect 68829 444410 68895 444413
rect 70166 444410 70226 444788
rect 583520 444668 584960 444908
rect 68185 444408 70226 444410
rect 68185 444352 68190 444408
rect 68246 444352 68834 444408
rect 68890 444352 70226 444408
rect 68185 444350 70226 444352
rect 68185 444347 68251 444350
rect 68829 444347 68895 444350
rect 68277 443866 68343 443869
rect 68921 443866 68987 443869
rect 70166 443866 70226 444108
rect 68277 443864 70226 443866
rect 68277 443808 68282 443864
rect 68338 443808 68926 443864
rect 68982 443808 70226 443864
rect 68277 443806 70226 443808
rect 99606 443866 99666 444108
rect 102225 443866 102291 443869
rect 99606 443864 102291 443866
rect 99606 443808 102230 443864
rect 102286 443808 102291 443864
rect 99606 443806 102291 443808
rect 68277 443803 68343 443806
rect 68921 443803 68987 443806
rect 102225 443803 102291 443806
rect 67633 443730 67699 443733
rect 67633 443728 70226 443730
rect 67633 443672 67638 443728
rect 67694 443672 70226 443728
rect 67633 443670 70226 443672
rect 67633 443667 67699 443670
rect 70166 443564 70226 443670
rect 99414 442988 99420 443052
rect 99484 443050 99490 443052
rect 99790 443050 99850 443428
rect 127617 443050 127683 443053
rect 99484 443048 127683 443050
rect 99484 442992 127622 443048
rect 127678 442992 127683 443048
rect 99484 442990 127683 442992
rect 99484 442988 99490 442990
rect 127617 442987 127683 442990
rect 67633 442506 67699 442509
rect 70166 442506 70226 442748
rect 67633 442504 70226 442506
rect 67633 442448 67638 442504
rect 67694 442448 70226 442504
rect 67633 442446 70226 442448
rect 99790 442506 99850 442748
rect 102225 442506 102291 442509
rect 99790 442504 102291 442506
rect 99790 442448 102230 442504
rect 102286 442448 102291 442504
rect 99790 442446 102291 442448
rect 67633 442443 67699 442446
rect 102225 442443 102291 442446
rect 46657 442370 46723 442373
rect 67633 442370 67699 442373
rect 101254 442370 101260 442372
rect 46657 442368 60750 442370
rect 46657 442312 46662 442368
rect 46718 442312 60750 442368
rect 46657 442310 60750 442312
rect 46657 442307 46723 442310
rect 60690 442234 60750 442310
rect 67633 442368 70226 442370
rect 67633 442312 67638 442368
rect 67694 442312 70226 442368
rect 67633 442310 70226 442312
rect 67633 442307 67699 442310
rect 69657 442234 69723 442237
rect 60690 442232 69723 442234
rect 60690 442176 69662 442232
rect 69718 442176 69723 442232
rect 70166 442204 70226 442310
rect 99790 442310 101260 442370
rect 99790 442204 99850 442310
rect 101254 442308 101260 442310
rect 101324 442308 101330 442372
rect 60690 442174 69723 442176
rect 69657 442171 69723 442174
rect 101254 441900 101260 441964
rect 101324 441962 101330 441964
rect 103605 441962 103671 441965
rect 101324 441960 103671 441962
rect 101324 441904 103610 441960
rect 103666 441904 103671 441960
rect 101324 441902 103671 441904
rect 101324 441900 101330 441902
rect 103605 441899 103671 441902
rect 67633 441146 67699 441149
rect 70350 441146 70410 441388
rect 67633 441144 70410 441146
rect 67633 441088 67638 441144
rect 67694 441088 70410 441144
rect 67633 441086 70410 441088
rect 99606 441146 99666 441388
rect 102225 441146 102291 441149
rect 99606 441144 102291 441146
rect 99606 441088 102230 441144
rect 102286 441088 102291 441144
rect 99606 441086 102291 441088
rect 67633 441083 67699 441086
rect 102225 441083 102291 441086
rect 67633 441010 67699 441013
rect 67633 441008 70226 441010
rect 67633 440952 67638 441008
rect 67694 440952 70226 441008
rect 67633 440950 70226 440952
rect 67633 440947 67699 440950
rect 70166 440844 70226 440950
rect 69606 440676 69612 440740
rect 69676 440738 69682 440740
rect 69749 440738 69815 440741
rect 69676 440736 69815 440738
rect 69676 440680 69754 440736
rect 69810 440680 69815 440736
rect 69676 440678 69815 440680
rect 69676 440676 69682 440678
rect 69749 440675 69815 440678
rect 69657 440058 69723 440061
rect 70158 440058 70164 440060
rect 69657 440056 70164 440058
rect 69657 440000 69662 440056
rect 69718 440000 70164 440056
rect 69657 439998 70164 440000
rect 69657 439995 69723 439998
rect 70158 439996 70164 439998
rect 70228 440058 70234 440060
rect 70393 440058 70459 440061
rect 70228 440056 70504 440058
rect 70228 440000 70398 440056
rect 70454 440000 70504 440056
rect 70228 439998 70504 440000
rect 70228 439996 70234 439998
rect 70393 439995 70459 439998
rect 99373 439786 99439 439789
rect 99606 439786 99666 440028
rect 100661 439786 100727 439789
rect 99373 439784 100727 439786
rect 99373 439728 99378 439784
rect 99434 439728 100666 439784
rect 100722 439728 100727 439784
rect 99373 439726 100727 439728
rect 99373 439723 99439 439726
rect 100661 439723 100727 439726
rect 92841 439242 92907 439245
rect 93209 439242 93275 439245
rect 98085 439242 98151 439245
rect 92841 439240 98151 439242
rect 92841 439184 92846 439240
rect 92902 439184 93214 439240
rect 93270 439184 98090 439240
rect 98146 439184 98151 439240
rect 92841 439182 98151 439184
rect 92841 439179 92907 439182
rect 93209 439179 93275 439182
rect 98085 439179 98151 439182
rect 106774 439106 106780 439108
rect 97950 439046 106780 439106
rect 96613 438970 96679 438973
rect 97717 438970 97783 438973
rect 97950 438970 98010 439046
rect 106774 439044 106780 439046
rect 106844 439044 106850 439108
rect 96613 438968 98010 438970
rect 96613 438912 96618 438968
rect 96674 438912 97722 438968
rect 97778 438912 98010 438968
rect 96613 438910 98010 438912
rect 98085 438970 98151 438973
rect 103830 438970 103836 438972
rect 98085 438968 103836 438970
rect 98085 438912 98090 438968
rect 98146 438912 103836 438968
rect 98085 438910 103836 438912
rect 96613 438907 96679 438910
rect 97717 438907 97783 438910
rect 98085 438907 98151 438910
rect 103830 438908 103836 438910
rect 103900 438908 103906 438972
rect 44030 438636 44036 438700
rect 44100 438698 44106 438700
rect 77477 438698 77543 438701
rect 44100 438696 77543 438698
rect 44100 438640 77482 438696
rect 77538 438640 77543 438696
rect 44100 438638 77543 438640
rect 44100 438636 44106 438638
rect 77477 438635 77543 438638
rect 87413 437474 87479 437477
rect 115974 437474 115980 437476
rect 87413 437472 115980 437474
rect 87413 437416 87418 437472
rect 87474 437416 115980 437472
rect 87413 437414 115980 437416
rect 87413 437411 87479 437414
rect 115974 437412 115980 437414
rect 116044 437412 116050 437476
rect 84561 437338 84627 437341
rect 105486 437338 105492 437340
rect 84561 437336 105492 437338
rect 84561 437280 84566 437336
rect 84622 437280 105492 437336
rect 84561 437278 105492 437280
rect 84561 437275 84627 437278
rect 105486 437276 105492 437278
rect 105556 437276 105562 437340
rect -960 436508 480 436748
rect 65926 436732 65932 436796
rect 65996 436794 66002 436796
rect 75269 436794 75335 436797
rect 65996 436792 75335 436794
rect 65996 436736 75274 436792
rect 75330 436736 75335 436792
rect 65996 436734 75335 436736
rect 65996 436732 66002 436734
rect 75269 436731 75335 436734
rect 87413 436522 87479 436525
rect 88241 436522 88307 436525
rect 87413 436520 88307 436522
rect 87413 436464 87418 436520
rect 87474 436464 88246 436520
rect 88302 436464 88307 436520
rect 87413 436462 88307 436464
rect 87413 436459 87479 436462
rect 88241 436459 88307 436462
rect 3417 435978 3483 435981
rect 99046 435978 99052 435980
rect 3417 435976 99052 435978
rect 3417 435920 3422 435976
rect 3478 435920 99052 435976
rect 3417 435918 99052 435920
rect 3417 435915 3483 435918
rect 99046 435916 99052 435918
rect 99116 435916 99122 435980
rect 53598 435780 53604 435844
rect 53668 435842 53674 435844
rect 76005 435842 76071 435845
rect 77109 435842 77175 435845
rect 53668 435840 77175 435842
rect 53668 435784 76010 435840
rect 76066 435784 77114 435840
rect 77170 435784 77175 435840
rect 53668 435782 77175 435784
rect 53668 435780 53674 435782
rect 76005 435779 76071 435782
rect 77109 435779 77175 435782
rect 69054 435236 69060 435300
rect 69124 435298 69130 435300
rect 77385 435298 77451 435301
rect 69124 435296 77451 435298
rect 69124 435240 77390 435296
rect 77446 435240 77451 435296
rect 69124 435238 77451 435240
rect 69124 435236 69130 435238
rect 77385 435235 77451 435238
rect 57830 434556 57836 434620
rect 57900 434618 57906 434620
rect 78673 434618 78739 434621
rect 79685 434618 79751 434621
rect 57900 434616 79751 434618
rect 57900 434560 78678 434616
rect 78734 434560 79690 434616
rect 79746 434560 79751 434616
rect 57900 434558 79751 434560
rect 57900 434556 57906 434558
rect 78673 434555 78739 434558
rect 79685 434555 79751 434558
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 92473 407826 92539 407829
rect 120022 407826 120028 407828
rect 92473 407824 120028 407826
rect 92473 407768 92478 407824
rect 92534 407768 120028 407824
rect 92473 407766 120028 407768
rect 92473 407763 92539 407766
rect 120022 407764 120028 407766
rect 120092 407764 120098 407828
rect 74625 407554 74691 407557
rect 75269 407554 75335 407557
rect 74625 407552 75335 407554
rect 74625 407496 74630 407552
rect 74686 407496 75274 407552
rect 75330 407496 75335 407552
rect 74625 407494 75335 407496
rect 74625 407491 74691 407494
rect 75269 407491 75335 407494
rect 75269 407146 75335 407149
rect 338246 407146 338252 407148
rect 75269 407144 338252 407146
rect 75269 407088 75274 407144
rect 75330 407088 338252 407144
rect 75269 407086 338252 407088
rect 75269 407083 75335 407086
rect 338246 407084 338252 407086
rect 338316 407084 338322 407148
rect 88241 405106 88307 405109
rect 122598 405106 122604 405108
rect 88241 405104 122604 405106
rect 88241 405048 88246 405104
rect 88302 405048 122604 405104
rect 88241 405046 122604 405048
rect 88241 405043 88307 405046
rect 122598 405044 122604 405046
rect 122668 405044 122674 405108
rect 47853 404970 47919 404973
rect 89713 404970 89779 404973
rect 47853 404968 89779 404970
rect 47853 404912 47858 404968
rect 47914 404912 89718 404968
rect 89774 404912 89779 404968
rect 47853 404910 89779 404912
rect 47853 404907 47919 404910
rect 89713 404907 89779 404910
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 89713 404426 89779 404429
rect 340086 404426 340092 404428
rect 89713 404424 340092 404426
rect 89713 404368 89718 404424
rect 89774 404368 340092 404424
rect 89713 404366 340092 404368
rect 89713 404363 89779 404366
rect 340086 404364 340092 404366
rect 340156 404364 340162 404428
rect 42517 403610 42583 403613
rect 85665 403610 85731 403613
rect 42517 403608 85731 403610
rect 42517 403552 42522 403608
rect 42578 403552 85670 403608
rect 85726 403552 85731 403608
rect 42517 403550 85731 403552
rect 42517 403547 42583 403550
rect 85665 403547 85731 403550
rect 85665 403066 85731 403069
rect 168966 403066 168972 403068
rect 85665 403064 168972 403066
rect 85665 403008 85670 403064
rect 85726 403008 168972 403064
rect 85665 403006 168972 403008
rect 85665 403003 85731 403006
rect 168966 403004 168972 403006
rect 169036 403004 169042 403068
rect 85113 401706 85179 401709
rect 85481 401706 85547 401709
rect 160686 401706 160692 401708
rect 85113 401704 160692 401706
rect 85113 401648 85118 401704
rect 85174 401648 85486 401704
rect 85542 401648 160692 401704
rect 85113 401646 160692 401648
rect 85113 401643 85179 401646
rect 85481 401643 85547 401646
rect 160686 401644 160692 401646
rect 160756 401644 160762 401708
rect 68686 401372 68692 401436
rect 68756 401434 68762 401436
rect 68921 401434 68987 401437
rect 68756 401432 68987 401434
rect 68756 401376 68926 401432
rect 68982 401376 68987 401432
rect 68756 401374 68987 401376
rect 68756 401372 68762 401374
rect 68921 401371 68987 401374
rect 67725 400346 67791 400349
rect 68870 400346 68876 400348
rect 67725 400344 68876 400346
rect 67725 400288 67730 400344
rect 67786 400288 68876 400344
rect 67725 400286 68876 400288
rect 67725 400283 67791 400286
rect 68870 400284 68876 400286
rect 68940 400284 68946 400348
rect 108941 399666 109007 399669
rect 117998 399666 118004 399668
rect 108941 399664 118004 399666
rect 108941 399608 108946 399664
rect 109002 399608 118004 399664
rect 108941 399606 118004 399608
rect 108941 399603 109007 399606
rect 117998 399604 118004 399606
rect 118068 399604 118074 399668
rect 93669 399530 93735 399533
rect 128670 399530 128676 399532
rect 93669 399528 128676 399530
rect 93669 399472 93674 399528
rect 93730 399472 128676 399528
rect 93669 399470 128676 399472
rect 93669 399467 93735 399470
rect 128670 399468 128676 399470
rect 128740 399468 128746 399532
rect 96613 398034 96679 398037
rect 124254 398034 124260 398036
rect 96613 398032 124260 398034
rect 96613 397976 96618 398032
rect 96674 397976 124260 398032
rect 96613 397974 124260 397976
rect 96613 397971 96679 397974
rect 124254 397972 124260 397974
rect 124324 397972 124330 398036
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 68870 396204 68876 396268
rect 68940 396266 68946 396268
rect 300117 396266 300183 396269
rect 68940 396264 300183 396266
rect 68940 396208 300122 396264
rect 300178 396208 300183 396264
rect 68940 396206 300183 396208
rect 68940 396204 68946 396206
rect 300117 396203 300183 396206
rect 286317 396130 286383 396133
rect 55170 396128 286383 396130
rect 55170 396072 286322 396128
rect 286378 396072 286383 396128
rect 55170 396070 286383 396072
rect 51717 395994 51783 395997
rect 53782 395994 53788 395996
rect 51717 395992 53788 395994
rect 51717 395936 51722 395992
rect 51778 395936 53788 395992
rect 51717 395934 53788 395936
rect 51717 395931 51783 395934
rect 53782 395932 53788 395934
rect 53852 395994 53858 395996
rect 55170 395994 55230 396070
rect 286317 396067 286383 396070
rect 53852 395934 55230 395994
rect 53852 395932 53858 395934
rect 133822 394844 133828 394908
rect 133892 394906 133898 394908
rect 134701 394906 134767 394909
rect 133892 394904 134767 394906
rect 133892 394848 134706 394904
rect 134762 394848 134767 394904
rect 133892 394846 134767 394848
rect 133892 394844 133898 394846
rect 134701 394843 134767 394846
rect 103421 392594 103487 392597
rect 114686 392594 114692 392596
rect 103421 392592 114692 392594
rect 103421 392536 103426 392592
rect 103482 392536 114692 392592
rect 103421 392534 114692 392536
rect 103421 392531 103487 392534
rect 114686 392532 114692 392534
rect 114756 392532 114762 392596
rect 583520 391628 584960 391868
rect 102133 391234 102199 391237
rect 119061 391234 119127 391237
rect 129774 391234 129780 391236
rect 102133 391232 129780 391234
rect 102133 391176 102138 391232
rect 102194 391176 119066 391232
rect 119122 391176 129780 391232
rect 102133 391174 129780 391176
rect 102133 391171 102199 391174
rect 119061 391171 119127 391174
rect 129774 391172 129780 391174
rect 129844 391172 129850 391236
rect 52269 390692 52335 390693
rect 52269 390688 52316 390692
rect 52380 390690 52386 390692
rect 52269 390632 52274 390688
rect 52269 390628 52316 390632
rect 52380 390630 52426 390690
rect 52380 390628 52386 390630
rect 68686 390628 68692 390692
rect 68756 390690 68762 390692
rect 335445 390690 335511 390693
rect 68756 390688 335511 390690
rect 68756 390632 335450 390688
rect 335506 390632 335511 390688
rect 68756 390630 335511 390632
rect 68756 390628 68762 390630
rect 52269 390627 52335 390628
rect 335445 390627 335511 390630
rect 109033 389874 109099 389877
rect 110321 389874 110387 389877
rect 115974 389874 115980 389876
rect 109033 389872 115980 389874
rect 109033 389816 109038 389872
rect 109094 389816 110326 389872
rect 110382 389816 115980 389872
rect 109033 389814 115980 389816
rect 109033 389811 109099 389814
rect 110321 389811 110387 389814
rect 115974 389812 115980 389814
rect 116044 389812 116050 389876
rect 136541 389874 136607 389877
rect 170254 389874 170260 389876
rect 136541 389872 170260 389874
rect 136541 389816 136546 389872
rect 136602 389816 170260 389872
rect 136541 389814 170260 389816
rect 136541 389811 136607 389814
rect 170254 389812 170260 389814
rect 170324 389812 170330 389876
rect 57881 389196 57947 389197
rect 57830 389194 57836 389196
rect 57790 389134 57836 389194
rect 57900 389192 57947 389196
rect 57942 389136 57947 389192
rect 57830 389132 57836 389134
rect 57900 389132 57947 389136
rect 57881 389131 57947 389132
rect 143574 388996 143580 389060
rect 143644 389058 143650 389060
rect 143901 389058 143967 389061
rect 143644 389056 143967 389058
rect 143644 389000 143906 389056
rect 143962 389000 143967 389056
rect 143644 388998 143967 389000
rect 143644 388996 143650 388998
rect 143901 388995 143967 388998
rect 108982 388860 108988 388924
rect 109052 388922 109058 388924
rect 109125 388922 109191 388925
rect 109052 388920 109191 388922
rect 109052 388864 109130 388920
rect 109186 388864 109191 388920
rect 109052 388862 109191 388864
rect 109052 388860 109058 388862
rect 109125 388859 109191 388862
rect 115749 387970 115815 387973
rect 122281 387970 122347 387973
rect 115749 387968 122347 387970
rect 115749 387912 115754 387968
rect 115810 387912 122286 387968
rect 122342 387912 122347 387968
rect 115749 387910 122347 387912
rect 115749 387907 115815 387910
rect 122281 387907 122347 387910
rect 101397 387834 101463 387837
rect 191230 387834 191236 387836
rect 101397 387832 191236 387834
rect 101397 387776 101402 387832
rect 101458 387776 191236 387832
rect 101397 387774 191236 387776
rect 101397 387771 101463 387774
rect 191230 387772 191236 387774
rect 191300 387772 191306 387836
rect 50838 387636 50844 387700
rect 50908 387698 50914 387700
rect 56501 387698 56567 387701
rect 50908 387696 56567 387698
rect 50908 387640 56506 387696
rect 56562 387640 56567 387696
rect 50908 387638 56567 387640
rect 50908 387636 50914 387638
rect 56501 387635 56567 387638
rect 118734 387636 118740 387700
rect 118804 387698 118810 387700
rect 120073 387698 120139 387701
rect 118804 387696 120139 387698
rect 118804 387640 120078 387696
rect 120134 387640 120139 387696
rect 118804 387638 120139 387640
rect 118804 387636 118810 387638
rect 120073 387635 120139 387638
rect 111793 387018 111859 387021
rect 118734 387018 118740 387020
rect 111793 387016 118740 387018
rect 111793 386960 111798 387016
rect 111854 386960 118740 387016
rect 111793 386958 118740 386960
rect 111793 386955 111859 386958
rect 118734 386956 118740 386958
rect 118804 386956 118810 387020
rect 112345 386610 112411 386613
rect 122189 386610 122255 386613
rect 112345 386608 122255 386610
rect 112345 386552 112350 386608
rect 112406 386552 122194 386608
rect 122250 386552 122255 386608
rect 112345 386550 122255 386552
rect 112345 386547 112411 386550
rect 122189 386547 122255 386550
rect 58617 386474 58683 386477
rect 328545 386474 328611 386477
rect 58617 386472 328611 386474
rect 58617 386416 58622 386472
rect 58678 386416 328550 386472
rect 328606 386416 328611 386472
rect 58617 386414 328611 386416
rect 58617 386411 58683 386414
rect 328545 386411 328611 386414
rect 58934 386276 58940 386340
rect 59004 386338 59010 386340
rect 64413 386338 64479 386341
rect 59004 386336 70226 386338
rect 59004 386280 64418 386336
rect 64474 386280 70226 386336
rect 59004 386278 70226 386280
rect 59004 386276 59010 386278
rect 64413 386275 64479 386278
rect 70166 385628 70226 386278
rect 80053 386066 80119 386069
rect 80053 386064 84210 386066
rect 80053 386008 80058 386064
rect 80114 386008 84210 386064
rect 80053 386006 84210 386008
rect 80053 386003 80119 386006
rect 84150 385658 84210 386006
rect 105537 385794 105603 385797
rect 121678 385794 121684 385796
rect 105537 385792 121684 385794
rect 105537 385736 105542 385792
rect 105598 385736 121684 385792
rect 105537 385734 121684 385736
rect 105537 385731 105603 385734
rect 121678 385732 121684 385734
rect 121748 385732 121754 385796
rect 340822 385658 340828 385660
rect 84150 385598 340828 385658
rect 340822 385596 340828 385598
rect 340892 385596 340898 385660
rect 69790 385324 69796 385388
rect 69860 385386 69866 385388
rect 77477 385386 77543 385389
rect 69860 385384 77543 385386
rect 69860 385328 77482 385384
rect 77538 385328 77543 385384
rect 69860 385326 77543 385328
rect 69860 385324 69866 385326
rect 77477 385323 77543 385326
rect 117405 384978 117471 384981
rect 118509 384978 118575 384981
rect 115828 384976 118575 384978
rect 67633 384706 67699 384709
rect 70166 384706 70226 384948
rect 115828 384920 117410 384976
rect 117466 384920 118514 384976
rect 118570 384920 118575 384976
rect 115828 384918 118575 384920
rect 117405 384915 117471 384918
rect 118509 384915 118575 384918
rect 116025 384706 116091 384709
rect 67633 384704 70226 384706
rect 67633 384648 67638 384704
rect 67694 384648 70226 384704
rect 67633 384646 70226 384648
rect 115798 384704 116091 384706
rect 115798 384648 116030 384704
rect 116086 384648 116091 384704
rect 115798 384646 116091 384648
rect 67633 384643 67699 384646
rect -960 384284 480 384524
rect 115798 384298 115858 384646
rect 116025 384643 116091 384646
rect 118049 384298 118115 384301
rect 115798 384296 118115 384298
rect 115798 384268 118054 384296
rect 115828 384240 118054 384268
rect 118110 384240 118115 384296
rect 115828 384238 118115 384240
rect 118049 384235 118115 384238
rect 118141 383618 118207 383621
rect 115828 383616 118207 383618
rect 69197 383482 69263 383485
rect 70166 383482 70226 383588
rect 115828 383560 118146 383616
rect 118202 383560 118207 383616
rect 115828 383558 118207 383560
rect 118141 383555 118207 383558
rect 69197 383480 70226 383482
rect 69197 383424 69202 383480
rect 69258 383424 70226 383480
rect 69197 383422 70226 383424
rect 69197 383419 69263 383422
rect 59077 383210 59143 383213
rect 69974 383210 69980 383212
rect 59077 383208 69980 383210
rect 59077 383152 59082 383208
rect 59138 383152 69980 383208
rect 59077 383150 69980 383152
rect 59077 383147 59143 383150
rect 69974 383148 69980 383150
rect 70044 383148 70050 383212
rect 67633 382530 67699 382533
rect 70166 382530 70226 382908
rect 67633 382528 70226 382530
rect 67633 382472 67638 382528
rect 67694 382472 70226 382528
rect 67633 382470 70226 382472
rect 67633 382467 67699 382470
rect 61694 382196 61700 382260
rect 61764 382258 61770 382260
rect 63125 382258 63191 382261
rect 118601 382258 118667 382261
rect 61764 382256 64890 382258
rect 61764 382200 63130 382256
rect 63186 382200 64890 382256
rect 115828 382256 118667 382258
rect 61764 382198 64890 382200
rect 61764 382196 61770 382198
rect 63125 382195 63191 382198
rect 64830 382122 64890 382198
rect 70166 382122 70226 382228
rect 115828 382200 118606 382256
rect 118662 382200 118667 382256
rect 115828 382198 118667 382200
rect 118601 382195 118667 382198
rect 64830 382062 70226 382122
rect 118601 381578 118667 381581
rect 115828 381576 118667 381578
rect 115828 381520 118606 381576
rect 118662 381520 118667 381576
rect 115828 381518 118667 381520
rect 118601 381515 118667 381518
rect 61469 381036 61535 381037
rect 61469 381032 61516 381036
rect 61580 381034 61586 381036
rect 61469 380976 61474 381032
rect 61469 380972 61516 380976
rect 61580 380974 61626 381034
rect 61580 380972 61586 380974
rect 61469 380971 61535 380972
rect 118601 380898 118667 380901
rect 115828 380896 118667 380898
rect 69105 380762 69171 380765
rect 69657 380762 69723 380765
rect 70166 380762 70226 380868
rect 115828 380840 118606 380896
rect 118662 380840 118667 380896
rect 115828 380838 118667 380840
rect 118601 380835 118667 380838
rect 69105 380760 70226 380762
rect 69105 380704 69110 380760
rect 69166 380704 69662 380760
rect 69718 380704 70226 380760
rect 69105 380702 70226 380704
rect 69105 380699 69171 380702
rect 69657 380699 69723 380702
rect 67725 379810 67791 379813
rect 70166 379810 70226 380188
rect 122046 380156 122052 380220
rect 122116 380218 122122 380220
rect 122465 380218 122531 380221
rect 140814 380218 140820 380220
rect 122116 380216 140820 380218
rect 122116 380160 122470 380216
rect 122526 380160 140820 380216
rect 122116 380158 140820 380160
rect 122116 380156 122122 380158
rect 122465 380155 122531 380158
rect 140814 380156 140820 380158
rect 140884 380156 140890 380220
rect 67725 379808 70226 379810
rect 67725 379752 67730 379808
rect 67786 379752 70226 379808
rect 67725 379750 70226 379752
rect 67725 379747 67791 379750
rect 66161 379676 66227 379677
rect 66110 379674 66116 379676
rect 66070 379614 66116 379674
rect 66180 379672 66227 379676
rect 66222 379616 66227 379672
rect 66110 379612 66116 379614
rect 66180 379612 66227 379616
rect 66161 379611 66227 379612
rect 67633 379674 67699 379677
rect 67633 379672 70226 379674
rect 67633 379616 67638 379672
rect 67694 379616 70226 379672
rect 67633 379614 70226 379616
rect 67633 379611 67699 379614
rect 70166 379508 70226 379614
rect 118325 379538 118391 379541
rect 115828 379536 118391 379538
rect 115828 379480 118330 379536
rect 118386 379480 118391 379536
rect 115828 379478 118391 379480
rect 118325 379475 118391 379478
rect 118601 378858 118667 378861
rect 115828 378856 118667 378858
rect 115828 378800 118606 378856
rect 118662 378800 118667 378856
rect 115828 378798 118667 378800
rect 118601 378795 118667 378798
rect 124121 378724 124187 378725
rect 124070 378722 124076 378724
rect 123994 378662 124076 378722
rect 124140 378722 124187 378724
rect 128670 378722 128676 378724
rect 124140 378720 128676 378722
rect 124182 378664 128676 378720
rect 124070 378660 124076 378662
rect 124140 378662 128676 378664
rect 124140 378660 124187 378662
rect 128670 378660 128676 378662
rect 128740 378660 128746 378724
rect 124121 378659 124187 378660
rect 115974 378586 115980 378588
rect 115798 378526 115980 378586
rect 69473 378314 69539 378317
rect 69841 378314 69907 378317
rect 69473 378312 70226 378314
rect 69473 378256 69478 378312
rect 69534 378256 69846 378312
rect 69902 378256 70226 378312
rect 69473 378254 70226 378256
rect 69473 378251 69539 378254
rect 69841 378251 69907 378254
rect 70166 378148 70226 378254
rect 115798 378178 115858 378526
rect 115974 378524 115980 378526
rect 116044 378524 116050 378588
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 118049 378178 118115 378181
rect 115798 378176 118115 378178
rect 115798 378148 118054 378176
rect 115828 378120 118054 378148
rect 118110 378120 118115 378176
rect 115828 378118 118115 378120
rect 118049 378115 118115 378118
rect 67541 377362 67607 377365
rect 70166 377362 70226 377468
rect 67541 377360 70226 377362
rect 67541 377304 67546 377360
rect 67602 377304 70226 377360
rect 67541 377302 70226 377304
rect 67541 377299 67607 377302
rect 115422 377300 115428 377364
rect 115492 377362 115498 377364
rect 115492 377302 115858 377362
rect 115492 377300 115498 377302
rect 67633 377226 67699 377229
rect 67633 377224 70226 377226
rect 67633 377168 67638 377224
rect 67694 377168 70226 377224
rect 67633 377166 70226 377168
rect 67633 377163 67699 377166
rect 70166 376788 70226 377166
rect 115798 376818 115858 377302
rect 117865 376818 117931 376821
rect 115798 376816 117931 376818
rect 115798 376788 117870 376816
rect 115828 376760 117870 376788
rect 117926 376760 117931 376816
rect 115828 376758 117931 376760
rect 117865 376755 117931 376758
rect 122046 376756 122052 376820
rect 122116 376818 122122 376820
rect 122189 376818 122255 376821
rect 244917 376818 244983 376821
rect 122116 376816 244983 376818
rect 122116 376760 122194 376816
rect 122250 376760 244922 376816
rect 244978 376760 244983 376816
rect 122116 376758 244983 376760
rect 122116 376756 122122 376758
rect 122189 376755 122255 376758
rect 244917 376755 244983 376758
rect 115473 376412 115539 376413
rect 115422 376410 115428 376412
rect 115382 376350 115428 376410
rect 115492 376408 115539 376412
rect 115534 376352 115539 376408
rect 115422 376348 115428 376350
rect 115492 376348 115539 376352
rect 115473 376347 115539 376348
rect 118509 376138 118575 376141
rect 115828 376136 118575 376138
rect 115828 376080 118514 376136
rect 118570 376080 118575 376136
rect 115828 376078 118575 376080
rect 118509 376075 118575 376078
rect 67633 375594 67699 375597
rect 67633 375592 70226 375594
rect 67633 375536 67638 375592
rect 67694 375536 70226 375592
rect 67633 375534 70226 375536
rect 67633 375531 67699 375534
rect 70166 375428 70226 375534
rect 118601 375458 118667 375461
rect 115828 375456 118667 375458
rect 115828 375400 118606 375456
rect 118662 375400 118667 375456
rect 115828 375398 118667 375400
rect 118601 375395 118667 375398
rect 154573 375458 154639 375461
rect 321502 375458 321508 375460
rect 154573 375456 321508 375458
rect 154573 375400 154578 375456
rect 154634 375400 321508 375456
rect 154573 375398 321508 375400
rect 154573 375395 154639 375398
rect 321502 375396 321508 375398
rect 321572 375396 321578 375460
rect 67633 374642 67699 374645
rect 70166 374642 70226 374748
rect 67633 374640 70226 374642
rect 67633 374584 67638 374640
rect 67694 374584 70226 374640
rect 67633 374582 70226 374584
rect 135161 374642 135227 374645
rect 188286 374642 188292 374644
rect 135161 374640 188292 374642
rect 135161 374584 135166 374640
rect 135222 374584 188292 374640
rect 135161 374582 188292 374584
rect 67633 374579 67699 374582
rect 135161 374579 135227 374582
rect 188286 374580 188292 374582
rect 188356 374580 188362 374644
rect 67633 374234 67699 374237
rect 67633 374232 70226 374234
rect 67633 374176 67638 374232
rect 67694 374176 70226 374232
rect 67633 374174 70226 374176
rect 67633 374171 67699 374174
rect 70166 374068 70226 374174
rect 118601 374098 118667 374101
rect 115828 374096 118667 374098
rect 115828 374040 118606 374096
rect 118662 374040 118667 374096
rect 115828 374038 118667 374040
rect 118601 374035 118667 374038
rect 117313 373418 117379 373421
rect 115828 373416 117379 373418
rect 115828 373360 117318 373416
rect 117374 373360 117379 373416
rect 115828 373358 117379 373360
rect 117313 373355 117379 373358
rect 67633 373010 67699 373013
rect 67633 373008 70226 373010
rect 67633 372952 67638 373008
rect 67694 372952 70226 373008
rect 67633 372950 70226 372952
rect 67633 372947 67699 372950
rect 70166 372708 70226 372950
rect 118049 372740 118115 372741
rect 117998 372738 118004 372740
rect 115828 372678 118004 372738
rect 118068 372736 118115 372740
rect 118110 372680 118115 372736
rect 117998 372676 118004 372678
rect 118068 372676 118115 372680
rect 118049 372675 118115 372676
rect 65926 371922 65932 371924
rect 64830 371862 65932 371922
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 62982 371316 62988 371380
rect 63052 371378 63058 371380
rect 64830 371378 64890 371862
rect 65926 371860 65932 371862
rect 65996 371922 66002 371924
rect 70166 371922 70226 372028
rect 65996 371862 70226 371922
rect 115473 371922 115539 371925
rect 115473 371920 115858 371922
rect 115473 371864 115478 371920
rect 115534 371864 115858 371920
rect 115473 371862 115858 371864
rect 65996 371860 66002 371862
rect 115473 371859 115539 371862
rect 67633 371786 67699 371789
rect 67633 371784 70226 371786
rect 67633 371728 67638 371784
rect 67694 371728 70226 371784
rect 67633 371726 70226 371728
rect 67633 371723 67699 371726
rect 63052 371318 64890 371378
rect 70166 371348 70226 371726
rect 115798 371378 115858 371862
rect 117865 371378 117931 371381
rect 115798 371376 117931 371378
rect 115798 371348 117870 371376
rect 115828 371320 117870 371348
rect 117926 371320 117931 371376
rect 115828 371318 117931 371320
rect 63052 371316 63058 371318
rect 117865 371315 117931 371318
rect 118601 370698 118667 370701
rect 115828 370696 118667 370698
rect 115828 370640 118606 370696
rect 118662 370640 118667 370696
rect 115828 370638 118667 370640
rect 118601 370635 118667 370638
rect 69289 370154 69355 370157
rect 69289 370152 70226 370154
rect 69289 370096 69294 370152
rect 69350 370096 70226 370152
rect 69289 370094 70226 370096
rect 69289 370091 69355 370094
rect 70166 369988 70226 370094
rect 116577 370018 116643 370021
rect 118233 370018 118299 370021
rect 115828 370016 118299 370018
rect 115828 369960 116582 370016
rect 116638 369960 118238 370016
rect 118294 369960 118299 370016
rect 115828 369958 118299 369960
rect 116577 369955 116643 369958
rect 118233 369955 118299 369958
rect 69790 369882 69796 369884
rect 66118 369822 69796 369882
rect 66118 369749 66178 369822
rect 69790 369820 69796 369822
rect 69860 369820 69866 369884
rect 282913 369882 282979 369885
rect 332910 369882 332916 369884
rect 282913 369880 332916 369882
rect 282913 369824 282918 369880
rect 282974 369824 332916 369880
rect 282913 369822 332916 369824
rect 282913 369819 282979 369822
rect 332910 369820 332916 369822
rect 332980 369820 332986 369884
rect 66118 369744 66227 369749
rect 66118 369688 66166 369744
rect 66222 369688 66227 369744
rect 66118 369686 66227 369688
rect 66161 369683 66227 369686
rect 68369 369474 68435 369477
rect 68737 369474 68803 369477
rect 68369 369472 70226 369474
rect 68369 369416 68374 369472
rect 68430 369416 68742 369472
rect 68798 369416 70226 369472
rect 68369 369414 70226 369416
rect 68369 369411 68435 369414
rect 68737 369411 68803 369414
rect 70166 369308 70226 369414
rect 118601 368658 118667 368661
rect 115828 368656 118667 368658
rect 67633 368522 67699 368525
rect 70166 368522 70226 368628
rect 115828 368600 118606 368656
rect 118662 368600 118667 368656
rect 115828 368598 118667 368600
rect 118601 368595 118667 368598
rect 67633 368520 70226 368522
rect 67633 368464 67638 368520
rect 67694 368464 70226 368520
rect 67633 368462 70226 368464
rect 67633 368459 67699 368462
rect 59169 368388 59235 368389
rect 59118 368324 59124 368388
rect 59188 368386 59235 368388
rect 59188 368384 59280 368386
rect 59230 368328 59280 368384
rect 59188 368326 59280 368328
rect 59188 368324 59235 368326
rect 59169 368323 59235 368324
rect 118601 367978 118667 367981
rect 115828 367976 118667 367978
rect 115828 367920 118606 367976
rect 118662 367920 118667 367976
rect 115828 367918 118667 367920
rect 118601 367915 118667 367918
rect 59169 367706 59235 367709
rect 115565 367706 115631 367709
rect 59169 367704 70226 367706
rect 59169 367648 59174 367704
rect 59230 367648 70226 367704
rect 59169 367646 70226 367648
rect 59169 367643 59235 367646
rect 70166 367268 70226 367646
rect 115565 367704 115674 367706
rect 115565 367648 115570 367704
rect 115626 367648 115674 367704
rect 115565 367643 115674 367648
rect 115614 367268 115674 367643
rect 60590 366964 60596 367028
rect 60660 367026 60666 367028
rect 62982 367026 62988 367028
rect 60660 366966 62988 367026
rect 60660 366964 60666 366966
rect 62982 366964 62988 366966
rect 63052 366964 63058 367028
rect 67633 367026 67699 367029
rect 67633 367024 70226 367026
rect 67633 366968 67638 367024
rect 67694 366968 70226 367024
rect 67633 366966 70226 366968
rect 67633 366963 67699 366966
rect 70166 366588 70226 366966
rect 118601 365938 118667 365941
rect 115828 365936 118667 365938
rect 62982 365740 62988 365804
rect 63052 365802 63058 365804
rect 70166 365802 70226 365908
rect 115828 365880 118606 365936
rect 118662 365880 118667 365936
rect 115828 365878 118667 365880
rect 118601 365875 118667 365878
rect 63052 365742 70226 365802
rect 63052 365740 63058 365742
rect 66069 365668 66135 365669
rect 66069 365664 66116 365668
rect 66180 365666 66186 365668
rect 66069 365608 66074 365664
rect 66069 365604 66116 365608
rect 66180 365606 66226 365666
rect 66180 365604 66186 365606
rect 66069 365603 66135 365604
rect 117405 365258 117471 365261
rect 115828 365256 117471 365258
rect 115828 365200 117410 365256
rect 117466 365200 117471 365256
rect 115828 365198 117471 365200
rect 117405 365195 117471 365198
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect 115289 364850 115355 364853
rect 115289 364848 115858 364850
rect 115289 364792 115294 364848
rect 115350 364792 115858 364848
rect 115289 364790 115858 364792
rect 115289 364787 115355 364790
rect 66110 364652 66116 364716
rect 66180 364714 66186 364716
rect 66180 364654 70226 364714
rect 66180 364652 66186 364654
rect 70166 364548 70226 364654
rect 115798 364578 115858 364790
rect 117865 364578 117931 364581
rect 115798 364576 117931 364578
rect 115798 364548 117870 364576
rect 115828 364520 117870 364548
rect 117926 364520 117931 364576
rect 115828 364518 117931 364520
rect 117865 364515 117931 364518
rect 206461 364442 206527 364445
rect 330334 364442 330340 364444
rect 206461 364440 330340 364442
rect 206461 364384 206466 364440
rect 206522 364384 330340 364440
rect 206461 364382 330340 364384
rect 206461 364379 206527 364382
rect 330334 364380 330340 364382
rect 330404 364380 330410 364444
rect 67633 363762 67699 363765
rect 70166 363762 70226 363868
rect 67633 363760 70226 363762
rect 67633 363704 67638 363760
rect 67694 363704 70226 363760
rect 67633 363702 70226 363704
rect 67633 363699 67699 363702
rect 69013 363626 69079 363629
rect 146385 363626 146451 363629
rect 184054 363626 184060 363628
rect 69013 363624 70226 363626
rect 69013 363568 69018 363624
rect 69074 363568 70226 363624
rect 69013 363566 70226 363568
rect 69013 363563 69079 363566
rect 70166 363188 70226 363566
rect 146385 363624 184060 363626
rect 146385 363568 146390 363624
rect 146446 363568 184060 363624
rect 146385 363566 184060 363568
rect 146385 363563 146451 363566
rect 184054 363564 184060 363566
rect 184124 363564 184130 363628
rect 118141 363218 118207 363221
rect 115828 363216 118207 363218
rect 115828 363160 118146 363216
rect 118202 363160 118207 363216
rect 115828 363158 118207 363160
rect 118141 363155 118207 363158
rect 293401 363218 293467 363221
rect 320214 363218 320220 363220
rect 293401 363216 320220 363218
rect 293401 363160 293406 363216
rect 293462 363160 320220 363216
rect 293401 363158 320220 363160
rect 293401 363155 293467 363158
rect 320214 363156 320220 363158
rect 320284 363156 320290 363220
rect 126329 363082 126395 363085
rect 126881 363082 126947 363085
rect 325693 363082 325759 363085
rect 126329 363080 325759 363082
rect 126329 363024 126334 363080
rect 126390 363024 126886 363080
rect 126942 363024 325698 363080
rect 325754 363024 325759 363080
rect 126329 363022 325759 363024
rect 126329 363019 126395 363022
rect 126881 363019 126947 363022
rect 325693 363019 325759 363022
rect 118601 362538 118667 362541
rect 115828 362536 118667 362538
rect 67541 361994 67607 361997
rect 70166 361994 70226 362508
rect 115828 362480 118606 362536
rect 118662 362480 118667 362536
rect 115828 362478 118667 362480
rect 118601 362475 118667 362478
rect 67541 361992 70226 361994
rect 67541 361936 67546 361992
rect 67602 361936 70226 361992
rect 67541 361934 70226 361936
rect 292481 361994 292547 361997
rect 345606 361994 345612 361996
rect 292481 361992 345612 361994
rect 292481 361936 292486 361992
rect 292542 361936 345612 361992
rect 292481 361934 345612 361936
rect 67541 361931 67607 361934
rect 292481 361931 292547 361934
rect 345606 361932 345612 361934
rect 345676 361932 345682 361996
rect 117589 361858 117655 361861
rect 118601 361858 118667 361861
rect 115828 361856 118667 361858
rect 115828 361800 117594 361856
rect 117650 361800 118606 361856
rect 118662 361800 118667 361856
rect 115828 361798 118667 361800
rect 117589 361795 117655 361798
rect 118601 361795 118667 361798
rect 199469 361858 199535 361861
rect 219341 361858 219407 361861
rect 199469 361856 219407 361858
rect 199469 361800 199474 361856
rect 199530 361800 219346 361856
rect 219402 361800 219407 361856
rect 199469 361798 219407 361800
rect 199469 361795 199535 361798
rect 219341 361795 219407 361798
rect 300117 361858 300183 361861
rect 320030 361858 320036 361860
rect 300117 361856 320036 361858
rect 300117 361800 300122 361856
rect 300178 361800 320036 361856
rect 300117 361798 320036 361800
rect 300117 361795 300183 361798
rect 320030 361796 320036 361798
rect 320100 361796 320106 361860
rect 200614 361660 200620 361724
rect 200684 361722 200690 361724
rect 248965 361722 249031 361725
rect 249701 361722 249767 361725
rect 200684 361720 249767 361722
rect 200684 361664 248970 361720
rect 249026 361664 249706 361720
rect 249762 361664 249767 361720
rect 200684 361662 249767 361664
rect 200684 361660 200690 361662
rect 248965 361659 249031 361662
rect 249701 361659 249767 361662
rect 319253 361722 319319 361725
rect 320081 361722 320147 361725
rect 319253 361720 320147 361722
rect 319253 361664 319258 361720
rect 319314 361664 320086 361720
rect 320142 361664 320147 361720
rect 319253 361662 320147 361664
rect 319253 361659 319319 361662
rect 320081 361659 320147 361662
rect 118049 361178 118115 361181
rect 115828 361176 118115 361178
rect 115828 361148 118054 361176
rect 67633 360906 67699 360909
rect 70166 360906 70226 361148
rect 67633 360904 70226 360906
rect 67633 360848 67638 360904
rect 67694 360848 70226 360904
rect 67633 360846 70226 360848
rect 115798 361120 118054 361148
rect 118110 361120 118115 361176
rect 115798 361118 118115 361120
rect 67633 360843 67699 360846
rect 68001 360634 68067 360637
rect 69105 360634 69171 360637
rect 115798 360634 115858 361118
rect 118049 361115 118115 361118
rect 116025 360634 116091 360637
rect 68001 360632 70226 360634
rect 68001 360576 68006 360632
rect 68062 360576 69110 360632
rect 69166 360576 70226 360632
rect 68001 360574 70226 360576
rect 115798 360632 116091 360634
rect 115798 360576 116030 360632
rect 116086 360576 116091 360632
rect 115798 360574 116091 360576
rect 68001 360571 68067 360574
rect 69105 360571 69171 360574
rect 70166 360468 70226 360574
rect 116025 360571 116091 360574
rect 146477 360364 146543 360365
rect 146477 360360 146524 360364
rect 146588 360362 146594 360364
rect 286593 360362 286659 360365
rect 334566 360362 334572 360364
rect 146477 360304 146482 360360
rect 146477 360300 146524 360304
rect 146588 360302 146634 360362
rect 286593 360360 334572 360362
rect 286593 360304 286598 360360
rect 286654 360304 334572 360360
rect 286593 360302 334572 360304
rect 146588 360300 146594 360302
rect 146477 360299 146543 360300
rect 286593 360299 286659 360302
rect 334566 360300 334572 360302
rect 334636 360300 334642 360364
rect 199326 360164 199332 360228
rect 199396 360226 199402 360228
rect 291469 360226 291535 360229
rect 292481 360226 292547 360229
rect 199396 360224 292547 360226
rect 199396 360168 291474 360224
rect 291530 360168 292486 360224
rect 292542 360168 292547 360224
rect 199396 360166 292547 360168
rect 199396 360164 199402 360166
rect 291469 360163 291535 360166
rect 292481 360163 292547 360166
rect 304349 360226 304415 360229
rect 414657 360226 414723 360229
rect 304349 360224 414723 360226
rect 304349 360168 304354 360224
rect 304410 360168 414662 360224
rect 414718 360168 414723 360224
rect 304349 360166 414723 360168
rect 304349 360163 304415 360166
rect 414657 360163 414723 360166
rect 118601 359818 118667 359821
rect 115828 359816 118667 359818
rect 67633 359546 67699 359549
rect 70166 359546 70226 359788
rect 115828 359760 118606 359816
rect 118662 359760 118667 359816
rect 115828 359758 118667 359760
rect 118601 359755 118667 359758
rect 316861 359682 316927 359685
rect 319345 359682 319411 359685
rect 316861 359680 319411 359682
rect 316861 359624 316866 359680
rect 316922 359624 319350 359680
rect 319406 359624 319411 359680
rect 316861 359622 319411 359624
rect 316861 359619 316927 359622
rect 319345 359619 319411 359622
rect 271965 359546 272031 359549
rect 67633 359544 70226 359546
rect 67633 359488 67638 359544
rect 67694 359488 70226 359544
rect 67633 359486 70226 359488
rect 258030 359544 272031 359546
rect 258030 359488 271970 359544
rect 272026 359488 272031 359544
rect 258030 359486 272031 359488
rect 67633 359483 67699 359486
rect 149697 359410 149763 359413
rect 173014 359410 173020 359412
rect 149697 359408 173020 359410
rect 149697 359352 149702 359408
rect 149758 359352 173020 359408
rect 149697 359350 173020 359352
rect 149697 359347 149763 359350
rect 173014 359348 173020 359350
rect 173084 359348 173090 359412
rect 122189 359274 122255 359277
rect 258030 359274 258090 359486
rect 271965 359483 272031 359486
rect 314837 359546 314903 359549
rect 499573 359546 499639 359549
rect 314837 359544 499639 359546
rect 314837 359488 314842 359544
rect 314898 359488 499578 359544
rect 499634 359488 499639 359544
rect 314837 359486 499639 359488
rect 314837 359483 314903 359486
rect 499573 359483 499639 359486
rect 319345 359410 319411 359413
rect 410517 359410 410583 359413
rect 319345 359408 410583 359410
rect 319345 359352 319350 359408
rect 319406 359352 410522 359408
rect 410578 359352 410583 359408
rect 319345 359350 410583 359352
rect 319345 359347 319411 359350
rect 410517 359347 410583 359350
rect 122189 359272 258090 359274
rect 122189 359216 122194 359272
rect 122250 359216 258090 359272
rect 122189 359214 258090 359216
rect 122189 359211 122255 359214
rect 118509 359138 118575 359141
rect 115828 359136 118575 359138
rect 115828 359080 118514 359136
rect 118570 359080 118575 359136
rect 115828 359078 118575 359080
rect 118509 359075 118575 359078
rect 321737 359002 321803 359005
rect 322197 359002 322263 359005
rect 319884 359000 322263 359002
rect 319884 358944 321742 359000
rect 321798 358944 322202 359000
rect 322258 358944 322263 359000
rect 319884 358942 322263 358944
rect 321737 358939 321803 358942
rect 322197 358939 322263 358942
rect 67633 358730 67699 358733
rect 67633 358728 70226 358730
rect 67633 358672 67638 358728
rect 67694 358672 70226 358728
rect 67633 358670 70226 358672
rect 67633 358667 67699 358670
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect 70166 358428 70226 358670
rect 120022 358668 120028 358732
rect 120092 358730 120098 358732
rect 120257 358730 120323 358733
rect 120092 358728 120323 358730
rect 120092 358672 120262 358728
rect 120318 358672 120323 358728
rect 120092 358670 120323 358672
rect 120092 358668 120098 358670
rect 120257 358667 120323 358670
rect 118601 358458 118667 358461
rect 115828 358456 118667 358458
rect -960 358398 3483 358400
rect 115828 358400 118606 358456
rect 118662 358400 118667 358456
rect 115828 358398 118667 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 118601 358395 118667 358398
rect 197854 358260 197860 358324
rect 197924 358322 197930 358324
rect 197924 358262 200100 358322
rect 197924 358260 197930 358262
rect 67633 358050 67699 358053
rect 322197 358050 322263 358053
rect 331254 358050 331260 358052
rect 67633 358048 70226 358050
rect 67633 357992 67638 358048
rect 67694 357992 70226 358048
rect 67633 357990 70226 357992
rect 67633 357987 67699 357990
rect 70166 357748 70226 357990
rect 322197 358048 331260 358050
rect 322197 357992 322202 358048
rect 322258 357992 331260 358048
rect 322197 357990 331260 357992
rect 322197 357987 322263 357990
rect 331254 357988 331260 357990
rect 331324 357988 331330 358052
rect 118601 357098 118667 357101
rect 115828 357096 118667 357098
rect 67909 356962 67975 356965
rect 68686 356962 68692 356964
rect 67909 356960 68692 356962
rect 67909 356904 67914 356960
rect 67970 356904 68692 356960
rect 67909 356902 68692 356904
rect 67909 356899 67975 356902
rect 68686 356900 68692 356902
rect 68756 356962 68762 356964
rect 70166 356962 70226 357068
rect 115828 357040 118606 357096
rect 118662 357040 118667 357096
rect 115828 357038 118667 357040
rect 118601 357035 118667 357038
rect 320265 356962 320331 356965
rect 68756 356902 70226 356962
rect 319884 356960 320331 356962
rect 319884 356904 320270 356960
rect 320326 356904 320331 356960
rect 319884 356902 320331 356904
rect 68756 356900 68762 356902
rect 320265 356899 320331 356902
rect 146201 356690 146267 356693
rect 195094 356690 195100 356692
rect 146201 356688 195100 356690
rect 146201 356632 146206 356688
rect 146262 356632 195100 356688
rect 146201 356630 195100 356632
rect 146201 356627 146267 356630
rect 195094 356628 195100 356630
rect 195164 356628 195170 356692
rect 319345 356690 319411 356693
rect 494053 356690 494119 356693
rect 319345 356688 494119 356690
rect 319345 356632 319350 356688
rect 319406 356632 494058 356688
rect 494114 356632 494119 356688
rect 319345 356630 494119 356632
rect 319345 356627 319411 356630
rect 494053 356627 494119 356630
rect 118601 356418 118667 356421
rect 115828 356416 118667 356418
rect 115828 356360 118606 356416
rect 118662 356360 118667 356416
rect 115828 356358 118667 356360
rect 118601 356355 118667 356358
rect 197353 356282 197419 356285
rect 198641 356282 198707 356285
rect 197353 356280 200100 356282
rect 197353 356224 197358 356280
rect 197414 356224 198646 356280
rect 198702 356224 200100 356280
rect 197353 356222 200100 356224
rect 197353 356219 197419 356222
rect 198641 356219 198707 356222
rect 116117 355738 116183 355741
rect 118141 355738 118207 355741
rect 115828 355736 118207 355738
rect 67725 355602 67791 355605
rect 70166 355602 70226 355708
rect 115828 355680 116122 355736
rect 116178 355680 118146 355736
rect 118202 355680 118207 355736
rect 115828 355678 118207 355680
rect 116117 355675 116183 355678
rect 118141 355675 118207 355678
rect 67725 355600 70226 355602
rect 67725 355544 67730 355600
rect 67786 355544 70226 355600
rect 67725 355542 70226 355544
rect 67725 355539 67791 355542
rect 53782 355404 53788 355468
rect 53852 355466 53858 355468
rect 54201 355466 54267 355469
rect 53852 355464 54267 355466
rect 53852 355408 54206 355464
rect 54262 355408 54267 355464
rect 53852 355406 54267 355408
rect 53852 355404 53858 355406
rect 54201 355403 54267 355406
rect 320030 355268 320036 355332
rect 320100 355330 320106 355332
rect 458173 355330 458239 355333
rect 320100 355328 458239 355330
rect 320100 355272 458178 355328
rect 458234 355272 458239 355328
rect 320100 355270 458239 355272
rect 320100 355268 320106 355270
rect 458173 355267 458239 355270
rect 67633 355194 67699 355197
rect 67633 355192 70226 355194
rect 67633 355136 67638 355192
rect 67694 355136 70226 355192
rect 67633 355134 70226 355136
rect 67633 355131 67699 355134
rect 70166 355028 70226 355134
rect 117773 354378 117839 354381
rect 323117 354378 323183 354381
rect 115828 354376 117839 354378
rect 70166 353426 70226 354348
rect 115828 354320 117778 354376
rect 117834 354320 117839 354376
rect 115828 354318 117839 354320
rect 319884 354376 325710 354378
rect 319884 354320 323122 354376
rect 323178 354320 325710 354376
rect 319884 354318 325710 354320
rect 117773 354315 117839 354318
rect 323117 354315 323183 354318
rect 325650 354242 325710 354318
rect 327022 354242 327028 354244
rect 325650 354182 327028 354242
rect 327022 354180 327028 354182
rect 327092 354180 327098 354244
rect 115933 353970 115999 353973
rect 115798 353968 115999 353970
rect 115798 353912 115938 353968
rect 115994 353912 115999 353968
rect 115798 353910 115999 353912
rect 115798 353668 115858 353910
rect 115933 353907 115999 353910
rect 137134 353908 137140 353972
rect 137204 353970 137210 353972
rect 137277 353970 137343 353973
rect 199326 353970 199332 353972
rect 137204 353968 199332 353970
rect 137204 353912 137282 353968
rect 137338 353912 199332 353968
rect 137204 353910 199332 353912
rect 137204 353908 137210 353910
rect 137277 353907 137343 353910
rect 199326 353908 199332 353910
rect 199396 353908 199402 353972
rect 197997 353698 198063 353701
rect 197997 353696 200100 353698
rect 197997 353640 198002 353696
rect 198058 353640 200100 353696
rect 197997 353638 200100 353640
rect 197997 353635 198063 353638
rect 67590 353366 70226 353426
rect 58617 353290 58683 353293
rect 66662 353290 66668 353292
rect 58617 353288 66668 353290
rect 58617 353232 58622 353288
rect 58678 353232 66668 353288
rect 58617 353230 66668 353232
rect 58617 353227 58683 353230
rect 66662 353228 66668 353230
rect 66732 353290 66738 353292
rect 67590 353290 67650 353366
rect 66732 353230 67650 353290
rect 66732 353228 66738 353230
rect 68553 353154 68619 353157
rect 68553 353152 70226 353154
rect 68553 353096 68558 353152
rect 68614 353096 70226 353152
rect 68553 353094 70226 353096
rect 68553 353091 68619 353094
rect 70166 352988 70226 353094
rect 118601 353018 118667 353021
rect 115828 353016 118667 353018
rect 115828 352960 118606 353016
rect 118662 352960 118667 353016
rect 115828 352958 118667 352960
rect 118601 352955 118667 352958
rect 67633 352202 67699 352205
rect 70166 352202 70226 352308
rect 321502 352202 321508 352204
rect 67633 352200 70226 352202
rect 67633 352144 67638 352200
rect 67694 352144 70226 352200
rect 67633 352142 70226 352144
rect 319884 352142 321508 352202
rect 67633 352139 67699 352142
rect 321502 352140 321508 352142
rect 321572 352202 321578 352204
rect 322105 352202 322171 352205
rect 321572 352200 322171 352202
rect 321572 352144 322110 352200
rect 322166 352144 322171 352200
rect 321572 352142 322171 352144
rect 321572 352140 321578 352142
rect 322105 352139 322171 352142
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 117497 351658 117563 351661
rect 118601 351658 118667 351661
rect 115828 351656 118667 351658
rect 67633 351114 67699 351117
rect 70166 351114 70226 351628
rect 115828 351600 117502 351656
rect 117558 351600 118606 351656
rect 118662 351600 118667 351656
rect 115828 351598 118667 351600
rect 117497 351595 117563 351598
rect 118601 351595 118667 351598
rect 198181 351522 198247 351525
rect 198181 351520 200100 351522
rect 198181 351464 198186 351520
rect 198242 351464 200100 351520
rect 198181 351462 200100 351464
rect 198181 351459 198247 351462
rect 67633 351112 70226 351114
rect 67633 351056 67638 351112
rect 67694 351056 70226 351112
rect 67633 351054 70226 351056
rect 147765 351114 147831 351117
rect 191046 351114 191052 351116
rect 147765 351112 191052 351114
rect 147765 351056 147770 351112
rect 147826 351056 191052 351112
rect 147765 351054 191052 351056
rect 67633 351051 67699 351054
rect 147765 351051 147831 351054
rect 191046 351052 191052 351054
rect 191116 351052 191122 351116
rect 118049 350978 118115 350981
rect 115828 350976 118115 350978
rect 115828 350920 118054 350976
rect 118110 350920 118115 350976
rect 115828 350918 118115 350920
rect 118049 350915 118115 350918
rect 118601 350298 118667 350301
rect 115828 350296 118667 350298
rect 68001 350162 68067 350165
rect 68870 350162 68876 350164
rect 68001 350160 68876 350162
rect 68001 350104 68006 350160
rect 68062 350104 68876 350160
rect 68001 350102 68876 350104
rect 68001 350099 68067 350102
rect 68870 350100 68876 350102
rect 68940 350162 68946 350164
rect 70166 350162 70226 350268
rect 115828 350240 118606 350296
rect 118662 350240 118667 350296
rect 115828 350238 118667 350240
rect 118601 350235 118667 350238
rect 322749 350162 322815 350165
rect 68940 350102 70226 350162
rect 319884 350160 322815 350162
rect 319884 350104 322754 350160
rect 322810 350104 322815 350160
rect 319884 350102 322815 350104
rect 68940 350100 68946 350102
rect 322749 350099 322815 350102
rect 64413 349892 64479 349893
rect 64413 349888 64460 349892
rect 64524 349890 64530 349892
rect 64413 349832 64418 349888
rect 64413 349828 64460 349832
rect 64524 349830 64570 349890
rect 64524 349828 64530 349830
rect 64413 349827 64479 349828
rect 64597 349756 64663 349757
rect 64597 349754 64644 349756
rect 64516 349752 64644 349754
rect 64708 349754 64714 349756
rect 64516 349696 64602 349752
rect 64516 349694 64644 349696
rect 64597 349692 64644 349694
rect 64708 349694 70226 349754
rect 64708 349692 64714 349694
rect 64597 349691 64663 349692
rect 70166 349588 70226 349694
rect 198089 349618 198155 349621
rect 198089 349616 200100 349618
rect 198089 349560 198094 349616
rect 198150 349560 200100 349616
rect 198089 349558 200100 349560
rect 198089 349555 198155 349558
rect 67633 349074 67699 349077
rect 67633 349072 70226 349074
rect 67633 349016 67638 349072
rect 67694 349016 70226 349072
rect 67633 349014 70226 349016
rect 67633 349011 67699 349014
rect 70166 348908 70226 349014
rect 118601 348938 118667 348941
rect 115828 348936 118667 348938
rect 115828 348880 118606 348936
rect 118662 348880 118667 348936
rect 115828 348878 118667 348880
rect 118601 348875 118667 348878
rect 153009 348394 153075 348397
rect 186814 348394 186820 348396
rect 153009 348392 186820 348394
rect 153009 348336 153014 348392
rect 153070 348336 186820 348392
rect 153009 348334 186820 348336
rect 153009 348331 153075 348334
rect 186814 348332 186820 348334
rect 186884 348332 186890 348396
rect 117681 348258 117747 348261
rect 115828 348256 117747 348258
rect 115828 348200 117686 348256
rect 117742 348200 117747 348256
rect 115828 348198 117747 348200
rect 117681 348195 117747 348198
rect 117405 347578 117471 347581
rect 321645 347578 321711 347581
rect 115828 347576 117471 347578
rect 70166 347170 70226 347548
rect 115828 347520 117410 347576
rect 117466 347520 117471 347576
rect 115828 347518 117471 347520
rect 319884 347576 321711 347578
rect 319884 347520 321650 347576
rect 321706 347520 321711 347576
rect 319884 347518 321711 347520
rect 117405 347515 117471 347518
rect 321645 347515 321711 347518
rect 197353 347442 197419 347445
rect 197353 347440 200100 347442
rect 197353 347384 197358 347440
rect 197414 347384 200100 347440
rect 197353 347382 200100 347384
rect 197353 347379 197419 347382
rect 64830 347110 70226 347170
rect 61878 346564 61884 346628
rect 61948 346626 61954 346628
rect 64830 346626 64890 347110
rect 67633 347034 67699 347037
rect 67633 347032 70226 347034
rect 67633 346976 67638 347032
rect 67694 346976 70226 347032
rect 67633 346974 70226 346976
rect 67633 346971 67699 346974
rect 70166 346868 70226 346974
rect 61948 346566 64890 346626
rect 61948 346564 61954 346566
rect 68829 346354 68895 346357
rect 144269 346354 144335 346357
rect 200614 346354 200620 346356
rect 68829 346352 70226 346354
rect 68829 346296 68834 346352
rect 68890 346296 70226 346352
rect 68829 346294 70226 346296
rect 68829 346291 68895 346294
rect 70166 346188 70226 346294
rect 144269 346352 200620 346354
rect 144269 346296 144274 346352
rect 144330 346296 200620 346352
rect 144269 346294 200620 346296
rect 144269 346291 144335 346294
rect 200614 346292 200620 346294
rect 200684 346292 200690 346356
rect 118509 346218 118575 346221
rect 115828 346216 118575 346218
rect 115828 346160 118514 346216
rect 118570 346160 118575 346216
rect 115828 346158 118575 346160
rect 118509 346155 118575 346158
rect 143441 345674 143507 345677
rect 189942 345674 189948 345676
rect 143441 345672 189948 345674
rect 143441 345616 143446 345672
rect 143502 345616 189948 345672
rect 143441 345614 189948 345616
rect 143441 345611 143507 345614
rect 189942 345612 189948 345614
rect 190012 345612 190018 345676
rect 118601 345538 118667 345541
rect 322473 345538 322539 345541
rect 115828 345536 118667 345538
rect -960 345402 480 345492
rect 115828 345480 118606 345536
rect 118662 345480 118667 345536
rect 115828 345478 118667 345480
rect 319884 345536 322539 345538
rect 319884 345480 322478 345536
rect 322534 345480 322539 345536
rect 319884 345478 322539 345480
rect 118601 345475 118667 345478
rect 322473 345475 322539 345478
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 68645 344994 68711 344997
rect 68645 344992 70226 344994
rect 68645 344936 68650 344992
rect 68706 344936 70226 344992
rect 68645 344934 70226 344936
rect 68645 344931 68711 344934
rect 70166 344828 70226 344934
rect 118601 344858 118667 344861
rect 115828 344856 118667 344858
rect 115828 344800 118606 344856
rect 118662 344800 118667 344856
rect 115828 344798 118667 344800
rect 118601 344795 118667 344798
rect 198089 344722 198155 344725
rect 198089 344720 200100 344722
rect 198089 344664 198094 344720
rect 198150 344664 200100 344720
rect 198089 344662 200100 344664
rect 198089 344659 198155 344662
rect 67633 343770 67699 343773
rect 70166 343770 70226 344148
rect 67633 343768 70226 343770
rect 67633 343712 67638 343768
rect 67694 343712 70226 343768
rect 67633 343710 70226 343712
rect 67633 343707 67699 343710
rect 67633 343634 67699 343637
rect 126789 343636 126855 343637
rect 67633 343632 70226 343634
rect 67633 343576 67638 343632
rect 67694 343576 70226 343632
rect 67633 343574 70226 343576
rect 67633 343571 67699 343574
rect 70166 343468 70226 343574
rect 126789 343632 126836 343636
rect 126900 343634 126906 343636
rect 126789 343576 126794 343632
rect 126789 343572 126836 343576
rect 126900 343574 126946 343634
rect 126900 343572 126906 343574
rect 126789 343571 126855 343572
rect 117497 343498 117563 343501
rect 115828 343496 117563 343498
rect 115828 343440 117502 343496
rect 117558 343440 117563 343496
rect 115828 343438 117563 343440
rect 117497 343435 117563 343438
rect 322473 343362 322539 343365
rect 319884 343360 322539 343362
rect 319884 343304 322478 343360
rect 322534 343304 322539 343360
rect 319884 343302 322539 343304
rect 322473 343299 322539 343302
rect 126789 342954 126855 342957
rect 133086 342954 133092 342956
rect 126789 342952 133092 342954
rect 126789 342896 126794 342952
rect 126850 342896 133092 342952
rect 126789 342894 133092 342896
rect 126789 342891 126855 342894
rect 133086 342892 133092 342894
rect 133156 342892 133162 342956
rect 150525 342954 150591 342957
rect 193806 342954 193812 342956
rect 150525 342952 193812 342954
rect 150525 342896 150530 342952
rect 150586 342896 193812 342952
rect 150525 342894 193812 342896
rect 150525 342891 150591 342894
rect 193806 342892 193812 342894
rect 193876 342892 193882 342956
rect 117865 342818 117931 342821
rect 115828 342816 117931 342818
rect 115828 342760 117870 342816
rect 117926 342760 117931 342816
rect 115828 342758 117931 342760
rect 117865 342755 117931 342758
rect 197997 342682 198063 342685
rect 197997 342680 200100 342682
rect 197997 342624 198002 342680
rect 198058 342624 200100 342680
rect 197997 342622 200100 342624
rect 197997 342619 198063 342622
rect 118601 342138 118667 342141
rect 120022 342138 120028 342140
rect 115828 342136 120028 342138
rect 68645 342002 68711 342005
rect 70534 342002 70594 342108
rect 115828 342080 118606 342136
rect 118662 342080 120028 342136
rect 115828 342078 120028 342080
rect 118601 342075 118667 342078
rect 120022 342076 120028 342078
rect 120092 342076 120098 342140
rect 68645 342000 70594 342002
rect 68645 341944 68650 342000
rect 68706 341944 70594 342000
rect 68645 341942 70594 341944
rect 68645 341939 68711 341942
rect 70534 341732 70594 341942
rect 70526 341668 70532 341732
rect 70596 341668 70602 341732
rect 322565 341458 322631 341461
rect 319884 341456 322631 341458
rect 67633 341050 67699 341053
rect 70166 341050 70226 341428
rect 319884 341400 322570 341456
rect 322626 341400 322631 341456
rect 319884 341398 322631 341400
rect 322565 341395 322631 341398
rect 67633 341048 70226 341050
rect 67633 340992 67638 341048
rect 67694 340992 70226 341048
rect 67633 340990 70226 340992
rect 67633 340987 67699 340990
rect 117313 340778 117379 340781
rect 115828 340776 117379 340778
rect 67633 340234 67699 340237
rect 70166 340234 70226 340748
rect 115828 340720 117318 340776
rect 117374 340720 117379 340776
rect 115828 340718 117379 340720
rect 117313 340715 117379 340718
rect 197353 340642 197419 340645
rect 197353 340640 200100 340642
rect 197353 340584 197358 340640
rect 197414 340584 200100 340640
rect 197353 340582 200100 340584
rect 197353 340579 197419 340582
rect 67633 340232 70226 340234
rect 67633 340176 67638 340232
rect 67694 340176 70226 340232
rect 67633 340174 70226 340176
rect 67633 340171 67699 340174
rect 69606 340036 69612 340100
rect 69676 340098 69682 340100
rect 69749 340098 69815 340101
rect 117405 340098 117471 340101
rect 69676 340096 69815 340098
rect 69676 340040 69754 340096
rect 69810 340040 69815 340096
rect 115828 340096 117471 340098
rect 115828 340068 117410 340096
rect 69676 340038 69815 340040
rect 69676 340036 69682 340038
rect 69749 340035 69815 340038
rect 115798 340040 117410 340068
rect 117466 340040 117471 340096
rect 115798 340038 117471 340040
rect 115105 339554 115171 339557
rect 115798 339554 115858 340038
rect 117405 340035 117471 340038
rect 115105 339552 115858 339554
rect 115105 339496 115110 339552
rect 115166 339496 115858 339552
rect 115105 339494 115858 339496
rect 115105 339491 115171 339494
rect 40953 339418 41019 339421
rect 75821 339418 75887 339421
rect 124254 339418 124260 339420
rect 40953 339416 75887 339418
rect 40953 339360 40958 339416
rect 41014 339360 75826 339416
rect 75882 339360 75887 339416
rect 40953 339358 75887 339360
rect 40953 339355 41019 339358
rect 75821 339355 75887 339358
rect 103470 339358 124260 339418
rect 102225 339282 102291 339285
rect 103470 339282 103530 339358
rect 124254 339356 124260 339358
rect 124324 339356 124330 339420
rect 102225 339280 103530 339282
rect 102225 339224 102230 339280
rect 102286 339224 103530 339280
rect 102225 339222 103530 339224
rect 102225 339219 102291 339222
rect 66662 338676 66668 338740
rect 66732 338738 66738 338740
rect 77293 338738 77359 338741
rect 322381 338738 322447 338741
rect 66732 338736 77359 338738
rect 66732 338680 77298 338736
rect 77354 338680 77359 338736
rect 66732 338678 77359 338680
rect 319884 338736 322447 338738
rect 319884 338680 322386 338736
rect 322442 338680 322447 338736
rect 319884 338678 322447 338680
rect 66732 338676 66738 338678
rect 77293 338675 77359 338678
rect 322381 338675 322447 338678
rect 583520 338452 584960 338692
rect 99281 338194 99347 338197
rect 102225 338194 102291 338197
rect 99281 338192 102291 338194
rect 99281 338136 99286 338192
rect 99342 338136 102230 338192
rect 102286 338136 102291 338192
rect 99281 338134 102291 338136
rect 99281 338131 99347 338134
rect 102225 338131 102291 338134
rect 142245 338060 142311 338061
rect 122598 338058 122604 338060
rect 93810 337998 122604 338058
rect 66161 337922 66227 337925
rect 79317 337922 79383 337925
rect 66161 337920 79383 337922
rect 66161 337864 66166 337920
rect 66222 337864 79322 337920
rect 79378 337864 79383 337920
rect 66161 337862 79383 337864
rect 66161 337859 66227 337862
rect 79317 337859 79383 337862
rect 89989 337786 90055 337789
rect 90909 337786 90975 337789
rect 93810 337786 93870 337998
rect 122598 337996 122604 337998
rect 122668 337996 122674 338060
rect 142245 338056 142292 338060
rect 142356 338058 142362 338060
rect 142245 338000 142250 338056
rect 142245 337996 142292 338000
rect 142356 337998 142402 338058
rect 142356 337996 142362 337998
rect 142245 337995 142311 337996
rect 111241 337922 111307 337925
rect 111609 337922 111675 337925
rect 121678 337922 121684 337924
rect 111241 337920 121684 337922
rect 111241 337864 111246 337920
rect 111302 337864 111614 337920
rect 111670 337864 121684 337920
rect 111241 337862 121684 337864
rect 111241 337859 111307 337862
rect 111609 337859 111675 337862
rect 121678 337860 121684 337862
rect 121748 337860 121754 337924
rect 197353 337922 197419 337925
rect 197353 337920 200100 337922
rect 197353 337864 197358 337920
rect 197414 337864 200100 337920
rect 197353 337862 200100 337864
rect 197353 337859 197419 337862
rect 89989 337784 93870 337786
rect 89989 337728 89994 337784
rect 90050 337728 90914 337784
rect 90970 337728 93870 337784
rect 89989 337726 93870 337728
rect 89989 337723 90055 337726
rect 90909 337723 90975 337726
rect 322473 336562 322539 336565
rect 319884 336560 322539 336562
rect 319884 336504 322478 336560
rect 322534 336504 322539 336560
rect 319884 336502 322539 336504
rect 322473 336499 322539 336502
rect 58985 336018 59051 336021
rect 77385 336018 77451 336021
rect 177389 336018 177455 336021
rect 58985 336016 177455 336018
rect 58985 335960 58990 336016
rect 59046 335960 77390 336016
rect 77446 335960 177394 336016
rect 177450 335960 177455 336016
rect 58985 335958 177455 335960
rect 58985 335955 59051 335958
rect 77385 335955 77451 335958
rect 177389 335955 177455 335958
rect 197721 335882 197787 335885
rect 197721 335880 200100 335882
rect 197721 335824 197726 335880
rect 197782 335824 200100 335880
rect 197721 335822 200100 335824
rect 197721 335819 197787 335822
rect 322473 334658 322539 334661
rect 319884 334656 322539 334658
rect 319884 334600 322478 334656
rect 322534 334600 322539 334656
rect 319884 334598 322539 334600
rect 322473 334595 322539 334598
rect 198917 333842 198983 333845
rect 198917 333840 200100 333842
rect 198917 333784 198922 333840
rect 198978 333784 200100 333840
rect 198917 333782 200100 333784
rect 198917 333779 198983 333782
rect 172421 333298 172487 333301
rect 197854 333298 197860 333300
rect 172421 333296 197860 333298
rect 172421 333240 172426 333296
rect 172482 333240 197860 333296
rect 172421 333238 197860 333240
rect 172421 333235 172487 333238
rect 197854 333236 197860 333238
rect 197924 333236 197930 333300
rect 70894 332556 70900 332620
rect 70964 332618 70970 332620
rect 172421 332618 172487 332621
rect 70964 332616 172487 332618
rect 70964 332560 172426 332616
rect 172482 332560 172487 332616
rect 70964 332558 172487 332560
rect 70964 332556 70970 332558
rect 172421 332555 172487 332558
rect -960 332196 480 332436
rect 107653 331802 107719 331805
rect 122046 331802 122052 331804
rect 107653 331800 122052 331802
rect 107653 331744 107658 331800
rect 107714 331744 122052 331800
rect 107653 331742 122052 331744
rect 107653 331739 107719 331742
rect 122046 331740 122052 331742
rect 122116 331740 122122 331804
rect 124806 331740 124812 331804
rect 124876 331802 124882 331804
rect 125501 331802 125567 331805
rect 133822 331802 133828 331804
rect 124876 331800 133828 331802
rect 124876 331744 125506 331800
rect 125562 331744 133828 331800
rect 124876 331742 133828 331744
rect 124876 331740 124882 331742
rect 125501 331739 125567 331742
rect 133822 331740 133828 331742
rect 133892 331740 133898 331804
rect 197353 331802 197419 331805
rect 321553 331802 321619 331805
rect 322197 331802 322263 331805
rect 197353 331800 200100 331802
rect 197353 331744 197358 331800
rect 197414 331744 200100 331800
rect 197353 331742 200100 331744
rect 319884 331800 322263 331802
rect 319884 331744 321558 331800
rect 321614 331744 322202 331800
rect 322258 331744 322263 331800
rect 319884 331742 322263 331744
rect 197353 331739 197419 331742
rect 321553 331739 321619 331742
rect 322197 331739 322263 331742
rect 96521 331122 96587 331125
rect 128854 331122 128860 331124
rect 96521 331120 128860 331122
rect 96521 331064 96526 331120
rect 96582 331064 128860 331120
rect 96521 331062 128860 331064
rect 96521 331059 96587 331062
rect 128854 331060 128860 331062
rect 128924 331060 128930 331124
rect 324313 331122 324379 331125
rect 324589 331122 324655 331125
rect 326654 331122 326660 331124
rect 324313 331120 326660 331122
rect 324313 331064 324318 331120
rect 324374 331064 324594 331120
rect 324650 331064 326660 331120
rect 324313 331062 326660 331064
rect 324313 331059 324379 331062
rect 324589 331059 324655 331062
rect 326654 331060 326660 331062
rect 326724 331060 326730 331124
rect 95785 330714 95851 330717
rect 96521 330714 96587 330717
rect 95785 330712 96587 330714
rect 95785 330656 95790 330712
rect 95846 330656 96526 330712
rect 96582 330656 96587 330712
rect 95785 330654 96587 330656
rect 95785 330651 95851 330654
rect 96521 330651 96587 330654
rect 322749 329898 322815 329901
rect 319884 329896 322815 329898
rect 319884 329840 322754 329896
rect 322810 329840 322815 329896
rect 319884 329838 322815 329840
rect 322749 329835 322815 329838
rect 197353 329082 197419 329085
rect 197353 329080 200100 329082
rect 197353 329024 197358 329080
rect 197414 329024 200100 329080
rect 197353 329022 200100 329024
rect 197353 329019 197419 329022
rect 322749 327722 322815 327725
rect 319884 327720 322815 327722
rect 319884 327664 322754 327720
rect 322810 327664 322815 327720
rect 319884 327662 322815 327664
rect 322749 327659 322815 327662
rect 197353 327178 197419 327181
rect 197353 327176 200100 327178
rect 197353 327120 197358 327176
rect 197414 327120 200100 327176
rect 197353 327118 200100 327120
rect 197353 327115 197419 327118
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 69054 324940 69060 325004
rect 69124 325002 69130 325004
rect 198273 325002 198339 325005
rect 320357 325002 320423 325005
rect 69124 324942 180810 325002
rect 69124 324940 69130 324942
rect 180750 324866 180810 324942
rect 198273 325000 200100 325002
rect 198273 324944 198278 325000
rect 198334 324944 200100 325000
rect 198273 324942 200100 324944
rect 319884 325000 320423 325002
rect 319884 324944 320362 325000
rect 320418 324944 320423 325000
rect 319884 324942 320423 324944
rect 198273 324939 198339 324942
rect 320357 324939 320423 324942
rect 198641 324866 198707 324869
rect 180750 324864 198707 324866
rect 180750 324808 198646 324864
rect 198702 324808 198707 324864
rect 180750 324806 198707 324808
rect 198641 324803 198707 324806
rect 322473 322962 322539 322965
rect 319884 322960 322539 322962
rect 319884 322904 322478 322960
rect 322534 322904 322539 322960
rect 319884 322902 322539 322904
rect 322473 322899 322539 322902
rect 197353 322418 197419 322421
rect 197353 322416 200100 322418
rect 197353 322360 197358 322416
rect 197414 322360 200100 322416
rect 197353 322358 200100 322360
rect 197353 322355 197419 322358
rect 71078 322084 71084 322148
rect 71148 322146 71154 322148
rect 140221 322146 140287 322149
rect 71148 322144 140287 322146
rect 71148 322088 140226 322144
rect 140282 322088 140287 322144
rect 71148 322086 140287 322088
rect 71148 322084 71154 322086
rect 140221 322083 140287 322086
rect 322841 320922 322907 320925
rect 319884 320920 322907 320922
rect 319884 320864 322846 320920
rect 322902 320864 322907 320920
rect 319884 320862 322907 320864
rect 322841 320859 322907 320862
rect 86401 320786 86467 320789
rect 178534 320786 178540 320788
rect 86401 320784 178540 320786
rect 86401 320728 86406 320784
rect 86462 320728 178540 320784
rect 86401 320726 178540 320728
rect 86401 320723 86467 320726
rect 178534 320724 178540 320726
rect 178604 320724 178610 320788
rect 197353 320242 197419 320245
rect 197353 320240 200100 320242
rect 197353 320184 197358 320240
rect 197414 320184 200100 320240
rect 197353 320182 200100 320184
rect 197353 320179 197419 320182
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 321502 318882 321508 318884
rect 319884 318822 321508 318882
rect 321502 318820 321508 318822
rect 321572 318820 321578 318884
rect 128629 318748 128695 318749
rect 128629 318744 128676 318748
rect 128740 318746 128746 318748
rect 128629 318688 128634 318744
rect 128629 318684 128676 318688
rect 128740 318686 128786 318746
rect 128740 318684 128746 318686
rect 128629 318683 128695 318684
rect 197353 318202 197419 318205
rect 197353 318200 200100 318202
rect 197353 318144 197358 318200
rect 197414 318144 200100 318200
rect 197353 318142 200100 318144
rect 197353 318139 197419 318142
rect 322473 316298 322539 316301
rect 319884 316296 322539 316298
rect 319884 316240 322478 316296
rect 322534 316240 322539 316296
rect 319884 316238 322539 316240
rect 322473 316235 322539 316238
rect 197353 315482 197419 315485
rect 197353 315480 200100 315482
rect 197353 315424 197358 315480
rect 197414 315424 200100 315480
rect 197353 315422 200100 315424
rect 197353 315419 197419 315422
rect 322473 314258 322539 314261
rect 319884 314256 322539 314258
rect 319884 314200 322478 314256
rect 322534 314200 322539 314256
rect 319884 314198 322539 314200
rect 322473 314195 322539 314198
rect 197353 313442 197419 313445
rect 198825 313442 198891 313445
rect 197353 313440 200100 313442
rect 197353 313384 197358 313440
rect 197414 313384 198830 313440
rect 198886 313384 200100 313440
rect 197353 313382 200100 313384
rect 197353 313379 197419 313382
rect 198825 313379 198891 313382
rect 322841 312218 322907 312221
rect 319884 312216 322907 312218
rect 319884 312160 322846 312216
rect 322902 312160 322907 312216
rect 319884 312158 322907 312160
rect 322841 312155 322907 312158
rect 580257 312082 580323 312085
rect 583520 312082 584960 312172
rect 580257 312080 584960 312082
rect 580257 312024 580262 312080
rect 580318 312024 584960 312080
rect 580257 312022 584960 312024
rect 580257 312019 580323 312022
rect 583520 311932 584960 312022
rect 197353 311402 197419 311405
rect 197353 311400 200100 311402
rect 197353 311344 197358 311400
rect 197414 311344 200100 311400
rect 197353 311342 200100 311344
rect 197353 311339 197419 311342
rect 322473 309498 322539 309501
rect 319884 309496 322539 309498
rect 319884 309440 322478 309496
rect 322534 309440 322539 309496
rect 319884 309438 322539 309440
rect 322473 309435 322539 309438
rect 197353 309362 197419 309365
rect 197353 309360 200100 309362
rect 197353 309304 197358 309360
rect 197414 309304 200100 309360
rect 197353 309302 200100 309304
rect 197353 309299 197419 309302
rect 125777 309228 125843 309229
rect 125726 309226 125732 309228
rect 125686 309166 125732 309226
rect 125796 309224 125843 309228
rect 125838 309168 125843 309224
rect 125726 309164 125732 309166
rect 125796 309164 125843 309168
rect 125777 309163 125843 309164
rect 69238 307804 69244 307868
rect 69308 307866 69314 307868
rect 165429 307866 165495 307869
rect 69308 307864 165495 307866
rect 69308 307808 165434 307864
rect 165490 307808 165495 307864
rect 69308 307806 165495 307808
rect 69308 307804 69314 307806
rect 165429 307803 165495 307806
rect 319529 307730 319595 307733
rect 321737 307730 321803 307733
rect 319302 307728 321803 307730
rect 319302 307672 319534 307728
rect 319590 307672 321742 307728
rect 321798 307672 321803 307728
rect 319302 307670 321803 307672
rect 319302 307428 319362 307670
rect 319529 307667 319595 307670
rect 321737 307667 321803 307670
rect 197261 306642 197327 306645
rect 197261 306640 200100 306642
rect 197261 306584 197266 306640
rect 197322 306584 200100 306640
rect 197261 306582 200100 306584
rect 197261 306579 197327 306582
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 322473 305282 322539 305285
rect 319884 305280 322539 305282
rect 319884 305224 322478 305280
rect 322534 305224 322539 305280
rect 319884 305222 322539 305224
rect 322473 305219 322539 305222
rect 197721 304602 197787 304605
rect 197721 304600 200100 304602
rect 197721 304544 197726 304600
rect 197782 304544 200100 304600
rect 197721 304542 200100 304544
rect 197721 304539 197787 304542
rect 322473 303242 322539 303245
rect 319884 303240 322539 303242
rect 319884 303184 322478 303240
rect 322534 303184 322539 303240
rect 319884 303182 322539 303184
rect 322473 303179 322539 303182
rect 197353 302562 197419 302565
rect 197353 302560 200100 302562
rect 197353 302504 197358 302560
rect 197414 302504 200100 302560
rect 197353 302502 200100 302504
rect 197353 302499 197419 302502
rect 71078 302228 71084 302292
rect 71148 302290 71154 302292
rect 186221 302290 186287 302293
rect 71148 302288 186287 302290
rect 71148 302232 186226 302288
rect 186282 302232 186287 302288
rect 71148 302230 186287 302232
rect 71148 302228 71154 302230
rect 186221 302227 186287 302230
rect 322565 300522 322631 300525
rect 319884 300520 322631 300522
rect 319884 300464 322570 300520
rect 322626 300464 322631 300520
rect 319884 300462 322631 300464
rect 322565 300459 322631 300462
rect 52177 300114 52243 300117
rect 125593 300114 125659 300117
rect 52177 300112 125659 300114
rect 52177 300056 52182 300112
rect 52238 300056 125598 300112
rect 125654 300056 125659 300112
rect 52177 300054 125659 300056
rect 52177 300051 52243 300054
rect 125593 300051 125659 300054
rect 197353 299978 197419 299981
rect 197353 299976 200100 299978
rect 197353 299920 197358 299976
rect 197414 299920 200100 299976
rect 197353 299918 200100 299920
rect 197353 299915 197419 299918
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 583520 298604 584960 298694
rect 319486 298213 319546 298452
rect 67541 298210 67607 298213
rect 147121 298210 147187 298213
rect 67541 298208 147187 298210
rect 67541 298152 67546 298208
rect 67602 298152 147126 298208
rect 147182 298152 147187 298208
rect 67541 298150 147187 298152
rect 319486 298208 319595 298213
rect 319486 298152 319534 298208
rect 319590 298152 319595 298208
rect 319486 298150 319595 298152
rect 67541 298147 67607 298150
rect 147121 298147 147187 298150
rect 319529 298147 319595 298150
rect 197353 297802 197419 297805
rect 197353 297800 200100 297802
rect 197353 297744 197358 297800
rect 197414 297744 200100 297800
rect 197353 297742 200100 297744
rect 197353 297739 197419 297742
rect 56501 297394 56567 297397
rect 91277 297394 91343 297397
rect 56501 297392 91343 297394
rect 56501 297336 56506 297392
rect 56562 297336 91282 297392
rect 91338 297336 91343 297392
rect 56501 297334 91343 297336
rect 56501 297331 56567 297334
rect 91277 297331 91343 297334
rect 91277 296850 91343 296853
rect 151169 296850 151235 296853
rect 91277 296848 151235 296850
rect 91277 296792 91282 296848
rect 91338 296792 151174 296848
rect 151230 296792 151235 296848
rect 91277 296790 151235 296792
rect 91277 296787 91343 296790
rect 151169 296787 151235 296790
rect 322473 296442 322539 296445
rect 319884 296440 322539 296442
rect 319884 296384 322478 296440
rect 322534 296384 322539 296440
rect 319884 296382 322539 296384
rect 322473 296379 322539 296382
rect 76557 296034 76623 296037
rect 120165 296034 120231 296037
rect 76557 296032 120231 296034
rect 76557 295976 76562 296032
rect 76618 295976 120170 296032
rect 120226 295976 120231 296032
rect 76557 295974 120231 295976
rect 76557 295971 76623 295974
rect 120165 295971 120231 295974
rect 197445 295762 197511 295765
rect 197445 295760 200100 295762
rect 197445 295704 197450 295760
rect 197506 295704 200100 295760
rect 197445 295702 200100 295704
rect 197445 295699 197511 295702
rect 107377 295354 107443 295357
rect 148593 295354 148659 295357
rect 107377 295352 148659 295354
rect 107377 295296 107382 295352
rect 107438 295296 148598 295352
rect 148654 295296 148659 295352
rect 107377 295294 148659 295296
rect 107377 295291 107443 295294
rect 148593 295291 148659 295294
rect 118969 295218 119035 295221
rect 123661 295218 123727 295221
rect 118969 295216 123727 295218
rect 118969 295160 118974 295216
rect 119030 295160 123666 295216
rect 123722 295160 123727 295216
rect 118969 295158 123727 295160
rect 118969 295155 119035 295158
rect 123661 295155 123727 295158
rect 114185 294674 114251 294677
rect 123477 294674 123543 294677
rect 114185 294672 123543 294674
rect 114185 294616 114190 294672
rect 114246 294616 123482 294672
rect 123538 294616 123543 294672
rect 114185 294614 123543 294616
rect 114185 294611 114251 294614
rect 123477 294611 123543 294614
rect 104157 294538 104223 294541
rect 195329 294538 195395 294541
rect 104157 294536 195395 294538
rect 104157 294480 104162 294536
rect 104218 294480 195334 294536
rect 195390 294480 195395 294536
rect 104157 294478 195395 294480
rect 104157 294475 104223 294478
rect 195329 294475 195395 294478
rect 196709 293722 196775 293725
rect 322841 293722 322907 293725
rect 196709 293720 200100 293722
rect 196709 293664 196714 293720
rect 196770 293664 200100 293720
rect 196709 293662 200100 293664
rect 319884 293720 322907 293722
rect 319884 293664 322846 293720
rect 322902 293664 322907 293720
rect 319884 293662 322907 293664
rect 196709 293659 196775 293662
rect 322841 293659 322907 293662
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 107469 293178 107535 293181
rect 124397 293178 124463 293181
rect 107469 293176 124463 293178
rect 107469 293120 107474 293176
rect 107530 293120 124402 293176
rect 124458 293120 124463 293176
rect 107469 293118 124463 293120
rect 107469 293115 107535 293118
rect 124397 293115 124463 293118
rect 97073 292634 97139 292637
rect 123334 292634 123340 292636
rect 97073 292632 123340 292634
rect 97073 292576 97078 292632
rect 97134 292576 123340 292632
rect 97073 292574 123340 292576
rect 97073 292571 97139 292574
rect 123334 292572 123340 292574
rect 123404 292572 123410 292636
rect 71681 292362 71747 292365
rect 70718 292360 71747 292362
rect 70718 292304 71686 292360
rect 71742 292304 71747 292360
rect 70718 292302 71747 292304
rect 70718 291788 70778 292302
rect 71681 292299 71747 292302
rect 103145 291954 103211 291957
rect 126421 291954 126487 291957
rect 103145 291952 126487 291954
rect 103145 291896 103150 291952
rect 103206 291896 126426 291952
rect 126482 291896 126487 291952
rect 103145 291894 126487 291896
rect 103145 291891 103211 291894
rect 126421 291891 126487 291894
rect 121453 291818 121519 291821
rect 119876 291816 121519 291818
rect 119876 291760 121458 291816
rect 121514 291760 121519 291816
rect 119876 291758 121519 291760
rect 121453 291755 121519 291758
rect 322473 291682 322539 291685
rect 319884 291680 322539 291682
rect 319884 291624 322478 291680
rect 322534 291624 322539 291680
rect 319884 291622 322539 291624
rect 322473 291619 322539 291622
rect 121545 291138 121611 291141
rect 119876 291136 121611 291138
rect 67633 290866 67699 290869
rect 70350 290866 70410 291108
rect 119876 291080 121550 291136
rect 121606 291080 121611 291136
rect 119876 291078 121611 291080
rect 121545 291075 121611 291078
rect 197445 291002 197511 291005
rect 197445 291000 200100 291002
rect 197445 290944 197450 291000
rect 197506 290944 200100 291000
rect 197445 290942 200100 290944
rect 197445 290939 197511 290942
rect 67633 290864 70410 290866
rect 67633 290808 67638 290864
rect 67694 290808 70410 290864
rect 67633 290806 70410 290808
rect 67633 290803 67699 290806
rect 121453 290458 121519 290461
rect 119876 290456 121519 290458
rect 67633 289914 67699 289917
rect 70166 289914 70226 290428
rect 119876 290400 121458 290456
rect 121514 290400 121519 290456
rect 119876 290398 121519 290400
rect 121453 290395 121519 290398
rect 67633 289912 70226 289914
rect 67633 289856 67638 289912
rect 67694 289856 70226 289912
rect 67633 289854 70226 289856
rect 67633 289851 67699 289854
rect 121453 289778 121519 289781
rect 119876 289776 121519 289778
rect 70534 289508 70594 289748
rect 119876 289720 121458 289776
rect 121514 289720 121519 289776
rect 119876 289718 121519 289720
rect 121453 289715 121519 289718
rect 321553 289642 321619 289645
rect 319884 289640 321619 289642
rect 319884 289584 321558 289640
rect 321614 289584 321619 289640
rect 319884 289582 321619 289584
rect 321553 289579 321619 289582
rect 70526 289444 70532 289508
rect 70596 289444 70602 289508
rect 121545 289098 121611 289101
rect 119876 289096 121611 289098
rect 67449 288554 67515 288557
rect 70166 288554 70226 289068
rect 119876 289040 121550 289096
rect 121606 289040 121611 289096
rect 119876 289038 121611 289040
rect 121545 289035 121611 289038
rect 197445 288962 197511 288965
rect 197445 288960 200100 288962
rect 197445 288904 197450 288960
rect 197506 288904 200100 288960
rect 197445 288902 200100 288904
rect 197445 288899 197511 288902
rect 67449 288552 70226 288554
rect 67449 288496 67454 288552
rect 67510 288496 70226 288552
rect 67449 288494 70226 288496
rect 67449 288491 67515 288494
rect 121453 288418 121519 288421
rect 119876 288416 121519 288418
rect 68829 288146 68895 288149
rect 70350 288146 70410 288388
rect 119876 288360 121458 288416
rect 121514 288360 121519 288416
rect 119876 288358 121519 288360
rect 121453 288355 121519 288358
rect 128854 288356 128860 288420
rect 128924 288418 128930 288420
rect 129733 288418 129799 288421
rect 181621 288418 181687 288421
rect 128924 288416 181687 288418
rect 128924 288360 129738 288416
rect 129794 288360 181626 288416
rect 181682 288360 181687 288416
rect 128924 288358 181687 288360
rect 128924 288356 128930 288358
rect 129733 288355 129799 288358
rect 181621 288355 181687 288358
rect 68829 288144 70410 288146
rect 68829 288088 68834 288144
rect 68890 288088 70410 288144
rect 68829 288086 70410 288088
rect 68829 288083 68895 288086
rect 121545 287738 121611 287741
rect 119876 287736 121611 287738
rect 67633 287194 67699 287197
rect 70166 287194 70226 287708
rect 119876 287680 121550 287736
rect 121606 287680 121611 287736
rect 119876 287678 121611 287680
rect 121545 287675 121611 287678
rect 67633 287192 70226 287194
rect 67633 287136 67638 287192
rect 67694 287136 70226 287192
rect 67633 287134 70226 287136
rect 67633 287131 67699 287134
rect 67817 287058 67883 287061
rect 69982 287058 70226 287070
rect 121453 287058 121519 287061
rect 67817 287056 70226 287058
rect 67817 287000 67822 287056
rect 67878 287010 70226 287056
rect 119876 287056 121519 287058
rect 67878 287000 70042 287010
rect 67817 286998 70042 287000
rect 119876 287000 121458 287056
rect 121514 287000 121519 287056
rect 119876 286998 121519 287000
rect 67817 286995 67883 286998
rect 121453 286995 121519 286998
rect 197445 286922 197511 286925
rect 322473 286922 322539 286925
rect 197445 286920 200100 286922
rect 197445 286864 197450 286920
rect 197506 286864 200100 286920
rect 197445 286862 200100 286864
rect 319884 286920 322539 286922
rect 319884 286864 322478 286920
rect 322534 286864 322539 286920
rect 319884 286862 322539 286864
rect 197445 286859 197511 286862
rect 322473 286859 322539 286862
rect 67725 286786 67791 286789
rect 67725 286784 70226 286786
rect 67725 286728 67730 286784
rect 67786 286728 70226 286784
rect 67725 286726 70226 286728
rect 67725 286723 67791 286726
rect 70166 286348 70226 286726
rect 121545 286378 121611 286381
rect 119876 286376 121611 286378
rect 119876 286320 121550 286376
rect 121606 286320 121611 286376
rect 119876 286318 121611 286320
rect 121545 286315 121611 286318
rect 68185 286106 68251 286109
rect 68185 286104 70226 286106
rect 68185 286048 68190 286104
rect 68246 286048 70226 286104
rect 68185 286046 70226 286048
rect 68185 286043 68251 286046
rect 70166 285668 70226 286046
rect 121637 285698 121703 285701
rect 119876 285696 121703 285698
rect 119876 285640 121642 285696
rect 121698 285640 121703 285696
rect 119876 285638 121703 285640
rect 121637 285635 121703 285638
rect 67633 285426 67699 285429
rect 67633 285424 70226 285426
rect 67633 285368 67638 285424
rect 67694 285368 70226 285424
rect 67633 285366 70226 285368
rect 67633 285363 67699 285366
rect 70166 284988 70226 285366
rect 583520 285276 584960 285516
rect 121453 285018 121519 285021
rect 322749 285018 322815 285021
rect 119876 285016 121519 285018
rect 119876 284960 121458 285016
rect 121514 284960 121519 285016
rect 119876 284958 121519 284960
rect 319884 285016 322815 285018
rect 319884 284960 322754 285016
rect 322810 284960 322815 285016
rect 319884 284958 322815 284960
rect 121453 284955 121519 284958
rect 322749 284955 322815 284958
rect 67633 284474 67699 284477
rect 67633 284472 70226 284474
rect 67633 284416 67638 284472
rect 67694 284416 70226 284472
rect 67633 284414 70226 284416
rect 67633 284411 67699 284414
rect 70166 284308 70226 284414
rect 121545 284338 121611 284341
rect 119876 284336 121611 284338
rect 119876 284280 121550 284336
rect 121606 284280 121611 284336
rect 119876 284278 121611 284280
rect 121545 284275 121611 284278
rect 197445 284202 197511 284205
rect 197445 284200 200100 284202
rect 197445 284144 197450 284200
rect 197506 284144 200100 284200
rect 197445 284142 200100 284144
rect 197445 284139 197511 284142
rect 70526 284004 70532 284068
rect 70596 284004 70602 284068
rect 70534 283628 70594 284004
rect 121453 283658 121519 283661
rect 119876 283656 121519 283658
rect 119876 283600 121458 283656
rect 121514 283600 121519 283656
rect 119876 283598 121519 283600
rect 121453 283595 121519 283598
rect 67725 283386 67791 283389
rect 67725 283384 70226 283386
rect 67725 283328 67730 283384
rect 67786 283328 70226 283384
rect 67725 283326 70226 283328
rect 67725 283323 67791 283326
rect 70166 282948 70226 283326
rect 121453 282978 121519 282981
rect 322473 282978 322539 282981
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 319884 282976 322539 282978
rect 319884 282920 322478 282976
rect 322534 282920 322539 282976
rect 319884 282918 322539 282920
rect 121453 282915 121519 282918
rect 322473 282915 322539 282918
rect 122189 282298 122255 282301
rect 119876 282296 122255 282298
rect 119876 282240 122194 282296
rect 122250 282240 122255 282296
rect 119876 282238 122255 282240
rect 122189 282235 122255 282238
rect 67633 282162 67699 282165
rect 197445 282162 197511 282165
rect 67633 282160 70226 282162
rect 67633 282104 67638 282160
rect 67694 282104 70226 282160
rect 67633 282102 70226 282104
rect 67633 282099 67699 282102
rect 70166 281588 70226 282102
rect 197445 282160 200100 282162
rect 197445 282104 197450 282160
rect 197506 282104 200100 282160
rect 197445 282102 200100 282104
rect 197445 282099 197511 282102
rect 121453 281618 121519 281621
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 121453 281555 121519 281558
rect 69105 281346 69171 281349
rect 69105 281344 70226 281346
rect 69105 281288 69110 281344
rect 69166 281288 70226 281344
rect 69105 281286 70226 281288
rect 69105 281283 69171 281286
rect 70166 280908 70226 281286
rect 121545 280938 121611 280941
rect 119876 280936 121611 280938
rect 119876 280880 121550 280936
rect 121606 280880 121611 280936
rect 119876 280878 121611 280880
rect 121545 280875 121611 280878
rect 322473 280802 322539 280805
rect 319884 280800 322539 280802
rect 319884 280744 322478 280800
rect 322534 280744 322539 280800
rect 319884 280742 322539 280744
rect 322473 280739 322539 280742
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121453 280258 121519 280261
rect 119876 280256 121519 280258
rect -960 279972 480 280212
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 121453 280195 121519 280198
rect 197445 280258 197511 280261
rect 197445 280256 200100 280258
rect 197445 280200 197450 280256
rect 197506 280200 200100 280256
rect 197445 280198 200100 280200
rect 197445 280195 197511 280198
rect 67725 279986 67791 279989
rect 67725 279984 70226 279986
rect 67725 279928 67730 279984
rect 67786 279928 70226 279984
rect 67725 279926 70226 279928
rect 67725 279923 67791 279926
rect 70166 279548 70226 279926
rect 121637 279578 121703 279581
rect 119876 279576 121703 279578
rect 119876 279520 121642 279576
rect 121698 279520 121703 279576
rect 119876 279518 121703 279520
rect 121637 279515 121703 279518
rect 67633 279306 67699 279309
rect 67633 279304 70226 279306
rect 67633 279248 67638 279304
rect 67694 279248 70226 279304
rect 67633 279246 70226 279248
rect 67633 279243 67699 279246
rect 70166 278868 70226 279246
rect 121453 278898 121519 278901
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 121453 278835 121519 278838
rect 67633 278626 67699 278629
rect 67633 278624 70226 278626
rect 67633 278568 67638 278624
rect 67694 278568 70226 278624
rect 67633 278566 70226 278568
rect 67633 278563 67699 278566
rect 70166 278188 70226 278566
rect 122741 278218 122807 278221
rect 119876 278216 122807 278218
rect 119876 278160 122746 278216
rect 122802 278160 122807 278216
rect 119876 278158 122807 278160
rect 122741 278155 122807 278158
rect 321829 278082 321895 278085
rect 319884 278080 321895 278082
rect 319884 278024 321834 278080
rect 321890 278024 321895 278080
rect 319884 278022 321895 278024
rect 321829 278019 321895 278022
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 121453 277538 121519 277541
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 121453 277475 121519 277478
rect 197445 277538 197511 277541
rect 197445 277536 200100 277538
rect 197445 277480 197450 277536
rect 197506 277480 200100 277536
rect 197445 277478 200100 277480
rect 197445 277475 197511 277478
rect 121453 276858 121519 276861
rect 119876 276856 121519 276858
rect 67725 276450 67791 276453
rect 70166 276450 70226 276828
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 119876 276798 121519 276800
rect 121453 276795 121519 276798
rect 67725 276448 70226 276450
rect 67725 276392 67730 276448
rect 67786 276392 70226 276448
rect 67725 276390 70226 276392
rect 67725 276387 67791 276390
rect 69054 276252 69060 276316
rect 69124 276314 69130 276316
rect 69124 276254 70226 276314
rect 69124 276252 69130 276254
rect 70166 276148 70226 276254
rect 121453 276178 121519 276181
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 121453 276115 121519 276118
rect 322197 276042 322263 276045
rect 319884 276040 322263 276042
rect 319884 275984 322202 276040
rect 322258 275984 322263 276040
rect 319884 275982 322263 275984
rect 322197 275979 322263 275982
rect 67633 275906 67699 275909
rect 67633 275904 70226 275906
rect 67633 275848 67638 275904
rect 67694 275848 70226 275904
rect 67633 275846 70226 275848
rect 67633 275843 67699 275846
rect 70166 275468 70226 275846
rect 120165 275498 120231 275501
rect 120717 275498 120783 275501
rect 119876 275496 120783 275498
rect 119876 275440 120170 275496
rect 120226 275440 120722 275496
rect 120778 275440 120783 275496
rect 119876 275438 120783 275440
rect 120165 275435 120231 275438
rect 120717 275435 120783 275438
rect 197445 275362 197511 275365
rect 197445 275360 200100 275362
rect 197445 275304 197450 275360
rect 197506 275304 200100 275360
rect 197445 275302 200100 275304
rect 197445 275299 197511 275302
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 121453 274818 121519 274821
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 121453 274755 121519 274758
rect 67725 274546 67791 274549
rect 67725 274544 70226 274546
rect 67725 274488 67730 274544
rect 67786 274488 70226 274544
rect 67725 274486 70226 274488
rect 67725 274483 67791 274486
rect 70166 274108 70226 274486
rect 121545 274138 121611 274141
rect 322381 274138 322447 274141
rect 119876 274136 121611 274138
rect 119876 274080 121550 274136
rect 121606 274080 121611 274136
rect 119876 274078 121611 274080
rect 319884 274136 322447 274138
rect 319884 274080 322386 274136
rect 322442 274080 322447 274136
rect 319884 274078 322447 274080
rect 121545 274075 121611 274078
rect 322381 274075 322447 274078
rect 67633 273594 67699 273597
rect 67633 273592 70226 273594
rect 67633 273536 67638 273592
rect 67694 273536 70226 273592
rect 67633 273534 70226 273536
rect 67633 273531 67699 273534
rect 70166 273428 70226 273534
rect 121453 273458 121519 273461
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 121453 273395 121519 273398
rect 197445 273322 197511 273325
rect 197445 273320 200100 273322
rect 197445 273264 197450 273320
rect 197506 273264 200100 273320
rect 197445 273262 200100 273264
rect 197445 273259 197511 273262
rect 121453 272778 121519 272781
rect 119876 272776 121519 272778
rect 67633 272370 67699 272373
rect 70166 272370 70226 272748
rect 119876 272720 121458 272776
rect 121514 272720 121519 272776
rect 119876 272718 121519 272720
rect 121453 272715 121519 272718
rect 67633 272368 70226 272370
rect 67633 272312 67638 272368
rect 67694 272312 70226 272368
rect 67633 272310 70226 272312
rect 67633 272307 67699 272310
rect 68829 272234 68895 272237
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 68829 272232 70226 272234
rect 68829 272176 68834 272232
rect 68890 272176 70226 272232
rect 68829 272174 70226 272176
rect 68829 272171 68895 272174
rect 70166 272068 70226 272174
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 122281 272098 122347 272101
rect 119876 272096 122347 272098
rect 119876 272040 122286 272096
rect 122342 272040 122347 272096
rect 583520 272084 584960 272174
rect 119876 272038 122347 272040
rect 122281 272035 122347 272038
rect 68093 271554 68159 271557
rect 68093 271552 70226 271554
rect 68093 271496 68098 271552
rect 68154 271496 70226 271552
rect 68093 271494 70226 271496
rect 68093 271491 68159 271494
rect 70166 271388 70226 271494
rect 121453 271418 121519 271421
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 121453 271355 121519 271358
rect 197445 271282 197511 271285
rect 198549 271282 198615 271285
rect 321645 271282 321711 271285
rect 197445 271280 200100 271282
rect 197445 271224 197450 271280
rect 197506 271224 198554 271280
rect 198610 271224 200100 271280
rect 197445 271222 200100 271224
rect 319884 271280 321711 271282
rect 319884 271224 321650 271280
rect 321706 271224 321711 271280
rect 319884 271222 321711 271224
rect 197445 271219 197511 271222
rect 198549 271219 198615 271222
rect 321645 271219 321711 271222
rect 67725 271146 67791 271149
rect 67725 271144 70226 271146
rect 67725 271088 67730 271144
rect 67786 271088 70226 271144
rect 67725 271086 70226 271088
rect 67725 271083 67791 271086
rect 70166 270708 70226 271086
rect 121453 270058 121519 270061
rect 119876 270056 121519 270058
rect 67633 269650 67699 269653
rect 70166 269650 70226 270028
rect 119876 270000 121458 270056
rect 121514 270000 121519 270056
rect 119876 269998 121519 270000
rect 121453 269995 121519 269998
rect 67633 269648 70226 269650
rect 67633 269592 67638 269648
rect 67694 269592 70226 269648
rect 67633 269590 70226 269592
rect 67633 269587 67699 269590
rect 69238 269452 69244 269516
rect 69308 269514 69314 269516
rect 69308 269454 70226 269514
rect 69308 269452 69314 269454
rect 70166 269348 70226 269454
rect 121453 269378 121519 269381
rect 119876 269376 121519 269378
rect 119876 269320 121458 269376
rect 121514 269320 121519 269376
rect 119876 269318 121519 269320
rect 121453 269315 121519 269318
rect 322841 269242 322907 269245
rect 319884 269240 322907 269242
rect 319884 269184 322846 269240
rect 322902 269184 322907 269240
rect 319884 269182 322907 269184
rect 322841 269179 322907 269182
rect 121545 268698 121611 268701
rect 119876 268696 121611 268698
rect 69105 268290 69171 268293
rect 70166 268290 70226 268668
rect 119876 268640 121550 268696
rect 121606 268640 121611 268696
rect 119876 268638 121611 268640
rect 121545 268635 121611 268638
rect 197445 268562 197511 268565
rect 197445 268560 200100 268562
rect 197445 268504 197450 268560
rect 197506 268504 200100 268560
rect 197445 268502 200100 268504
rect 197445 268499 197511 268502
rect 69105 268288 70226 268290
rect 69105 268232 69110 268288
rect 69166 268232 70226 268288
rect 69105 268230 70226 268232
rect 69105 268227 69171 268230
rect 67633 268154 67699 268157
rect 67633 268152 70226 268154
rect 67633 268096 67638 268152
rect 67694 268096 70226 268152
rect 67633 268094 70226 268096
rect 67633 268091 67699 268094
rect 70166 267988 70226 268094
rect 121453 268018 121519 268021
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 121453 267955 121519 267958
rect 121545 267338 121611 267341
rect 322473 267338 322539 267341
rect 119876 267336 121611 267338
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 67633 267066 67699 267069
rect 70166 267066 70226 267308
rect 119876 267280 121550 267336
rect 121606 267280 121611 267336
rect 119876 267278 121611 267280
rect 319884 267336 322539 267338
rect 319884 267280 322478 267336
rect 322534 267280 322539 267336
rect 319884 267278 322539 267280
rect 121545 267275 121611 267278
rect 322473 267275 322539 267278
rect 67633 267064 70226 267066
rect 67633 267008 67638 267064
rect 67694 267008 70226 267064
rect 67633 267006 70226 267008
rect 67633 267003 67699 267006
rect 123334 267004 123340 267068
rect 123404 267066 123410 267068
rect 179413 267066 179479 267069
rect 123404 267064 179479 267066
rect 123404 267008 179418 267064
rect 179474 267008 179479 267064
rect 123404 267006 179479 267008
rect 123404 267004 123410 267006
rect 179413 267003 179479 267006
rect 67725 266930 67791 266933
rect 67725 266928 70226 266930
rect 67725 266872 67730 266928
rect 67786 266872 70226 266928
rect 67725 266870 70226 266872
rect 67725 266867 67791 266870
rect 70166 266628 70226 266870
rect 121453 266658 121519 266661
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 121453 266595 121519 266598
rect 197353 266522 197419 266525
rect 197353 266520 200100 266522
rect 197353 266464 197358 266520
rect 197414 266464 200100 266520
rect 197353 266462 200100 266464
rect 197353 266459 197419 266462
rect 68737 266250 68803 266253
rect 68737 266248 70226 266250
rect 68737 266192 68742 266248
rect 68798 266192 70226 266248
rect 68737 266190 70226 266192
rect 68737 266187 68803 266190
rect 70166 265948 70226 266190
rect 121545 265978 121611 265981
rect 119876 265976 121611 265978
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 121545 265915 121611 265918
rect 67633 265706 67699 265709
rect 67633 265704 70226 265706
rect 67633 265648 67638 265704
rect 67694 265648 70226 265704
rect 67633 265646 70226 265648
rect 67633 265643 67699 265646
rect 70166 265268 70226 265646
rect 121453 265298 121519 265301
rect 119876 265296 121519 265298
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 121453 265235 121519 265238
rect 322473 265162 322539 265165
rect 319884 265160 322539 265162
rect 319884 265104 322478 265160
rect 322534 265104 322539 265160
rect 319884 265102 322539 265104
rect 322473 265099 322539 265102
rect 121453 264618 121519 264621
rect 119876 264616 121519 264618
rect 67725 264210 67791 264213
rect 70166 264210 70226 264588
rect 119876 264560 121458 264616
rect 121514 264560 121519 264616
rect 119876 264558 121519 264560
rect 121453 264555 121519 264558
rect 197353 264482 197419 264485
rect 197353 264480 200100 264482
rect 197353 264424 197358 264480
rect 197414 264424 200100 264480
rect 197353 264422 200100 264424
rect 197353 264419 197419 264422
rect 67725 264208 70226 264210
rect 67725 264152 67730 264208
rect 67786 264152 70226 264208
rect 67725 264150 70226 264152
rect 67725 264147 67791 264150
rect 121453 263938 121519 263941
rect 119876 263936 121519 263938
rect 67633 263666 67699 263669
rect 70350 263666 70410 263908
rect 119876 263880 121458 263936
rect 121514 263880 121519 263936
rect 119876 263878 121519 263880
rect 121453 263875 121519 263878
rect 67633 263664 70410 263666
rect 67633 263608 67638 263664
rect 67694 263608 70410 263664
rect 67633 263606 70410 263608
rect 67633 263603 67699 263606
rect 67633 263530 67699 263533
rect 67633 263528 70226 263530
rect 67633 263472 67638 263528
rect 67694 263472 70226 263528
rect 67633 263470 70226 263472
rect 67633 263467 67699 263470
rect 70166 263228 70226 263470
rect 121453 263258 121519 263261
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 121453 263195 121519 263198
rect 121545 262578 121611 262581
rect 119876 262576 121611 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121550 262576
rect 121606 262520 121611 262576
rect 119876 262518 121611 262520
rect 121545 262515 121611 262518
rect 322473 262442 322539 262445
rect 319884 262440 322539 262442
rect 319884 262384 322478 262440
rect 322534 262384 322539 262440
rect 319884 262382 322539 262384
rect 322473 262379 322539 262382
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121453 261898 121519 261901
rect 119876 261896 121519 261898
rect 67725 261490 67791 261493
rect 70166 261490 70226 261868
rect 119876 261840 121458 261896
rect 121514 261840 121519 261896
rect 119876 261838 121519 261840
rect 121453 261835 121519 261838
rect 197353 261762 197419 261765
rect 197353 261760 200100 261762
rect 197353 261704 197358 261760
rect 197414 261704 200100 261760
rect 197353 261702 200100 261704
rect 197353 261699 197419 261702
rect 67725 261488 70226 261490
rect 67725 261432 67730 261488
rect 67786 261432 70226 261488
rect 67725 261430 70226 261432
rect 67725 261427 67791 261430
rect 67817 261354 67883 261357
rect 67817 261352 70226 261354
rect 67817 261296 67822 261352
rect 67878 261296 70226 261352
rect 67817 261294 70226 261296
rect 67817 261291 67883 261294
rect 70166 261188 70226 261294
rect 121545 261218 121611 261221
rect 119876 261216 121611 261218
rect 119876 261160 121550 261216
rect 121606 261160 121611 261216
rect 119876 261158 121611 261160
rect 121545 261155 121611 261158
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121453 260538 121519 260541
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 121453 260475 121519 260478
rect 322473 260402 322539 260405
rect 319884 260400 322539 260402
rect 319884 260344 322478 260400
rect 322534 260344 322539 260400
rect 319884 260342 322539 260344
rect 322473 260339 322539 260342
rect 69197 260266 69263 260269
rect 69197 260264 70226 260266
rect 69197 260208 69202 260264
rect 69258 260208 70226 260264
rect 69197 260206 70226 260208
rect 69197 260203 69263 260206
rect 70166 259828 70226 260206
rect 121453 259858 121519 259861
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 121453 259795 121519 259798
rect 197353 259722 197419 259725
rect 197353 259720 200100 259722
rect 197353 259664 197358 259720
rect 197414 259664 200100 259720
rect 197353 259662 200100 259664
rect 197353 259659 197419 259662
rect 121637 259178 121703 259181
rect 119876 259176 121703 259178
rect 67633 258634 67699 258637
rect 70166 258634 70226 259148
rect 119876 259120 121642 259176
rect 121698 259120 121703 259176
rect 119876 259118 121703 259120
rect 121637 259115 121703 259118
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect 67633 258632 70226 258634
rect 67633 258576 67638 258632
rect 67694 258576 70226 258632
rect 67633 258574 70226 258576
rect 67633 258571 67699 258574
rect 121545 258498 121611 258501
rect 119876 258496 121611 258498
rect 67725 258226 67791 258229
rect 70350 258226 70410 258468
rect 119876 258440 121550 258496
rect 121606 258440 121611 258496
rect 119876 258438 121611 258440
rect 121545 258435 121611 258438
rect 322841 258362 322907 258365
rect 319884 258360 322907 258362
rect 319884 258304 322846 258360
rect 322902 258304 322907 258360
rect 319884 258302 322907 258304
rect 322841 258299 322907 258302
rect 67725 258224 70410 258226
rect 67725 258168 67730 258224
rect 67786 258168 70410 258224
rect 67725 258166 70410 258168
rect 67725 258163 67791 258166
rect 67633 257954 67699 257957
rect 67633 257952 70226 257954
rect 67633 257896 67638 257952
rect 67694 257896 70226 257952
rect 67633 257894 70226 257896
rect 67633 257891 67699 257894
rect 70166 257788 70226 257894
rect 121545 257818 121611 257821
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 121545 257755 121611 257758
rect 197353 257682 197419 257685
rect 197353 257680 200100 257682
rect 197353 257624 197358 257680
rect 197414 257624 200100 257680
rect 197353 257622 200100 257624
rect 197353 257619 197419 257622
rect 121453 257138 121519 257141
rect 119876 257136 121519 257138
rect 67633 256866 67699 256869
rect 70350 256866 70410 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 121453 257075 121519 257078
rect 67633 256864 70410 256866
rect 67633 256808 67638 256864
rect 67694 256808 70410 256864
rect 67633 256806 70410 256808
rect 67633 256803 67699 256806
rect 133086 256668 133092 256732
rect 133156 256730 133162 256732
rect 133873 256730 133939 256733
rect 133156 256728 133939 256730
rect 133156 256672 133878 256728
rect 133934 256672 133939 256728
rect 133156 256670 133939 256672
rect 133156 256668 133162 256670
rect 133873 256667 133939 256670
rect 68737 255914 68803 255917
rect 70166 255914 70226 256428
rect 68737 255912 70226 255914
rect 68737 255856 68742 255912
rect 68798 255856 70226 255912
rect 68737 255854 70226 255856
rect 119846 255914 119906 256428
rect 128854 255914 128860 255916
rect 119846 255854 128860 255914
rect 68737 255851 68803 255854
rect 128854 255852 128860 255854
rect 128924 255852 128930 255916
rect 121453 255778 121519 255781
rect 119876 255776 121519 255778
rect 67633 255370 67699 255373
rect 70166 255370 70226 255748
rect 119876 255720 121458 255776
rect 121514 255720 121519 255776
rect 119876 255718 121519 255720
rect 121453 255715 121519 255718
rect 197353 255642 197419 255645
rect 321829 255642 321895 255645
rect 197353 255640 200100 255642
rect 197353 255584 197358 255640
rect 197414 255584 200100 255640
rect 197353 255582 200100 255584
rect 319884 255640 321895 255642
rect 319884 255584 321834 255640
rect 321890 255584 321895 255640
rect 319884 255582 321895 255584
rect 197353 255579 197419 255582
rect 321829 255579 321895 255582
rect 67633 255368 70226 255370
rect 67633 255312 67638 255368
rect 67694 255312 70226 255368
rect 67633 255310 70226 255312
rect 67633 255307 67699 255310
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 121453 255098 121519 255101
rect 119876 255096 121519 255098
rect 119876 255040 121458 255096
rect 121514 255040 121519 255096
rect 119876 255038 121519 255040
rect 121453 255035 121519 255038
rect 67725 254826 67791 254829
rect 67725 254824 70226 254826
rect 67725 254768 67730 254824
rect 67786 254768 70226 254824
rect 67725 254766 70226 254768
rect 67725 254763 67791 254766
rect 70166 254388 70226 254766
rect 122097 254418 122163 254421
rect 119876 254416 122163 254418
rect 119876 254360 122102 254416
rect 122158 254360 122163 254416
rect 119876 254358 122163 254360
rect 122097 254355 122163 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 67633 253874 67699 253877
rect 67633 253872 70226 253874
rect 67633 253816 67638 253872
rect 67694 253816 70226 253872
rect 67633 253814 70226 253816
rect 67633 253811 67699 253814
rect 70166 253708 70226 253814
rect 122189 253738 122255 253741
rect 119876 253736 122255 253738
rect 119876 253680 122194 253736
rect 122250 253680 122255 253736
rect 119876 253678 122255 253680
rect 122189 253675 122255 253678
rect 322841 253602 322907 253605
rect 319884 253600 322907 253602
rect 319884 253544 322846 253600
rect 322902 253544 322907 253600
rect 319884 253542 322907 253544
rect 322841 253539 322907 253542
rect 67725 253466 67791 253469
rect 67725 253464 70226 253466
rect 67725 253408 67730 253464
rect 67786 253408 70226 253464
rect 67725 253406 70226 253408
rect 67725 253403 67791 253406
rect 70166 253028 70226 253406
rect 121453 253058 121519 253061
rect 119876 253056 121519 253058
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 121453 252995 121519 252998
rect 197353 252922 197419 252925
rect 197353 252920 200100 252922
rect 197353 252864 197358 252920
rect 197414 252864 200100 252920
rect 197353 252862 200100 252864
rect 197353 252859 197419 252862
rect 197118 252452 197124 252516
rect 197188 252514 197194 252516
rect 197445 252514 197511 252517
rect 197188 252512 197511 252514
rect 197188 252456 197450 252512
rect 197506 252456 197511 252512
rect 197188 252454 197511 252456
rect 197188 252452 197194 252454
rect 197445 252451 197511 252454
rect 121453 252378 121519 252381
rect 119876 252376 121519 252378
rect 69197 251834 69263 251837
rect 70166 251834 70226 252348
rect 119876 252320 121458 252376
rect 121514 252320 121519 252376
rect 119876 252318 121519 252320
rect 121453 252315 121519 252318
rect 69197 251832 70226 251834
rect 69197 251776 69202 251832
rect 69258 251776 70226 251832
rect 69197 251774 70226 251776
rect 69197 251771 69263 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 68921 251426 68987 251429
rect 70350 251426 70410 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 323577 251562 323643 251565
rect 319884 251560 323643 251562
rect 319884 251504 323582 251560
rect 323638 251504 323643 251560
rect 319884 251502 323643 251504
rect 323577 251499 323643 251502
rect 68921 251424 70410 251426
rect 68921 251368 68926 251424
rect 68982 251368 70410 251424
rect 68921 251366 70410 251368
rect 68921 251363 68987 251366
rect 130561 251290 130627 251293
rect 192334 251290 192340 251292
rect 130561 251288 192340 251290
rect 130561 251232 130566 251288
rect 130622 251232 192340 251288
rect 130561 251230 192340 251232
rect 130561 251227 130627 251230
rect 192334 251228 192340 251230
rect 192404 251290 192410 251292
rect 192845 251290 192911 251293
rect 192404 251288 192911 251290
rect 192404 251232 192850 251288
rect 192906 251232 192911 251288
rect 192404 251230 192911 251232
rect 192404 251228 192410 251230
rect 192845 251227 192911 251230
rect 67633 251154 67699 251157
rect 119797 251154 119863 251157
rect 67633 251152 70226 251154
rect 67633 251096 67638 251152
rect 67694 251096 70226 251152
rect 67633 251094 70226 251096
rect 67633 251091 67699 251094
rect 70166 250988 70226 251094
rect 119797 251152 119906 251154
rect 119797 251096 119802 251152
rect 119858 251096 119906 251152
rect 119797 251091 119906 251096
rect 119846 251018 119906 251091
rect 120165 251018 120231 251021
rect 119846 251016 120231 251018
rect 119846 250988 120170 251016
rect 119876 250960 120170 250988
rect 120226 250960 120231 251016
rect 119876 250958 120231 250960
rect 120165 250955 120231 250958
rect 197353 250882 197419 250885
rect 197353 250880 200100 250882
rect 197353 250824 197358 250880
rect 197414 250824 200100 250880
rect 197353 250822 200100 250824
rect 197353 250819 197419 250822
rect 121453 250338 121519 250341
rect 119876 250336 121519 250338
rect 68553 249930 68619 249933
rect 70166 249930 70226 250308
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 121453 250275 121519 250278
rect 68553 249928 70226 249930
rect 68553 249872 68558 249928
rect 68614 249872 70226 249928
rect 68553 249870 70226 249872
rect 68553 249867 68619 249870
rect 121545 249658 121611 249661
rect 119876 249656 121611 249658
rect 67633 249114 67699 249117
rect 70166 249114 70226 249628
rect 119876 249600 121550 249656
rect 121606 249600 121611 249656
rect 119876 249598 121611 249600
rect 121545 249595 121611 249598
rect 67633 249112 70226 249114
rect 67633 249056 67638 249112
rect 67694 249056 70226 249112
rect 67633 249054 70226 249056
rect 67633 249051 67699 249054
rect 121453 248978 121519 248981
rect 119876 248976 121519 248978
rect 68369 248706 68435 248709
rect 70166 248706 70226 248948
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 121453 248915 121519 248918
rect 197353 248978 197419 248981
rect 197353 248976 200100 248978
rect 197353 248920 197358 248976
rect 197414 248920 200100 248976
rect 197353 248918 200100 248920
rect 197353 248915 197419 248918
rect 322473 248842 322539 248845
rect 319884 248840 322539 248842
rect 319884 248784 322478 248840
rect 322534 248784 322539 248840
rect 319884 248782 322539 248784
rect 322473 248779 322539 248782
rect 68369 248704 70226 248706
rect 68369 248648 68374 248704
rect 68430 248648 70226 248704
rect 68369 248646 70226 248648
rect 68369 248643 68435 248646
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67633 247754 67699 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67633 247752 70226 247754
rect 67633 247696 67638 247752
rect 67694 247696 70226 247752
rect 67633 247694 70226 247696
rect 67633 247691 67699 247694
rect 119286 247692 119292 247756
rect 119356 247754 119362 247756
rect 119356 247694 119906 247754
rect 119356 247692 119362 247694
rect 119846 247618 119906 247694
rect 121545 247618 121611 247621
rect 119846 247616 121611 247618
rect 119846 247588 121550 247616
rect 69841 247074 69907 247077
rect 70166 247074 70226 247588
rect 119876 247560 121550 247588
rect 121606 247560 121611 247616
rect 119876 247558 121611 247560
rect 121545 247555 121611 247558
rect 69841 247072 70226 247074
rect 69841 247016 69846 247072
rect 69902 247016 70226 247072
rect 69841 247014 70226 247016
rect 69841 247011 69907 247014
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 67357 246394 67423 246397
rect 70166 246396 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 322473 246802 322539 246805
rect 319884 246800 322539 246802
rect 319884 246744 322478 246800
rect 322534 246744 322539 246800
rect 319884 246742 322539 246744
rect 322473 246739 322539 246742
rect 70158 246394 70164 246396
rect 67357 246392 70164 246394
rect 67357 246336 67362 246392
rect 67418 246336 70164 246392
rect 67357 246334 70164 246336
rect 67357 246331 67423 246334
rect 70158 246332 70164 246334
rect 70228 246332 70234 246396
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 67541 245714 67607 245717
rect 70166 245714 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 198089 246122 198155 246125
rect 198089 246120 200100 246122
rect 198089 246064 198094 246120
rect 198150 246064 200100 246120
rect 198089 246062 200100 246064
rect 198089 246059 198155 246062
rect 67541 245712 70226 245714
rect 67541 245656 67546 245712
rect 67602 245656 70226 245712
rect 67541 245654 70226 245656
rect 67541 245651 67607 245654
rect 121545 245578 121611 245581
rect 119876 245576 121611 245578
rect 67633 245306 67699 245309
rect 70350 245306 70410 245548
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 121545 245515 121611 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 120022 245306 120028 245308
rect 67633 245304 70410 245306
rect 67633 245248 67638 245304
rect 67694 245248 70410 245304
rect 67633 245246 70410 245248
rect 119846 245246 120028 245306
rect 67633 245243 67699 245246
rect 119846 244868 119906 245246
rect 120022 245244 120028 245246
rect 120092 245244 120098 245308
rect 67357 244354 67423 244357
rect 70166 244354 70226 244868
rect 321737 244762 321803 244765
rect 319884 244760 321803 244762
rect 319884 244732 321742 244760
rect 319854 244704 321742 244732
rect 321798 244704 321803 244760
rect 319854 244702 321803 244704
rect 67357 244352 70226 244354
rect 67357 244296 67362 244352
rect 67418 244296 70226 244352
rect 67357 244294 70226 244296
rect 319345 244354 319411 244357
rect 319854 244354 319914 244702
rect 321737 244699 321803 244702
rect 319345 244352 319914 244354
rect 319345 244296 319350 244352
rect 319406 244296 319914 244352
rect 319345 244294 319914 244296
rect 67357 244291 67423 244294
rect 319345 244291 319411 244294
rect 121545 244218 121611 244221
rect 119876 244216 121611 244218
rect 67633 243810 67699 243813
rect 70350 243810 70410 244188
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 121545 244155 121611 244158
rect 198273 244082 198339 244085
rect 198273 244080 200100 244082
rect 198273 244024 198278 244080
rect 198334 244024 200100 244080
rect 198273 244022 200100 244024
rect 198273 244019 198339 244022
rect 67633 243808 70410 243810
rect 67633 243752 67638 243808
rect 67694 243752 70410 243808
rect 67633 243750 70410 243752
rect 67633 243747 67699 243750
rect 67725 243674 67791 243677
rect 67725 243672 70226 243674
rect 67725 243616 67730 243672
rect 67786 243616 70226 243672
rect 67725 243614 70226 243616
rect 67725 243611 67791 243614
rect 70166 243508 70226 243614
rect 121453 243538 121519 243541
rect 119876 243536 121519 243538
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 121453 243475 121519 243478
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70534 242452 70594 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 140681 242858 140747 242861
rect 140814 242858 140820 242860
rect 140681 242856 140820 242858
rect 140681 242800 140686 242856
rect 140742 242800 140820 242856
rect 140681 242798 140820 242800
rect 140681 242795 140747 242798
rect 140814 242796 140820 242798
rect 140884 242796 140890 242860
rect 320357 242858 320423 242861
rect 321461 242858 321527 242861
rect 319884 242856 321527 242858
rect 319884 242800 320362 242856
rect 320418 242800 321466 242856
rect 321522 242800 321527 242856
rect 319884 242798 321527 242800
rect 320357 242795 320423 242798
rect 321461 242795 321527 242798
rect 70526 242388 70532 242452
rect 70596 242388 70602 242452
rect 121453 242178 121519 242181
rect 119876 242176 121519 242178
rect 70534 241636 70594 242148
rect 119876 242120 121458 242176
rect 121514 242120 121519 242176
rect 119876 242118 121519 242120
rect 121453 242115 121519 242118
rect 196566 242116 196572 242180
rect 196636 242178 196642 242180
rect 196801 242178 196867 242181
rect 196636 242176 200100 242178
rect 196636 242120 196806 242176
rect 196862 242120 200100 242176
rect 196636 242118 200100 242120
rect 196636 242116 196642 242118
rect 196801 242115 196867 242118
rect 70526 241572 70532 241636
rect 70596 241572 70602 241636
rect 120073 241498 120139 241501
rect 119876 241496 120139 241498
rect 119876 241468 120078 241496
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 70350 240956 70410 241468
rect 119846 241440 120078 241468
rect 120134 241440 120139 241496
rect 119846 241438 120139 241440
rect 119846 241226 119906 241438
rect 120073 241435 120139 241438
rect 120022 241226 120028 241228
rect 119846 241166 120028 241226
rect 120022 241164 120028 241166
rect 120092 241164 120098 241228
rect 70342 240892 70348 240956
rect 70412 240892 70418 240956
rect 121453 240818 121519 240821
rect 529933 240818 529999 240821
rect 580257 240818 580323 240821
rect 119876 240816 121519 240818
rect 69054 240212 69060 240276
rect 69124 240274 69130 240276
rect 70166 240274 70226 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 528510 240816 580323 240818
rect 528510 240760 529938 240816
rect 529994 240760 580262 240816
rect 580318 240760 580323 240816
rect 528510 240758 580323 240760
rect 320030 240348 320036 240412
rect 320100 240410 320106 240412
rect 528510 240410 528570 240758
rect 529933 240755 529999 240758
rect 580257 240755 580323 240758
rect 320100 240350 528570 240410
rect 320100 240348 320106 240350
rect 69124 240214 70226 240274
rect 195697 240274 195763 240277
rect 200614 240274 200620 240276
rect 195697 240272 200620 240274
rect 195697 240216 195702 240272
rect 195758 240216 200620 240272
rect 195697 240214 200620 240216
rect 69124 240212 69130 240214
rect 195697 240211 195763 240214
rect 200614 240212 200620 240214
rect 200684 240212 200690 240276
rect 121453 240138 121519 240141
rect 119876 240136 121519 240138
rect 119876 240080 121458 240136
rect 121514 240080 121519 240136
rect 119876 240078 121519 240080
rect 121453 240075 121519 240078
rect 320081 240002 320147 240005
rect 319884 240000 320147 240002
rect 319884 239944 320086 240000
rect 320142 239944 320147 240000
rect 319884 239942 320147 239944
rect 320081 239939 320147 239942
rect 70158 239804 70164 239868
rect 70228 239866 70234 239868
rect 72417 239866 72483 239869
rect 70228 239864 72483 239866
rect 70228 239808 72422 239864
rect 72478 239808 72483 239864
rect 70228 239806 72483 239808
rect 70228 239804 70234 239806
rect 72417 239803 72483 239806
rect 120717 239866 120783 239869
rect 320817 239866 320883 239869
rect 120717 239864 320883 239866
rect 120717 239808 120722 239864
rect 120778 239808 320822 239864
rect 320878 239808 320883 239864
rect 120717 239806 320883 239808
rect 120717 239803 120783 239806
rect 320817 239803 320883 239806
rect 117037 239730 117103 239733
rect 124806 239730 124812 239732
rect 117037 239728 124812 239730
rect 117037 239672 117042 239728
rect 117098 239672 124812 239728
rect 117037 239670 124812 239672
rect 117037 239667 117103 239670
rect 124806 239668 124812 239670
rect 124876 239668 124882 239732
rect 195881 239730 195947 239733
rect 200941 239730 201007 239733
rect 195881 239728 201007 239730
rect 195881 239672 195886 239728
rect 195942 239672 200946 239728
rect 201002 239672 201007 239728
rect 195881 239670 201007 239672
rect 195881 239667 195947 239670
rect 200941 239667 201007 239670
rect 155401 238778 155467 238781
rect 210233 238778 210299 238781
rect 155401 238776 210299 238778
rect 155401 238720 155406 238776
rect 155462 238720 210238 238776
rect 210294 238720 210299 238776
rect 155401 238718 210299 238720
rect 155401 238715 155467 238718
rect 210233 238715 210299 238718
rect 70342 238580 70348 238644
rect 70412 238642 70418 238644
rect 129774 238642 129780 238644
rect 70412 238582 129780 238642
rect 70412 238580 70418 238582
rect 129774 238580 129780 238582
rect 129844 238580 129850 238644
rect 146293 238642 146359 238645
rect 305637 238642 305703 238645
rect 146293 238640 305703 238642
rect 146293 238584 146298 238640
rect 146354 238584 305642 238640
rect 305698 238584 305703 238640
rect 146293 238582 305703 238584
rect 146293 238579 146359 238582
rect 305637 238579 305703 238582
rect 176101 238506 176167 238509
rect 201585 238506 201651 238509
rect 176101 238504 201651 238506
rect 176101 238448 176106 238504
rect 176162 238448 201590 238504
rect 201646 238448 201651 238504
rect 176101 238446 201651 238448
rect 176101 238443 176167 238446
rect 201585 238443 201651 238446
rect 299197 238506 299263 238509
rect 320030 238506 320036 238508
rect 299197 238504 320036 238506
rect 299197 238448 299202 238504
rect 299258 238448 320036 238504
rect 299197 238446 320036 238448
rect 299197 238443 299263 238446
rect 320030 238444 320036 238446
rect 320100 238444 320106 238508
rect 190361 237962 190427 237965
rect 203517 237962 203583 237965
rect 190361 237960 203583 237962
rect 190361 237904 190366 237960
rect 190422 237904 203522 237960
rect 203578 237904 203583 237960
rect 190361 237902 203583 237904
rect 190361 237899 190427 237902
rect 203517 237899 203583 237902
rect 71078 237220 71084 237284
rect 71148 237282 71154 237284
rect 126329 237282 126395 237285
rect 71148 237280 126395 237282
rect 71148 237224 126334 237280
rect 126390 237224 126395 237280
rect 71148 237222 126395 237224
rect 71148 237220 71154 237222
rect 126329 237219 126395 237222
rect 169201 237282 169267 237285
rect 324497 237282 324563 237285
rect 169201 237280 324563 237282
rect 169201 237224 169206 237280
rect 169262 237224 324502 237280
rect 324558 237224 324563 237280
rect 169201 237222 324563 237224
rect 169201 237219 169267 237222
rect 324497 237219 324563 237222
rect 107377 237146 107443 237149
rect 125726 237146 125732 237148
rect 107377 237144 125732 237146
rect 107377 237088 107382 237144
rect 107438 237088 125732 237144
rect 107377 237086 125732 237088
rect 107377 237083 107443 237086
rect 125726 237084 125732 237086
rect 125796 237084 125802 237148
rect 195973 236738 196039 236741
rect 211889 236738 211955 236741
rect 195973 236736 211955 236738
rect 195973 236680 195978 236736
rect 196034 236680 211894 236736
rect 211950 236680 211955 236736
rect 195973 236678 211955 236680
rect 195973 236675 196039 236678
rect 211889 236675 211955 236678
rect 195053 236602 195119 236605
rect 304901 236602 304967 236605
rect 321502 236602 321508 236604
rect 195053 236600 321508 236602
rect 195053 236544 195058 236600
rect 195114 236544 304906 236600
rect 304962 236544 321508 236600
rect 195053 236542 321508 236544
rect 195053 236539 195119 236542
rect 304901 236539 304967 236542
rect 321502 236540 321508 236542
rect 321572 236540 321578 236604
rect 195881 236058 195947 236061
rect 196566 236058 196572 236060
rect 195881 236056 196572 236058
rect 195881 236000 195886 236056
rect 195942 236000 196572 236056
rect 195881 235998 196572 236000
rect 195881 235995 195947 235998
rect 196566 235996 196572 235998
rect 196636 235996 196642 236060
rect 57830 235860 57836 235924
rect 57900 235922 57906 235924
rect 98361 235922 98427 235925
rect 57900 235920 98427 235922
rect 57900 235864 98366 235920
rect 98422 235864 98427 235920
rect 57900 235862 98427 235864
rect 57900 235860 57906 235862
rect 98361 235859 98427 235862
rect 106733 235922 106799 235925
rect 123661 235922 123727 235925
rect 106733 235920 123727 235922
rect 106733 235864 106738 235920
rect 106794 235864 123666 235920
rect 123722 235864 123727 235920
rect 106733 235862 123727 235864
rect 106733 235859 106799 235862
rect 123661 235859 123727 235862
rect 155309 235922 155375 235925
rect 227069 235922 227135 235925
rect 155309 235920 227135 235922
rect 155309 235864 155314 235920
rect 155370 235864 227074 235920
rect 227130 235864 227135 235920
rect 155309 235862 227135 235864
rect 155309 235859 155375 235862
rect 227069 235859 227135 235862
rect 195145 235242 195211 235245
rect 324313 235242 324379 235245
rect 195145 235240 324379 235242
rect 195145 235184 195150 235240
rect 195206 235184 324318 235240
rect 324374 235184 324379 235240
rect 195145 235182 324379 235184
rect 195145 235179 195211 235182
rect 324313 235179 324379 235182
rect 86125 234562 86191 234565
rect 324589 234562 324655 234565
rect 86125 234560 324655 234562
rect 86125 234504 86130 234560
rect 86186 234504 324594 234560
rect 324650 234504 324655 234560
rect 86125 234502 324655 234504
rect 86125 234499 86191 234502
rect 324589 234499 324655 234502
rect 140681 234426 140747 234429
rect 244457 234426 244523 234429
rect 140681 234424 244523 234426
rect 140681 234368 140686 234424
rect 140742 234368 244462 234424
rect 244518 234368 244523 234424
rect 140681 234366 244523 234368
rect 140681 234363 140747 234366
rect 244457 234363 244523 234366
rect 193121 233882 193187 233885
rect 206277 233882 206343 233885
rect 193121 233880 206343 233882
rect 193121 233824 193126 233880
rect 193182 233824 206282 233880
rect 206338 233824 206343 233880
rect 193121 233822 206343 233824
rect 193121 233819 193187 233822
rect 206277 233819 206343 233822
rect 129774 233140 129780 233204
rect 129844 233202 129850 233204
rect 289445 233202 289511 233205
rect 129844 233200 289511 233202
rect 129844 233144 289450 233200
rect 289506 233144 289511 233200
rect 129844 233142 289511 233144
rect 129844 233140 129850 233142
rect 289445 233139 289511 233142
rect 75821 233066 75887 233069
rect 137134 233066 137140 233068
rect 75821 233064 137140 233066
rect 75821 233008 75826 233064
rect 75882 233008 137140 233064
rect 75821 233006 137140 233008
rect 75821 233003 75887 233006
rect 137134 233004 137140 233006
rect 137204 233004 137210 233068
rect 122741 232522 122807 232525
rect 328494 232522 328500 232524
rect 122741 232520 328500 232522
rect 122741 232464 122746 232520
rect 122802 232464 328500 232520
rect 122741 232462 328500 232464
rect 122741 232459 122807 232462
rect 328494 232460 328500 232462
rect 328564 232460 328570 232524
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 68829 231162 68895 231165
rect 255262 231162 255268 231164
rect 68829 231160 255268 231162
rect 68829 231104 68834 231160
rect 68890 231104 255268 231160
rect 68829 231102 255268 231104
rect 68829 231099 68895 231102
rect 255262 231100 255268 231102
rect 255332 231100 255338 231164
rect 161013 230482 161079 230485
rect 320357 230482 320423 230485
rect 161013 230480 320423 230482
rect 161013 230424 161018 230480
rect 161074 230424 320362 230480
rect 320418 230424 320423 230480
rect 161013 230422 320423 230424
rect 161013 230419 161079 230422
rect 320357 230419 320423 230422
rect 69054 228924 69060 228988
rect 69124 228986 69130 228988
rect 255957 228986 256023 228989
rect 69124 228984 256023 228986
rect 69124 228928 255962 228984
rect 256018 228928 256023 228984
rect 69124 228926 256023 228928
rect 69124 228924 69130 228926
rect 255957 228923 256023 228926
rect 192334 228244 192340 228308
rect 192404 228306 192410 228308
rect 216121 228306 216187 228309
rect 192404 228304 216187 228306
rect 192404 228248 216126 228304
rect 216182 228248 216187 228304
rect 192404 228246 216187 228248
rect 192404 228244 192410 228246
rect 216121 228243 216187 228246
rect -960 227884 480 228124
rect 151169 227626 151235 227629
rect 324405 227626 324471 227629
rect 151169 227624 324471 227626
rect 151169 227568 151174 227624
rect 151230 227568 324410 227624
rect 324466 227568 324471 227624
rect 151169 227566 324471 227568
rect 151169 227563 151235 227566
rect 324405 227563 324471 227566
rect 126329 226266 126395 226269
rect 292021 226266 292087 226269
rect 126329 226264 292087 226266
rect 126329 226208 126334 226264
rect 126390 226208 292026 226264
rect 292082 226208 292087 226264
rect 126329 226206 292087 226208
rect 126329 226203 126395 226206
rect 292021 226203 292087 226206
rect 321502 224436 321508 224500
rect 321572 224498 321578 224500
rect 321645 224498 321711 224501
rect 321572 224496 321711 224498
rect 321572 224440 321650 224496
rect 321706 224440 321711 224496
rect 321572 224438 321711 224440
rect 321572 224436 321578 224438
rect 321645 224435 321711 224438
rect 211889 224226 211955 224229
rect 499849 224226 499915 224229
rect 211889 224224 499915 224226
rect 211889 224168 211894 224224
rect 211950 224168 499854 224224
rect 499910 224168 499915 224224
rect 211889 224166 499915 224168
rect 211889 224163 211955 224166
rect 499849 224163 499915 224166
rect 164877 222866 164943 222869
rect 353385 222866 353451 222869
rect 164877 222864 353451 222866
rect 164877 222808 164882 222864
rect 164938 222808 353390 222864
rect 353446 222808 353451 222864
rect 164877 222806 353451 222808
rect 164877 222803 164943 222806
rect 353385 222803 353451 222806
rect 178534 221444 178540 221508
rect 178604 221506 178610 221508
rect 362953 221506 363019 221509
rect 178604 221504 363019 221506
rect 178604 221448 362958 221504
rect 363014 221448 363019 221504
rect 178604 221446 363019 221448
rect 178604 221444 178610 221446
rect 362953 221443 363019 221446
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 1301 217290 1367 217293
rect 120022 217290 120028 217292
rect 1301 217288 120028 217290
rect 1301 217232 1306 217288
rect 1362 217232 120028 217288
rect 1301 217230 120028 217232
rect 1301 217227 1367 217230
rect 120022 217228 120028 217230
rect 120092 217228 120098 217292
rect 160686 215868 160692 215932
rect 160756 215930 160762 215932
rect 268326 215930 268332 215932
rect 160756 215870 268332 215930
rect 160756 215868 160762 215870
rect 268326 215868 268332 215870
rect 268396 215868 268402 215932
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 52177 206274 52243 206277
rect 263542 206274 263548 206276
rect 52177 206272 263548 206274
rect 52177 206216 52182 206272
rect 52238 206216 263548 206272
rect 52177 206214 263548 206216
rect 52177 206211 52243 206214
rect 263542 206212 263548 206214
rect 263612 206212 263618 206276
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 173157 204914 173223 204917
rect 258574 204914 258580 204916
rect 173157 204912 258580 204914
rect 173157 204856 173162 204912
rect 173218 204856 258580 204912
rect 173157 204854 258580 204856
rect 173157 204851 173223 204854
rect 258574 204852 258580 204854
rect 258644 204852 258650 204916
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 78673 200698 78739 200701
rect 259494 200698 259500 200700
rect 78673 200696 259500 200698
rect 78673 200640 78678 200696
rect 78734 200640 259500 200696
rect 78673 200638 259500 200640
rect 78673 200635 78739 200638
rect 259494 200636 259500 200638
rect 259564 200636 259570 200700
rect 68921 198114 68987 198117
rect 254526 198114 254532 198116
rect 68921 198112 254532 198114
rect 68921 198056 68926 198112
rect 68982 198056 254532 198112
rect 68921 198054 254532 198056
rect 68921 198051 68987 198054
rect 254526 198052 254532 198054
rect 254596 198052 254602 198116
rect 148409 197978 148475 197981
rect 336038 197978 336044 197980
rect 148409 197976 336044 197978
rect 148409 197920 148414 197976
rect 148470 197920 336044 197976
rect 148409 197918 336044 197920
rect 148409 197915 148475 197918
rect 336038 197916 336044 197918
rect 336108 197916 336114 197980
rect 123477 195394 123543 195397
rect 266302 195394 266308 195396
rect 123477 195392 266308 195394
rect 123477 195336 123482 195392
rect 123538 195336 266308 195392
rect 123477 195334 266308 195336
rect 123477 195331 123543 195334
rect 266302 195332 266308 195334
rect 266372 195332 266378 195396
rect 65926 195196 65932 195260
rect 65996 195258 66002 195260
rect 271137 195258 271203 195261
rect 65996 195256 271203 195258
rect 65996 195200 271142 195256
rect 271198 195200 271203 195256
rect 65996 195198 271203 195200
rect 65996 195196 66002 195198
rect 271137 195195 271203 195198
rect 240869 192538 240935 192541
rect 403709 192538 403775 192541
rect 240869 192536 403775 192538
rect 240869 192480 240874 192536
rect 240930 192480 403714 192536
rect 403770 192480 403775 192536
rect 240869 192478 403775 192480
rect 240869 192475 240935 192478
rect 403709 192475 403775 192478
rect 580257 192538 580323 192541
rect 583520 192538 584960 192628
rect 580257 192536 584960 192538
rect 580257 192480 580262 192536
rect 580318 192480 584960 192536
rect 580257 192478 584960 192480
rect 580257 192475 580323 192478
rect 583520 192388 584960 192478
rect 128997 191178 129063 191181
rect 258390 191178 258396 191180
rect 128997 191176 258396 191178
rect 128997 191120 129002 191176
rect 129058 191120 258396 191176
rect 128997 191118 258396 191120
rect 128997 191115 129063 191118
rect 258390 191116 258396 191118
rect 258460 191116 258466 191180
rect 129181 191042 129247 191045
rect 259678 191042 259684 191044
rect 129181 191040 259684 191042
rect 129181 190984 129186 191040
rect 129242 190984 259684 191040
rect 129181 190982 259684 190984
rect 129181 190979 129247 190982
rect 259678 190980 259684 190982
rect 259748 190980 259754 191044
rect 66161 189682 66227 189685
rect 262254 189682 262260 189684
rect 66161 189680 262260 189682
rect 66161 189624 66166 189680
rect 66222 189624 262260 189680
rect 66161 189622 262260 189624
rect 66161 189619 66227 189622
rect 262254 189620 262260 189622
rect 262324 189620 262330 189684
rect 292021 189682 292087 189685
rect 502374 189682 502380 189684
rect 292021 189680 502380 189682
rect 292021 189624 292026 189680
rect 292082 189624 502380 189680
rect 292021 189622 502380 189624
rect 292021 189619 292087 189622
rect 502374 189620 502380 189622
rect 502444 189620 502450 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 232589 187098 232655 187101
rect 263726 187098 263732 187100
rect 232589 187096 263732 187098
rect 232589 187040 232594 187096
rect 232650 187040 263732 187096
rect 232589 187038 263732 187040
rect 232589 187035 232655 187038
rect 263726 187036 263732 187038
rect 263796 187036 263802 187100
rect 69013 186962 69079 186965
rect 249190 186962 249196 186964
rect 69013 186960 249196 186962
rect 69013 186904 69018 186960
rect 69074 186904 249196 186960
rect 69013 186902 249196 186904
rect 69013 186899 69079 186902
rect 249190 186900 249196 186902
rect 249260 186900 249266 186964
rect 200614 185540 200620 185604
rect 200684 185602 200690 185604
rect 332685 185602 332751 185605
rect 200684 185600 332751 185602
rect 200684 185544 332690 185600
rect 332746 185544 332751 185600
rect 200684 185542 332751 185544
rect 200684 185540 200690 185542
rect 332685 185539 332751 185542
rect 226977 184378 227043 184381
rect 256734 184378 256740 184380
rect 226977 184376 256740 184378
rect 226977 184320 226982 184376
rect 227038 184320 256740 184376
rect 226977 184318 256740 184320
rect 226977 184315 227043 184318
rect 256734 184316 256740 184318
rect 256804 184316 256810 184380
rect 70894 184180 70900 184244
rect 70964 184242 70970 184244
rect 270585 184242 270651 184245
rect 70964 184240 270651 184242
rect 70964 184184 270590 184240
rect 270646 184184 270651 184240
rect 70964 184182 270651 184184
rect 70964 184180 70970 184182
rect 270585 184179 270651 184182
rect 100661 183698 100727 183701
rect 166206 183698 166212 183700
rect 100661 183696 166212 183698
rect 100661 183640 100666 183696
rect 100722 183640 166212 183696
rect 100661 183638 166212 183640
rect 100661 183635 100727 183638
rect 166206 183636 166212 183638
rect 166276 183636 166282 183700
rect 232497 183018 232563 183021
rect 343725 183018 343791 183021
rect 232497 183016 343791 183018
rect 232497 182960 232502 183016
rect 232558 182960 343730 183016
rect 343786 182960 343791 183016
rect 232497 182958 343791 182960
rect 232497 182955 232563 182958
rect 343725 182955 343791 182958
rect 170397 182882 170463 182885
rect 347037 182882 347103 182885
rect 170397 182880 347103 182882
rect 170397 182824 170402 182880
rect 170458 182824 347042 182880
rect 347098 182824 347103 182880
rect 170397 182822 347103 182824
rect 170397 182819 170463 182822
rect 347037 182819 347103 182822
rect 168966 181460 168972 181524
rect 169036 181522 169042 181524
rect 207657 181522 207723 181525
rect 169036 181520 207723 181522
rect 169036 181464 207662 181520
rect 207718 181464 207723 181520
rect 169036 181462 207723 181464
rect 169036 181460 169042 181462
rect 207657 181459 207723 181462
rect 209221 181522 209287 181525
rect 321318 181522 321324 181524
rect 209221 181520 321324 181522
rect 209221 181464 209226 181520
rect 209282 181464 321324 181520
rect 209221 181462 321324 181464
rect 209221 181459 209287 181462
rect 321318 181460 321324 181462
rect 321388 181460 321394 181524
rect 133229 181386 133295 181389
rect 252502 181386 252508 181388
rect 133229 181384 252508 181386
rect 133229 181328 133234 181384
rect 133290 181328 252508 181384
rect 133229 181326 252508 181328
rect 133229 181323 133295 181326
rect 252502 181324 252508 181326
rect 252572 181324 252578 181388
rect 105721 180842 105787 180845
rect 166390 180842 166396 180844
rect 105721 180840 166396 180842
rect 105721 180784 105726 180840
rect 105782 180784 166396 180840
rect 105721 180782 166396 180784
rect 105721 180779 105787 180782
rect 166390 180780 166396 180782
rect 166460 180780 166466 180844
rect 239397 180298 239463 180301
rect 255446 180298 255452 180300
rect 239397 180296 255452 180298
rect 239397 180240 239402 180296
rect 239458 180240 255452 180296
rect 239397 180238 255452 180240
rect 239397 180235 239463 180238
rect 255446 180236 255452 180238
rect 255516 180236 255522 180300
rect 233877 180162 233943 180165
rect 262438 180162 262444 180164
rect 233877 180160 262444 180162
rect 233877 180104 233882 180160
rect 233938 180104 262444 180160
rect 233877 180102 262444 180104
rect 233877 180099 233943 180102
rect 262438 180100 262444 180102
rect 262508 180100 262514 180164
rect 197118 179964 197124 180028
rect 197188 180026 197194 180028
rect 346577 180026 346643 180029
rect 197188 180024 346643 180026
rect 197188 179968 346582 180024
rect 346638 179968 346643 180024
rect 197188 179966 346643 179968
rect 197188 179964 197194 179966
rect 346577 179963 346643 179966
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 492581 179074 492647 179077
rect 492581 179072 493610 179074
rect 492581 179016 492586 179072
rect 492642 179016 493610 179072
rect 583520 179060 584960 179150
rect 492581 179014 493610 179016
rect 492581 179011 492647 179014
rect 493550 178938 493610 179014
rect 493550 178878 493764 178938
rect 245009 178802 245075 178805
rect 269062 178802 269068 178804
rect 245009 178800 269068 178802
rect 245009 178744 245014 178800
rect 245070 178744 269068 178800
rect 245009 178742 269068 178744
rect 245009 178739 245075 178742
rect 269062 178740 269068 178742
rect 269132 178740 269138 178804
rect 130377 178666 130443 178669
rect 249374 178666 249380 178668
rect 130377 178664 249380 178666
rect 130377 178608 130382 178664
rect 130438 178608 249380 178664
rect 130377 178606 249380 178608
rect 130377 178603 130443 178606
rect 249374 178604 249380 178606
rect 249444 178604 249450 178668
rect 307017 178666 307083 178669
rect 331438 178666 331444 178668
rect 307017 178664 331444 178666
rect 307017 178608 307022 178664
rect 307078 178608 331444 178664
rect 307017 178606 331444 178608
rect 307017 178603 307083 178606
rect 331438 178604 331444 178606
rect 331508 178604 331514 178668
rect 342846 178060 342852 178124
rect 342916 178122 342922 178124
rect 420134 178122 420194 178636
rect 342916 178062 420194 178122
rect 342916 178060 342922 178062
rect 100702 177652 100708 177716
rect 100772 177714 100778 177716
rect 102041 177714 102107 177717
rect 105721 177716 105787 177717
rect 105670 177714 105676 177716
rect 100772 177712 102107 177714
rect 100772 177656 102046 177712
rect 102102 177656 102107 177712
rect 100772 177654 102107 177656
rect 105630 177654 105676 177714
rect 105740 177712 105787 177716
rect 105782 177656 105787 177712
rect 100772 177652 100778 177654
rect 102041 177651 102107 177654
rect 105670 177652 105676 177654
rect 105740 177652 105787 177656
rect 106958 177652 106964 177716
rect 107028 177714 107034 177716
rect 107561 177714 107627 177717
rect 110689 177716 110755 177717
rect 110638 177714 110644 177716
rect 107028 177712 107627 177714
rect 107028 177656 107566 177712
rect 107622 177656 107627 177712
rect 107028 177654 107627 177656
rect 110598 177654 110644 177714
rect 110708 177712 110755 177716
rect 110750 177656 110755 177712
rect 107028 177652 107034 177654
rect 105721 177651 105787 177652
rect 107561 177651 107627 177654
rect 110638 177652 110644 177654
rect 110708 177652 110755 177656
rect 112110 177652 112116 177716
rect 112180 177714 112186 177716
rect 112437 177714 112503 177717
rect 118417 177716 118483 177717
rect 119521 177716 119587 177717
rect 118366 177714 118372 177716
rect 112180 177712 112503 177714
rect 112180 177656 112442 177712
rect 112498 177656 112503 177712
rect 112180 177654 112503 177656
rect 118326 177654 118372 177714
rect 118436 177712 118483 177716
rect 119470 177714 119476 177716
rect 118478 177656 118483 177712
rect 112180 177652 112186 177654
rect 110689 177651 110755 177652
rect 112437 177651 112503 177654
rect 118366 177652 118372 177654
rect 118436 177652 118483 177656
rect 119430 177654 119476 177714
rect 119540 177712 119587 177716
rect 119582 177656 119587 177712
rect 119470 177652 119476 177654
rect 119540 177652 119587 177656
rect 123150 177652 123156 177716
rect 123220 177714 123226 177716
rect 124029 177714 124095 177717
rect 123220 177712 124095 177714
rect 123220 177656 124034 177712
rect 124090 177656 124095 177712
rect 123220 177654 124095 177656
rect 123220 177652 123226 177654
rect 118417 177651 118483 177652
rect 119521 177651 119587 177652
rect 124029 177651 124095 177654
rect 124438 177652 124444 177716
rect 124508 177714 124514 177716
rect 125501 177714 125567 177717
rect 129457 177716 129523 177717
rect 132401 177716 132467 177717
rect 129406 177714 129412 177716
rect 124508 177712 125567 177714
rect 124508 177656 125506 177712
rect 125562 177656 125567 177712
rect 124508 177654 125567 177656
rect 129366 177654 129412 177714
rect 129476 177712 129523 177716
rect 132350 177714 132356 177716
rect 129518 177656 129523 177712
rect 124508 177652 124514 177654
rect 125501 177651 125567 177654
rect 129406 177652 129412 177654
rect 129476 177652 129523 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 129457 177651 129523 177652
rect 132401 177651 132467 177652
rect 319437 177442 319503 177445
rect 338297 177442 338363 177445
rect 319437 177440 338363 177442
rect 319437 177384 319442 177440
rect 319498 177384 338302 177440
rect 338358 177384 338363 177440
rect 319437 177382 338363 177384
rect 319437 177379 319503 177382
rect 338297 177379 338363 177382
rect 162117 177306 162183 177309
rect 204897 177306 204963 177309
rect 162117 177304 204963 177306
rect 162117 177248 162122 177304
rect 162178 177248 204902 177304
rect 204958 177248 204963 177304
rect 162117 177246 204963 177248
rect 162117 177243 162183 177246
rect 204897 177243 204963 177246
rect 316769 177306 316835 177309
rect 336825 177306 336891 177309
rect 494102 177308 494162 177820
rect 316769 177304 336891 177306
rect 316769 177248 316774 177304
rect 316830 177248 336830 177304
rect 336886 177248 336891 177304
rect 316769 177246 336891 177248
rect 316769 177243 316835 177246
rect 336825 177243 336891 177246
rect 494094 177244 494100 177308
rect 494164 177244 494170 177308
rect 97022 176972 97028 177036
rect 97092 177034 97098 177036
rect 97809 177034 97875 177037
rect 115841 177036 115907 177037
rect 115790 177034 115796 177036
rect 97092 177032 97875 177034
rect 97092 176976 97814 177032
rect 97870 176976 97875 177032
rect 97092 176974 97875 176976
rect 115750 176974 115796 177034
rect 115860 177032 115907 177036
rect 115902 176976 115907 177032
rect 97092 176972 97098 176974
rect 97809 176971 97875 176974
rect 115790 176972 115796 176974
rect 115860 176972 115907 176976
rect 125726 176972 125732 177036
rect 125796 177034 125802 177036
rect 126605 177034 126671 177037
rect 125796 177032 126671 177034
rect 125796 176976 126610 177032
rect 126666 176976 126671 177032
rect 125796 176974 126671 176976
rect 125796 176972 125802 176974
rect 115841 176971 115907 176972
rect 126605 176971 126671 176974
rect 134374 176972 134380 177036
rect 134444 177034 134450 177036
rect 134701 177034 134767 177037
rect 134444 177032 134767 177034
rect 134444 176976 134706 177032
rect 134762 176976 134767 177032
rect 134444 176974 134767 176976
rect 134444 176972 134450 176974
rect 134701 176971 134767 176974
rect 416773 177034 416839 177037
rect 416773 177032 420164 177034
rect 416773 176976 416778 177032
rect 416834 176976 420164 177032
rect 416773 176974 420164 176976
rect 416773 176971 416839 176974
rect 114318 176836 114324 176900
rect 114388 176898 114394 176900
rect 214414 176898 214420 176900
rect 114388 176838 214420 176898
rect 114388 176836 114394 176838
rect 214414 176836 214420 176838
rect 214484 176836 214490 176900
rect 98310 176700 98316 176764
rect 98380 176762 98386 176764
rect 98729 176762 98795 176765
rect 100661 176762 100727 176765
rect 103329 176762 103395 176765
rect 104617 176764 104683 176765
rect 108113 176764 108179 176765
rect 104566 176762 104572 176764
rect 98380 176760 98795 176762
rect 98380 176704 98734 176760
rect 98790 176704 98795 176760
rect 98380 176702 98795 176704
rect 98380 176700 98386 176702
rect 98729 176699 98795 176702
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 104526 176702 104572 176762
rect 104636 176760 104683 176764
rect 108062 176762 108068 176764
rect 104678 176704 104683 176760
rect 104566 176700 104572 176702
rect 104636 176700 104683 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 110321 176762 110387 176765
rect 109604 176760 110387 176762
rect 109604 176704 110326 176760
rect 110382 176704 110387 176760
rect 109604 176702 110387 176704
rect 109604 176700 109610 176702
rect 104617 176699 104683 176700
rect 108113 176699 108179 176700
rect 110321 176699 110387 176702
rect 113214 176700 113220 176764
rect 113284 176762 113290 176764
rect 113725 176762 113791 176765
rect 127065 176764 127131 176765
rect 133137 176764 133203 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 127014 176762 127020 176764
rect 113284 176760 113791 176762
rect 113284 176704 113730 176760
rect 113786 176704 113791 176760
rect 113284 176702 113791 176704
rect 126974 176702 127020 176762
rect 127084 176760 127131 176764
rect 133086 176762 133092 176764
rect 127126 176704 127131 176760
rect 113284 176700 113290 176702
rect 113725 176699 113791 176702
rect 127014 176700 127020 176702
rect 127084 176700 127131 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 136030 176762 136036 176764
rect 133198 176704 133203 176760
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 159909 176762 159975 176765
rect 499798 176762 499804 176764
rect 158916 176760 159975 176762
rect 158916 176704 159914 176760
rect 159970 176704 159975 176760
rect 158916 176702 159975 176704
rect 494316 176702 499804 176762
rect 158916 176700 158922 176702
rect 127065 176699 127131 176700
rect 133137 176699 133203 176700
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 159909 176699 159975 176702
rect 499798 176700 499804 176702
rect 499868 176700 499874 176764
rect 103286 176492 103346 176699
rect 128169 176492 128235 176493
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176490 128124 176492
rect 128078 176430 128124 176490
rect 128188 176488 128235 176492
rect 128230 176432 128235 176488
rect 128118 176428 128124 176430
rect 128188 176428 128235 176432
rect 128169 176427 128235 176428
rect 213913 176218 213979 176221
rect 321686 176218 321692 176220
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 217182 175644 217242 176158
rect 315990 176158 321692 176218
rect 235257 175946 235323 175949
rect 256877 175946 256943 175949
rect 235257 175944 256943 175946
rect 235257 175888 235262 175944
rect 235318 175888 256882 175944
rect 256938 175888 256943 175944
rect 235257 175886 256943 175888
rect 235257 175883 235323 175886
rect 256877 175883 256943 175886
rect 266997 175946 267063 175949
rect 315990 175946 316050 176158
rect 321686 176156 321692 176158
rect 321756 176156 321762 176220
rect 266997 175944 316050 175946
rect 266997 175888 267002 175944
rect 267058 175888 316050 175944
rect 266997 175886 316050 175888
rect 266997 175883 267063 175886
rect 247953 175810 248019 175813
rect 247953 175808 248338 175810
rect 247953 175752 247958 175808
rect 248014 175752 248338 175808
rect 247953 175750 248338 175752
rect 247953 175747 248019 175750
rect 248278 175644 248338 175750
rect 320214 175748 320220 175812
rect 320284 175810 320290 175812
rect 321369 175810 321435 175813
rect 320284 175808 321435 175810
rect 320284 175752 321374 175808
rect 321430 175752 321435 175808
rect 320284 175750 321435 175752
rect 320284 175748 320290 175750
rect 321369 175747 321435 175750
rect 307017 175674 307083 175677
rect 313917 175674 313983 175677
rect 498101 175674 498167 175677
rect 307017 175672 310132 175674
rect 307017 175616 307022 175672
rect 307078 175616 310132 175672
rect 307017 175614 310132 175616
rect 313917 175672 321386 175674
rect 313917 175616 313922 175672
rect 313978 175616 321386 175672
rect 313917 175614 321386 175616
rect 494316 175672 498167 175674
rect 494316 175616 498106 175672
rect 498162 175616 498167 175672
rect 494316 175614 498167 175616
rect 307017 175611 307083 175614
rect 313917 175611 313983 175614
rect 321326 175508 321386 175614
rect 498101 175611 498167 175614
rect 102041 175404 102107 175405
rect 116945 175404 117011 175405
rect 120809 175404 120875 175405
rect 121913 175404 121979 175405
rect 130745 175404 130811 175405
rect 101990 175402 101996 175404
rect 101950 175342 101996 175402
rect 102060 175400 102107 175404
rect 116894 175402 116900 175404
rect 102102 175344 102107 175400
rect 101990 175340 101996 175342
rect 102060 175340 102107 175344
rect 116854 175342 116900 175402
rect 116964 175400 117011 175404
rect 120758 175402 120764 175404
rect 117006 175344 117011 175400
rect 116894 175340 116900 175342
rect 116964 175340 117011 175344
rect 120718 175342 120764 175402
rect 120828 175400 120875 175404
rect 121862 175402 121868 175404
rect 120870 175344 120875 175400
rect 120758 175340 120764 175342
rect 120828 175340 120875 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 130694 175402 130700 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 130654 175342 130700 175402
rect 130764 175400 130811 175404
rect 130806 175344 130811 175400
rect 130694 175340 130700 175342
rect 130764 175340 130811 175344
rect 102041 175339 102107 175340
rect 116945 175339 117011 175340
rect 120809 175339 120875 175340
rect 121913 175339 121979 175340
rect 130745 175339 130811 175340
rect 249149 175266 249215 175269
rect 248952 175264 249215 175266
rect 248952 175208 249154 175264
rect 249210 175208 249215 175264
rect 248952 175206 249215 175208
rect 249149 175203 249215 175206
rect 307293 175266 307359 175269
rect 307293 175264 310040 175266
rect 307293 175208 307298 175264
rect 307354 175208 310040 175264
rect 307293 175206 310040 175208
rect 307293 175203 307359 175206
rect 332910 175204 332916 175268
rect 332980 175266 332986 175268
rect 336917 175266 336983 175269
rect 332980 175264 336983 175266
rect 332980 175208 336922 175264
rect 336978 175208 336983 175264
rect 332980 175206 336983 175208
rect 332980 175204 332986 175206
rect 336917 175203 336983 175206
rect 416773 175266 416839 175269
rect 416773 175264 420164 175266
rect 416773 175208 416778 175264
rect 416834 175208 420164 175264
rect 416773 175206 420164 175208
rect 416773 175203 416839 175206
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 217182 174964 217242 175070
rect 307569 174858 307635 174861
rect 307569 174856 310040 174858
rect 307569 174800 307574 174856
rect 307630 174800 310040 174856
rect 307569 174798 310040 174800
rect 307569 174795 307635 174798
rect 214005 174722 214071 174725
rect 249374 174722 249380 174724
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 248952 174662 249380 174722
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 249374 174660 249380 174662
rect 249444 174660 249450 174724
rect 322933 174722 322999 174725
rect 321908 174720 322999 174722
rect 321908 174664 322938 174720
rect 322994 174664 322999 174720
rect 321908 174662 322999 174664
rect 322933 174659 322999 174662
rect 307661 174450 307727 174453
rect 496854 174450 496860 174452
rect 307661 174448 310040 174450
rect 307661 174392 307666 174448
rect 307722 174392 310040 174448
rect 307661 174390 310040 174392
rect 494316 174390 496860 174450
rect 307661 174387 307727 174390
rect 496854 174388 496860 174390
rect 496924 174388 496930 174452
rect 249190 174314 249196 174316
rect 248952 174254 249196 174314
rect 249190 174252 249196 174254
rect 249260 174252 249266 174316
rect 307109 174042 307175 174045
rect 324497 174042 324563 174045
rect 307109 174040 310040 174042
rect 307109 173984 307114 174040
rect 307170 173984 310040 174040
rect 307109 173982 310040 173984
rect 321908 174040 324563 174042
rect 321908 173984 324502 174040
rect 324558 173984 324563 174040
rect 321908 173982 324563 173984
rect 307109 173979 307175 173982
rect 324497 173979 324563 173982
rect 213913 173770 213979 173773
rect 249333 173770 249399 173773
rect 321369 173770 321435 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 248952 173768 249399 173770
rect 248952 173712 249338 173768
rect 249394 173712 249399 173768
rect 248952 173710 249399 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 249333 173707 249399 173710
rect 321326 173768 321435 173770
rect 321326 173712 321374 173768
rect 321430 173712 321435 173768
rect 321326 173707 321435 173712
rect 307569 173634 307635 173637
rect 307569 173632 310040 173634
rect 307569 173576 307574 173632
rect 307630 173576 310040 173632
rect 307569 173574 310040 173576
rect 307569 173571 307635 173574
rect 214097 173362 214163 173365
rect 252461 173362 252527 173365
rect 214097 173360 217242 173362
rect 214097 173304 214102 173360
rect 214158 173304 217242 173360
rect 214097 173302 217242 173304
rect 248952 173360 252527 173362
rect 248952 173304 252466 173360
rect 252522 173304 252527 173360
rect 248952 173302 252527 173304
rect 214097 173299 214163 173302
rect 217182 172924 217242 173302
rect 252461 173299 252527 173302
rect 307109 173226 307175 173229
rect 307109 173224 310040 173226
rect 307109 173168 307114 173224
rect 307170 173168 310040 173224
rect 321326 173196 321386 173707
rect 307109 173166 310040 173168
rect 307109 173163 307175 173166
rect 249241 172818 249307 172821
rect 248952 172816 249307 172818
rect 248952 172760 249246 172816
rect 249302 172760 249307 172816
rect 248952 172758 249307 172760
rect 249241 172755 249307 172758
rect 307661 172682 307727 172685
rect 321277 172682 321343 172685
rect 307661 172680 310040 172682
rect 307661 172624 307666 172680
rect 307722 172624 310040 172680
rect 307661 172622 310040 172624
rect 321277 172680 321386 172682
rect 321277 172624 321282 172680
rect 321338 172624 321386 172680
rect 307661 172619 307727 172622
rect 321277 172619 321386 172624
rect 213913 172410 213979 172413
rect 252461 172410 252527 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 248952 172408 252527 172410
rect 248952 172352 252466 172408
rect 252522 172352 252527 172408
rect 321326 172380 321386 172619
rect 332910 172484 332916 172548
rect 332980 172546 332986 172548
rect 420134 172546 420194 173604
rect 496905 173362 496971 173365
rect 494316 173360 496971 173362
rect 494316 173304 496910 173360
rect 496966 173304 496971 173360
rect 494316 173302 496971 173304
rect 496905 173299 496971 173302
rect 332980 172486 420194 172546
rect 332980 172484 332986 172486
rect 248952 172350 252527 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 252461 172347 252527 172350
rect 306925 172274 306991 172277
rect 306925 172272 310040 172274
rect 306925 172216 306930 172272
rect 306986 172216 310040 172272
rect 306925 172214 310040 172216
rect 306925 172211 306991 172214
rect 214189 172002 214255 172005
rect 214189 172000 217242 172002
rect 214189 171944 214194 172000
rect 214250 171944 217242 172000
rect 214189 171942 217242 171944
rect 214189 171939 214255 171942
rect 167637 171594 167703 171597
rect 164694 171592 167703 171594
rect 164694 171536 167642 171592
rect 167698 171536 167703 171592
rect 217182 171564 217242 171942
rect 252461 171866 252527 171869
rect 248952 171864 252527 171866
rect 248952 171808 252466 171864
rect 252522 171808 252527 171864
rect 248952 171806 252527 171808
rect 252461 171803 252527 171806
rect 307661 171866 307727 171869
rect 307661 171864 310040 171866
rect 307661 171808 307666 171864
rect 307722 171808 310040 171864
rect 307661 171806 310040 171808
rect 307661 171803 307727 171806
rect 324313 171730 324379 171733
rect 321908 171728 324379 171730
rect 321908 171672 324318 171728
rect 324374 171672 324379 171728
rect 321908 171670 324379 171672
rect 324313 171667 324379 171670
rect 164694 171534 167703 171536
rect 167637 171531 167703 171534
rect 252093 171458 252159 171461
rect 248952 171456 252159 171458
rect 248952 171400 252098 171456
rect 252154 171400 252159 171456
rect 248952 171398 252159 171400
rect 252093 171395 252159 171398
rect 306741 171458 306807 171461
rect 306741 171456 310040 171458
rect 306741 171400 306746 171456
rect 306802 171400 310040 171456
rect 306741 171398 310040 171400
rect 306741 171395 306807 171398
rect 216998 171126 217242 171186
rect 216998 171050 217058 171126
rect 215250 170990 217058 171050
rect 217182 171020 217242 171126
rect 334750 171124 334756 171188
rect 334820 171186 334826 171188
rect 420134 171186 420194 171836
rect 494286 171733 494346 172244
rect 494237 171728 494346 171733
rect 494237 171672 494242 171728
rect 494298 171672 494346 171728
rect 494237 171670 494346 171672
rect 494237 171667 494303 171670
rect 494462 171458 494468 171460
rect 334820 171126 420194 171186
rect 494286 171398 494468 171458
rect 494286 171156 494346 171398
rect 494462 171396 494468 171398
rect 494532 171396 494538 171460
rect 334820 171124 334826 171126
rect 307293 171050 307359 171053
rect 307293 171048 310040 171050
rect 307293 170992 307298 171048
rect 307354 170992 310040 171048
rect 307293 170990 310040 170992
rect 214557 170914 214623 170917
rect 215250 170914 215310 170990
rect 307293 170987 307359 170990
rect 256734 170914 256740 170916
rect 214557 170912 215310 170914
rect 214557 170856 214562 170912
rect 214618 170856 215310 170912
rect 214557 170854 215310 170856
rect 248952 170854 256740 170914
rect 214557 170851 214623 170854
rect 256734 170852 256740 170854
rect 256804 170852 256810 170916
rect 324313 170914 324379 170917
rect 321908 170912 324379 170914
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 324313 170851 324379 170854
rect 213913 170778 213979 170781
rect 213913 170776 217242 170778
rect 213913 170720 213918 170776
rect 213974 170720 217242 170776
rect 213913 170718 217242 170720
rect 213913 170715 213979 170718
rect 217182 170340 217242 170718
rect 307661 170642 307727 170645
rect 307661 170640 310040 170642
rect 307661 170584 307666 170640
rect 307722 170584 310040 170640
rect 307661 170582 310040 170584
rect 307661 170579 307727 170582
rect 321318 170580 321324 170644
rect 321388 170580 321394 170644
rect 252461 170506 252527 170509
rect 248952 170504 252527 170506
rect 248952 170448 252466 170504
rect 252522 170448 252527 170504
rect 248952 170446 252527 170448
rect 252461 170443 252527 170446
rect 306557 170234 306623 170237
rect 306557 170232 310040 170234
rect 306557 170176 306562 170232
rect 306618 170176 310040 170232
rect 306557 170174 310040 170176
rect 306557 170171 306623 170174
rect 252369 170098 252435 170101
rect 248952 170096 252435 170098
rect 248952 170040 252374 170096
rect 252430 170040 252435 170096
rect 321326 170068 321386 170580
rect 248952 170038 252435 170040
rect 252369 170035 252435 170038
rect 307477 169826 307543 169829
rect 216998 169766 217242 169826
rect 214649 169690 214715 169693
rect 216998 169690 217058 169766
rect 214649 169688 217058 169690
rect 214649 169632 214654 169688
rect 214710 169632 217058 169688
rect 217182 169660 217242 169766
rect 307477 169824 310040 169826
rect 307477 169768 307482 169824
rect 307538 169768 310040 169824
rect 307477 169766 310040 169768
rect 307477 169763 307543 169766
rect 335854 169764 335860 169828
rect 335924 169826 335930 169828
rect 420134 169826 420194 170204
rect 495525 169962 495591 169965
rect 494316 169960 495591 169962
rect 494316 169904 495530 169960
rect 495586 169904 495591 169960
rect 494316 169902 495591 169904
rect 495525 169899 495591 169902
rect 335924 169766 420194 169826
rect 335924 169764 335930 169766
rect 214649 169630 217058 169632
rect 214649 169627 214715 169630
rect 249977 169554 250043 169557
rect 248952 169552 250043 169554
rect 248952 169496 249982 169552
rect 250038 169496 250043 169552
rect 248952 169494 250043 169496
rect 249977 169491 250043 169494
rect 213913 169418 213979 169421
rect 324313 169418 324379 169421
rect 213913 169416 217242 169418
rect 213913 169360 213918 169416
rect 213974 169360 217242 169416
rect 213913 169358 217242 169360
rect 321908 169416 324379 169418
rect 321908 169360 324318 169416
rect 324374 169360 324379 169416
rect 321908 169358 324379 169360
rect 213913 169355 213979 169358
rect 217182 168980 217242 169358
rect 324313 169355 324379 169358
rect 307109 169282 307175 169285
rect 307109 169280 310040 169282
rect 307109 169224 307114 169280
rect 307170 169224 310040 169280
rect 307109 169222 310040 169224
rect 307109 169219 307175 169222
rect 252461 169146 252527 169149
rect 248952 169144 252527 169146
rect 248952 169088 252466 169144
rect 252522 169088 252527 169144
rect 248952 169086 252527 169088
rect 252461 169083 252527 169086
rect 307661 168874 307727 168877
rect 495617 168874 495683 168877
rect 307661 168872 310040 168874
rect 307661 168816 307666 168872
rect 307722 168816 310040 168872
rect 307661 168814 310040 168816
rect 494316 168872 495683 168874
rect 494316 168816 495622 168872
rect 495678 168816 495683 168872
rect 494316 168814 495683 168816
rect 307661 168811 307727 168814
rect 495617 168811 495683 168814
rect 252369 168602 252435 168605
rect 324497 168602 324563 168605
rect 248952 168600 252435 168602
rect 248952 168544 252374 168600
rect 252430 168544 252435 168600
rect 248952 168542 252435 168544
rect 321908 168600 324563 168602
rect 321908 168544 324502 168600
rect 324558 168544 324563 168600
rect 321908 168542 324563 168544
rect 252369 168539 252435 168542
rect 324497 168539 324563 168542
rect 306557 168466 306623 168469
rect 416773 168466 416839 168469
rect 216998 168406 217242 168466
rect 213913 168330 213979 168333
rect 216998 168330 217058 168406
rect 213913 168328 217058 168330
rect 213913 168272 213918 168328
rect 213974 168272 217058 168328
rect 217182 168300 217242 168406
rect 306557 168464 310040 168466
rect 306557 168408 306562 168464
rect 306618 168408 310040 168464
rect 306557 168406 310040 168408
rect 416773 168464 420164 168466
rect 416773 168408 416778 168464
rect 416834 168408 420164 168464
rect 416773 168406 420164 168408
rect 306557 168403 306623 168406
rect 416773 168403 416839 168406
rect 213913 168270 217058 168272
rect 213913 168267 213979 168270
rect 252461 168194 252527 168197
rect 248952 168192 252527 168194
rect 248952 168136 252466 168192
rect 252522 168136 252527 168192
rect 248952 168134 252527 168136
rect 252461 168131 252527 168134
rect 214005 168058 214071 168061
rect 307477 168058 307543 168061
rect 214005 168056 217242 168058
rect 214005 168000 214010 168056
rect 214066 168000 217242 168056
rect 214005 167998 217242 168000
rect 214005 167995 214071 167998
rect 217182 167620 217242 167998
rect 307477 168056 310040 168058
rect 307477 168000 307482 168056
rect 307538 168000 310040 168056
rect 307477 167998 310040 168000
rect 307477 167995 307543 167998
rect 324313 167786 324379 167789
rect 496905 167786 496971 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 494316 167784 496971 167786
rect 494316 167728 496910 167784
rect 496966 167728 496971 167784
rect 494316 167726 496971 167728
rect 324313 167723 324379 167726
rect 496905 167723 496971 167726
rect 252461 167650 252527 167653
rect 248952 167648 252527 167650
rect 248952 167592 252466 167648
rect 252522 167592 252527 167648
rect 248952 167590 252527 167592
rect 252461 167587 252527 167590
rect 307385 167650 307451 167653
rect 307385 167648 310040 167650
rect 307385 167592 307390 167648
rect 307446 167592 310040 167648
rect 307385 167590 310040 167592
rect 307385 167587 307451 167590
rect 252737 167242 252803 167245
rect 248952 167240 252803 167242
rect 248952 167184 252742 167240
rect 252798 167184 252803 167240
rect 248952 167182 252803 167184
rect 252737 167179 252803 167182
rect 307293 167242 307359 167245
rect 307293 167240 310040 167242
rect 307293 167184 307298 167240
rect 307354 167184 310040 167240
rect 307293 167182 310040 167184
rect 307293 167179 307359 167182
rect 324497 167106 324563 167109
rect 321908 167104 324563 167106
rect 321908 167048 324502 167104
rect 324558 167048 324563 167104
rect 321908 167046 324563 167048
rect 324497 167043 324563 167046
rect 213913 166970 213979 166973
rect 216998 166970 217242 167010
rect 213913 166968 217242 166970
rect 213913 166912 213918 166968
rect 213974 166950 217242 166968
rect 213974 166912 217058 166950
rect 217182 166940 217242 166950
rect 213913 166910 217058 166912
rect 213913 166907 213979 166910
rect 307661 166834 307727 166837
rect 416773 166834 416839 166837
rect 307661 166832 310040 166834
rect 307661 166776 307666 166832
rect 307722 166776 310040 166832
rect 307661 166774 310040 166776
rect 416773 166832 420164 166834
rect 416773 166776 416778 166832
rect 416834 166776 420164 166832
rect 416773 166774 420164 166776
rect 307661 166771 307727 166774
rect 416773 166771 416839 166774
rect 214005 166698 214071 166701
rect 252461 166698 252527 166701
rect 496905 166698 496971 166701
rect 214005 166696 217242 166698
rect 214005 166640 214010 166696
rect 214066 166640 217242 166696
rect 214005 166638 217242 166640
rect 248952 166696 252527 166698
rect 248952 166640 252466 166696
rect 252522 166640 252527 166696
rect 248952 166638 252527 166640
rect 494316 166696 496971 166698
rect 494316 166640 496910 166696
rect 496966 166640 496971 166696
rect 494316 166638 496971 166640
rect 214005 166635 214071 166638
rect 217182 166396 217242 166638
rect 252461 166635 252527 166638
rect 496905 166635 496971 166638
rect 307477 166426 307543 166429
rect 307477 166424 310040 166426
rect 307477 166368 307482 166424
rect 307538 166368 310040 166424
rect 307477 166366 310040 166368
rect 307477 166363 307543 166366
rect 252369 166290 252435 166293
rect 324313 166290 324379 166293
rect 248952 166288 252435 166290
rect 248952 166232 252374 166288
rect 252430 166232 252435 166288
rect 248952 166230 252435 166232
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 252369 166227 252435 166230
rect 324313 166227 324379 166230
rect 214097 166154 214163 166157
rect 214097 166152 217242 166154
rect 214097 166096 214102 166152
rect 214158 166096 217242 166152
rect 214097 166094 217242 166096
rect 214097 166091 214163 166094
rect 217182 165716 217242 166094
rect 306741 165882 306807 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 306741 165880 310040 165882
rect 306741 165824 306746 165880
rect 306802 165824 310040 165880
rect 306741 165822 310040 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 306741 165819 306807 165822
rect 580165 165819 580231 165822
rect 252277 165746 252343 165749
rect 248952 165744 252343 165746
rect 248952 165688 252282 165744
rect 252338 165688 252343 165744
rect 583520 165732 584960 165822
rect 248952 165686 252343 165688
rect 252277 165683 252343 165686
rect 307201 165474 307267 165477
rect 324313 165474 324379 165477
rect 496905 165474 496971 165477
rect 307201 165472 310040 165474
rect 307201 165416 307206 165472
rect 307262 165416 310040 165472
rect 307201 165414 310040 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 494316 165472 496971 165474
rect 494316 165416 496910 165472
rect 496966 165416 496971 165472
rect 494316 165414 496971 165416
rect 307201 165411 307267 165414
rect 324313 165411 324379 165414
rect 496905 165411 496971 165414
rect 213913 165338 213979 165341
rect 252461 165338 252527 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 248952 165336 252527 165338
rect 248952 165280 252466 165336
rect 252522 165280 252527 165336
rect 248952 165278 252527 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 252461 165275 252527 165278
rect 307017 165066 307083 165069
rect 416773 165066 416839 165069
rect 307017 165064 310040 165066
rect 307017 165008 307022 165064
rect 307078 165008 310040 165064
rect 307017 165006 310040 165008
rect 416773 165064 420164 165066
rect 416773 165008 416778 165064
rect 416834 165008 420164 165064
rect 416773 165006 420164 165008
rect 307017 165003 307083 165006
rect 416773 165003 416839 165006
rect 214414 164732 214420 164796
rect 214484 164794 214490 164796
rect 252369 164794 252435 164797
rect 324497 164794 324563 164797
rect 214484 164734 217242 164794
rect 248952 164792 252435 164794
rect 248952 164736 252374 164792
rect 252430 164736 252435 164792
rect 248952 164734 252435 164736
rect 321908 164792 324563 164794
rect 321908 164736 324502 164792
rect 324558 164736 324563 164792
rect 321908 164734 324563 164736
rect 214484 164732 214490 164734
rect 217182 164356 217242 164734
rect 252369 164731 252435 164734
rect 324497 164731 324563 164734
rect 307661 164658 307727 164661
rect 307661 164656 310040 164658
rect 307661 164600 307666 164656
rect 307722 164600 310040 164656
rect 307661 164598 310040 164600
rect 307661 164595 307727 164598
rect 252277 164386 252343 164389
rect 496997 164386 497063 164389
rect 248952 164384 252343 164386
rect 248952 164328 252282 164384
rect 252338 164328 252343 164384
rect 248952 164326 252343 164328
rect 494316 164384 497063 164386
rect 494316 164328 497002 164384
rect 497058 164328 497063 164384
rect 494316 164326 497063 164328
rect 252277 164323 252343 164326
rect 496997 164323 497063 164326
rect 307109 164250 307175 164253
rect 307109 164248 310040 164250
rect 307109 164192 307114 164248
rect 307170 164192 310040 164248
rect 307109 164190 310040 164192
rect 307109 164187 307175 164190
rect 213913 164114 213979 164117
rect 213913 164112 217242 164114
rect 213913 164056 213918 164112
rect 213974 164056 217242 164112
rect 213913 164054 217242 164056
rect 213913 164051 213979 164054
rect 217182 163676 217242 164054
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 248952 163976 252527 163978
rect 248952 163920 252466 163976
rect 252522 163920 252527 163976
rect 248952 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 307569 163842 307635 163845
rect 307569 163840 310040 163842
rect 307569 163784 307574 163840
rect 307630 163784 310040 163840
rect 307569 163782 310040 163784
rect 307569 163779 307635 163782
rect 214005 163434 214071 163437
rect 306741 163434 306807 163437
rect 214005 163432 217242 163434
rect 214005 163376 214010 163432
rect 214066 163376 217242 163432
rect 306741 163432 310040 163434
rect 214005 163374 217242 163376
rect 214005 163371 214071 163374
rect 217182 162996 217242 163374
rect 248860 163330 249442 163390
rect 306741 163376 306746 163432
rect 306802 163376 310040 163432
rect 306741 163374 310040 163376
rect 306741 163371 306807 163374
rect 249382 163162 249442 163330
rect 263726 163162 263732 163164
rect 249382 163102 263732 163162
rect 263726 163100 263732 163102
rect 263796 163100 263802 163164
rect 323117 163162 323183 163165
rect 321908 163160 323183 163162
rect 321908 163104 323122 163160
rect 323178 163104 323183 163160
rect 321908 163102 323183 163104
rect 323117 163099 323183 163102
rect 252369 163026 252435 163029
rect 248952 163024 252435 163026
rect -960 162890 480 162980
rect 248952 162968 252374 163024
rect 252430 162968 252435 163024
rect 248952 162966 252435 162968
rect 252369 162963 252435 162966
rect 307661 163026 307727 163029
rect 307661 163024 310040 163026
rect 307661 162968 307666 163024
rect 307722 162968 310040 163024
rect 307661 162966 310040 162968
rect 307661 162963 307727 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 305637 162890 305703 162893
rect 307569 162890 307635 162893
rect 305637 162888 307635 162890
rect 305637 162832 305642 162888
rect 305698 162832 307574 162888
rect 307630 162832 307635 162888
rect 305637 162830 307635 162832
rect 305637 162827 305703 162830
rect 307569 162827 307635 162830
rect 340270 162828 340276 162892
rect 340340 162890 340346 162892
rect 420134 162890 420194 163404
rect 496905 163298 496971 163301
rect 494316 163296 496971 163298
rect 494316 163240 496910 163296
rect 496966 163240 496971 163296
rect 494316 163238 496971 163240
rect 496905 163235 496971 163238
rect 340340 162830 420194 162890
rect 340340 162828 340346 162830
rect 213913 162618 213979 162621
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 252461 162482 252527 162485
rect 248952 162480 252527 162482
rect 248952 162424 252466 162480
rect 252522 162424 252527 162480
rect 248952 162422 252527 162424
rect 252461 162419 252527 162422
rect 307477 162482 307543 162485
rect 324313 162482 324379 162485
rect 307477 162480 310040 162482
rect 307477 162424 307482 162480
rect 307538 162424 310040 162480
rect 307477 162422 310040 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307477 162419 307543 162422
rect 324313 162419 324379 162422
rect 321737 162210 321803 162213
rect 496905 162210 496971 162213
rect 321694 162208 321803 162210
rect 321694 162152 321742 162208
rect 321798 162152 321803 162208
rect 321694 162147 321803 162152
rect 494316 162208 496971 162210
rect 494316 162152 496910 162208
rect 496966 162152 496971 162208
rect 494316 162150 496971 162152
rect 496905 162147 496971 162150
rect 214005 162074 214071 162077
rect 252369 162074 252435 162077
rect 214005 162072 217242 162074
rect 214005 162016 214010 162072
rect 214066 162016 217242 162072
rect 214005 162014 217242 162016
rect 248952 162072 252435 162074
rect 248952 162016 252374 162072
rect 252430 162016 252435 162072
rect 248952 162014 252435 162016
rect 214005 162011 214071 162014
rect 217182 161772 217242 162014
rect 252369 162011 252435 162014
rect 307569 162074 307635 162077
rect 307569 162072 310040 162074
rect 307569 162016 307574 162072
rect 307630 162016 310040 162072
rect 307569 162014 310040 162016
rect 307569 162011 307635 162014
rect 307661 161666 307727 161669
rect 307661 161664 310040 161666
rect 307661 161608 307666 161664
rect 307722 161608 310040 161664
rect 321694 161636 321754 162147
rect 416773 161802 416839 161805
rect 416773 161800 420164 161802
rect 416773 161744 416778 161800
rect 416834 161744 420164 161800
rect 416773 161742 420164 161744
rect 416773 161739 416839 161742
rect 307661 161606 310040 161608
rect 307661 161603 307727 161606
rect 252829 161530 252895 161533
rect 248952 161528 252895 161530
rect 248952 161472 252834 161528
rect 252890 161472 252895 161528
rect 248952 161470 252895 161472
rect 252829 161467 252895 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 307477 161258 307543 161261
rect 307477 161256 310040 161258
rect 307477 161200 307482 161256
rect 307538 161200 310040 161256
rect 307477 161198 310040 161200
rect 307477 161195 307543 161198
rect 248860 161018 249442 161078
rect 249382 160986 249442 161018
rect 258390 160986 258396 160988
rect 249382 160926 258396 160986
rect 258390 160924 258396 160926
rect 258460 160924 258466 160988
rect 496905 160986 496971 160989
rect 494316 160984 496971 160986
rect 494316 160928 496910 160984
rect 496966 160928 496971 160984
rect 494316 160926 496971 160928
rect 496905 160923 496971 160926
rect 214005 160850 214071 160853
rect 307569 160850 307635 160853
rect 323025 160850 323091 160853
rect 214005 160848 217242 160850
rect 214005 160792 214010 160848
rect 214066 160792 217242 160848
rect 214005 160790 217242 160792
rect 214005 160787 214071 160790
rect 217182 160412 217242 160790
rect 307569 160848 310040 160850
rect 307569 160792 307574 160848
rect 307630 160792 310040 160848
rect 307569 160790 310040 160792
rect 321908 160848 323091 160850
rect 321908 160792 323030 160848
rect 323086 160792 323091 160848
rect 321908 160790 323091 160792
rect 307569 160787 307635 160790
rect 323025 160787 323091 160790
rect 252461 160578 252527 160581
rect 248952 160576 252527 160578
rect 248952 160520 252466 160576
rect 252522 160520 252527 160576
rect 248952 160518 252527 160520
rect 252461 160515 252527 160518
rect 307661 160442 307727 160445
rect 307661 160440 310040 160442
rect 307661 160384 307666 160440
rect 307722 160384 310040 160440
rect 307661 160382 310040 160384
rect 307661 160379 307727 160382
rect 251449 160170 251515 160173
rect 324313 160170 324379 160173
rect 248952 160168 251515 160170
rect 248952 160112 251454 160168
rect 251510 160112 251515 160168
rect 248952 160110 251515 160112
rect 321908 160168 324379 160170
rect 321908 160112 324318 160168
rect 324374 160112 324379 160168
rect 321908 160110 324379 160112
rect 251449 160107 251515 160110
rect 324313 160107 324379 160110
rect 306557 160034 306623 160037
rect 306557 160032 310040 160034
rect 306557 159976 306562 160032
rect 306618 159976 310040 160032
rect 306557 159974 310040 159976
rect 306557 159971 306623 159974
rect 217182 159218 217242 159732
rect 251173 159626 251239 159629
rect 248952 159624 251239 159626
rect 248952 159568 251178 159624
rect 251234 159568 251239 159624
rect 248952 159566 251239 159568
rect 251173 159563 251239 159566
rect 307569 159626 307635 159629
rect 307569 159624 310040 159626
rect 307569 159568 307574 159624
rect 307630 159568 310040 159624
rect 307569 159566 310040 159568
rect 307569 159563 307635 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 251357 159218 251423 159221
rect 200070 159158 217242 159218
rect 248952 159216 251423 159218
rect 248952 159160 251362 159216
rect 251418 159160 251423 159216
rect 248952 159158 251423 159160
rect 166390 158748 166396 158812
rect 166460 158810 166466 158812
rect 200070 158810 200130 159158
rect 251357 159155 251423 159158
rect 307661 159082 307727 159085
rect 307661 159080 310040 159082
rect 166460 158750 200130 158810
rect 214465 158810 214531 158813
rect 217366 158810 217426 159052
rect 307661 159024 307666 159080
rect 307722 159024 310040 159080
rect 307661 159022 310040 159024
rect 307661 159019 307727 159022
rect 251265 158810 251331 158813
rect 214465 158808 217426 158810
rect 214465 158752 214470 158808
rect 214526 158752 217426 158808
rect 214465 158750 217426 158752
rect 248952 158808 251331 158810
rect 248952 158752 251270 158808
rect 251326 158752 251331 158808
rect 248952 158750 251331 158752
rect 166460 158748 166466 158750
rect 214465 158747 214531 158750
rect 251265 158747 251331 158750
rect 338614 158748 338620 158812
rect 338684 158810 338690 158812
rect 420134 158810 420194 160004
rect 496905 159898 496971 159901
rect 494316 159896 496971 159898
rect 494316 159840 496910 159896
rect 496966 159840 496971 159896
rect 494316 159838 496971 159840
rect 496905 159835 496971 159838
rect 496997 158810 497063 158813
rect 338684 158750 420194 158810
rect 494316 158808 497063 158810
rect 494316 158752 497002 158808
rect 497058 158752 497063 158808
rect 494316 158750 497063 158752
rect 338684 158748 338690 158750
rect 496997 158747 497063 158750
rect 214005 158674 214071 158677
rect 306557 158674 306623 158677
rect 322197 158674 322263 158677
rect 214005 158672 217242 158674
rect 214005 158616 214010 158672
rect 214066 158616 217242 158672
rect 214005 158614 217242 158616
rect 214005 158611 214071 158614
rect 217182 158372 217242 158614
rect 306557 158672 310040 158674
rect 306557 158616 306562 158672
rect 306618 158616 310040 158672
rect 306557 158614 310040 158616
rect 321878 158672 322263 158674
rect 321878 158616 322202 158672
rect 322258 158616 322263 158672
rect 321878 158614 322263 158616
rect 306557 158611 306623 158614
rect 321878 158508 321938 158614
rect 322197 158611 322263 158614
rect 416773 158402 416839 158405
rect 416773 158400 420164 158402
rect 416773 158344 416778 158400
rect 416834 158344 420164 158400
rect 416773 158342 420164 158344
rect 416773 158339 416839 158342
rect 252185 158266 252251 158269
rect 248952 158264 252251 158266
rect 248952 158208 252190 158264
rect 252246 158208 252251 158264
rect 248952 158206 252251 158208
rect 252185 158203 252251 158206
rect 307661 158266 307727 158269
rect 307661 158264 310040 158266
rect 307661 158208 307666 158264
rect 307722 158208 310040 158264
rect 307661 158206 310040 158208
rect 307661 158203 307727 158206
rect 213913 158130 213979 158133
rect 213913 158128 217242 158130
rect 213913 158072 213918 158128
rect 213974 158072 217242 158128
rect 213913 158070 217242 158072
rect 213913 158067 213979 158070
rect 217182 157692 217242 158070
rect 251357 157858 251423 157861
rect 248952 157856 251423 157858
rect 248952 157800 251362 157856
rect 251418 157800 251423 157856
rect 248952 157798 251423 157800
rect 251357 157795 251423 157798
rect 307477 157858 307543 157861
rect 324313 157858 324379 157861
rect 307477 157856 310040 157858
rect 307477 157800 307482 157856
rect 307538 157800 310040 157856
rect 307477 157798 310040 157800
rect 321908 157856 324379 157858
rect 321908 157800 324318 157856
rect 324374 157800 324379 157856
rect 321908 157798 324379 157800
rect 307477 157795 307543 157798
rect 324313 157795 324379 157798
rect 496905 157722 496971 157725
rect 494316 157720 496971 157722
rect 494316 157664 496910 157720
rect 496966 157664 496971 157720
rect 494316 157662 496971 157664
rect 496905 157659 496971 157662
rect 307385 157450 307451 157453
rect 307385 157448 310040 157450
rect 307385 157392 307390 157448
rect 307446 157392 310040 157448
rect 307385 157390 310040 157392
rect 307385 157387 307451 157390
rect 213913 157314 213979 157317
rect 252461 157314 252527 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 248952 157312 252527 157314
rect 248952 157256 252466 157312
rect 252522 157256 252527 157312
rect 248952 157254 252527 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 252461 157251 252527 157254
rect 307661 157042 307727 157045
rect 324313 157042 324379 157045
rect 307661 157040 310040 157042
rect 307661 156984 307666 157040
rect 307722 156984 310040 157040
rect 307661 156982 310040 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 307661 156979 307727 156982
rect 324313 156979 324379 156982
rect 252369 156906 252435 156909
rect 248952 156904 252435 156906
rect 248952 156848 252374 156904
rect 252430 156848 252435 156904
rect 248952 156846 252435 156848
rect 252369 156843 252435 156846
rect 307569 156634 307635 156637
rect 416773 156634 416839 156637
rect 307569 156632 310040 156634
rect 307569 156576 307574 156632
rect 307630 156576 310040 156632
rect 307569 156574 310040 156576
rect 416773 156632 420164 156634
rect 416773 156576 416778 156632
rect 416834 156576 420164 156632
rect 416773 156574 420164 156576
rect 307569 156571 307635 156574
rect 416773 156571 416839 156574
rect 496905 156498 496971 156501
rect 494316 156496 496971 156498
rect 166206 156028 166212 156092
rect 166276 156090 166282 156092
rect 217182 156090 217242 156468
rect 494316 156440 496910 156496
rect 496966 156440 496971 156496
rect 494316 156438 496971 156440
rect 496905 156435 496971 156438
rect 255262 156362 255268 156364
rect 248952 156302 255268 156362
rect 255262 156300 255268 156302
rect 255332 156300 255338 156364
rect 324405 156362 324471 156365
rect 321908 156360 324471 156362
rect 321908 156304 324410 156360
rect 324466 156304 324471 156360
rect 321908 156302 324471 156304
rect 324405 156299 324471 156302
rect 306557 156226 306623 156229
rect 306557 156224 310040 156226
rect 306557 156168 306562 156224
rect 306618 156168 310040 156224
rect 306557 156166 310040 156168
rect 306557 156163 306623 156166
rect 166276 156030 217242 156090
rect 166276 156028 166282 156030
rect 213913 155954 213979 155957
rect 252553 155954 252619 155957
rect 213913 155952 217242 155954
rect 213913 155896 213918 155952
rect 213974 155896 217242 155952
rect 213913 155894 217242 155896
rect 248952 155952 252619 155954
rect 248952 155896 252558 155952
rect 252614 155896 252619 155952
rect 248952 155894 252619 155896
rect 213913 155891 213979 155894
rect 217182 155788 217242 155894
rect 252553 155891 252619 155894
rect 307569 155682 307635 155685
rect 307569 155680 310040 155682
rect 307569 155624 307574 155680
rect 307630 155624 310040 155680
rect 307569 155622 310040 155624
rect 307569 155619 307635 155622
rect 214005 155546 214071 155549
rect 324313 155546 324379 155549
rect 214005 155544 217242 155546
rect 214005 155488 214010 155544
rect 214066 155488 217242 155544
rect 214005 155486 217242 155488
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 214005 155483 214071 155486
rect 217182 155108 217242 155486
rect 324313 155483 324379 155486
rect 250253 155410 250319 155413
rect 496905 155410 496971 155413
rect 248952 155408 250319 155410
rect 248952 155352 250258 155408
rect 250314 155352 250319 155408
rect 248952 155350 250319 155352
rect 494316 155408 496971 155410
rect 494316 155352 496910 155408
rect 496966 155352 496971 155408
rect 494316 155350 496971 155352
rect 250253 155347 250319 155350
rect 496905 155347 496971 155350
rect 307477 155274 307543 155277
rect 307477 155272 310040 155274
rect 307477 155216 307482 155272
rect 307538 155216 310040 155272
rect 307477 155214 310040 155216
rect 307477 155211 307543 155214
rect 321686 155212 321692 155276
rect 321756 155212 321762 155276
rect 248860 154898 249442 154958
rect 249382 154594 249442 154898
rect 307661 154866 307727 154869
rect 307661 154864 310040 154866
rect 307661 154808 307666 154864
rect 307722 154808 310040 154864
rect 307661 154806 310040 154808
rect 307661 154803 307727 154806
rect 321694 154700 321754 155212
rect 416773 155002 416839 155005
rect 416773 155000 420164 155002
rect 416773 154944 416778 155000
rect 416834 154944 420164 155000
rect 416773 154942 420164 154944
rect 416773 154939 416839 154942
rect 262438 154594 262444 154596
rect 249382 154534 262444 154594
rect 262438 154532 262444 154534
rect 262508 154532 262514 154596
rect 252461 154458 252527 154461
rect 248952 154456 252527 154458
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 248952 154400 252466 154456
rect 252522 154400 252527 154456
rect 248952 154398 252527 154400
rect 252461 154395 252527 154398
rect 306557 154458 306623 154461
rect 306557 154456 310040 154458
rect 306557 154400 306562 154456
rect 306618 154400 310040 154456
rect 306557 154398 310040 154400
rect 306557 154395 306623 154398
rect 496997 154322 497063 154325
rect 494316 154320 497063 154322
rect 494316 154264 497002 154320
rect 497058 154264 497063 154320
rect 494316 154262 497063 154264
rect 496997 154259 497063 154262
rect 252369 154050 252435 154053
rect 248952 154048 252435 154050
rect 248952 153992 252374 154048
rect 252430 153992 252435 154048
rect 248952 153990 252435 153992
rect 252369 153987 252435 153990
rect 307661 154050 307727 154053
rect 324313 154050 324379 154053
rect 307661 154048 310040 154050
rect 307661 153992 307666 154048
rect 307722 153992 310040 154048
rect 307661 153990 310040 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307661 153987 307727 153990
rect 324313 153987 324379 153990
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 214005 153851 214071 153854
rect 213913 153506 213979 153509
rect 217182 153506 217242 153748
rect 306649 153642 306715 153645
rect 306649 153640 310040 153642
rect 306649 153584 306654 153640
rect 306710 153584 310040 153640
rect 306649 153582 310040 153584
rect 306649 153579 306715 153582
rect 251541 153506 251607 153509
rect 213913 153504 217242 153506
rect 213913 153448 213918 153504
rect 213974 153448 217242 153504
rect 213913 153446 217242 153448
rect 248952 153504 251607 153506
rect 248952 153448 251546 153504
rect 251602 153448 251607 153504
rect 248952 153446 251607 153448
rect 213913 153443 213979 153446
rect 251541 153443 251607 153446
rect 307661 153234 307727 153237
rect 324405 153234 324471 153237
rect 307661 153232 310040 153234
rect 307661 153176 307666 153232
rect 307722 153176 310040 153232
rect 307661 153174 310040 153176
rect 321908 153232 324471 153234
rect 321908 153176 324410 153232
rect 324466 153176 324471 153232
rect 321908 153174 324471 153176
rect 307661 153171 307727 153174
rect 324405 153171 324471 153174
rect 416773 153234 416839 153237
rect 496905 153234 496971 153237
rect 416773 153232 420164 153234
rect 416773 153176 416778 153232
rect 416834 153176 420164 153232
rect 416773 153174 420164 153176
rect 494316 153232 496971 153234
rect 494316 153176 496910 153232
rect 496966 153176 496971 153232
rect 494316 153174 496971 153176
rect 416773 153171 416839 153174
rect 496905 153171 496971 153174
rect 252369 153098 252435 153101
rect 248952 153096 252435 153098
rect 213361 152690 213427 152693
rect 217182 152690 217242 153068
rect 248952 153040 252374 153096
rect 252430 153040 252435 153096
rect 248952 153038 252435 153040
rect 252369 153035 252435 153038
rect 252461 152690 252527 152693
rect 213361 152688 217242 152690
rect 213361 152632 213366 152688
rect 213422 152632 217242 152688
rect 213361 152630 217242 152632
rect 248952 152688 252527 152690
rect 248952 152632 252466 152688
rect 252522 152632 252527 152688
rect 248952 152630 252527 152632
rect 213361 152627 213427 152630
rect 252461 152627 252527 152630
rect 308489 152690 308555 152693
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 308489 152688 310040 152690
rect 308489 152632 308494 152688
rect 308550 152632 310040 152688
rect 308489 152630 310040 152632
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 308489 152627 308555 152630
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 307109 152282 307175 152285
rect 307109 152280 310040 152282
rect 307109 152224 307114 152280
rect 307170 152224 310040 152280
rect 307109 152222 310040 152224
rect 307109 152219 307175 152222
rect 252277 152146 252343 152149
rect 496905 152146 496971 152149
rect 248952 152144 252343 152146
rect 248952 152088 252282 152144
rect 252338 152088 252343 152144
rect 248952 152086 252343 152088
rect 494316 152144 496971 152146
rect 494316 152088 496910 152144
rect 496966 152088 496971 152144
rect 494316 152086 496971 152088
rect 252277 152083 252343 152086
rect 496905 152083 496971 152086
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 213913 151947 213979 151950
rect 214649 151874 214715 151877
rect 307661 151874 307727 151877
rect 214649 151872 217058 151874
rect 214649 151816 214654 151872
rect 214710 151830 217058 151872
rect 307661 151872 310040 151874
rect 217182 151830 217242 151844
rect 214710 151816 217242 151830
rect 214649 151814 217242 151816
rect 214649 151811 214715 151814
rect 216998 151770 217242 151814
rect 307661 151816 307666 151872
rect 307722 151816 310040 151872
rect 307661 151814 310040 151816
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324957 151738 325023 151741
rect 248952 151736 252527 151738
rect 248952 151680 252466 151736
rect 252522 151680 252527 151736
rect 248952 151678 252527 151680
rect 321908 151736 325023 151738
rect 321908 151680 324962 151736
rect 325018 151680 325023 151736
rect 321908 151678 325023 151680
rect 252461 151675 252527 151678
rect 324957 151675 325023 151678
rect 416773 151602 416839 151605
rect 416773 151600 420164 151602
rect 416773 151544 416778 151600
rect 416834 151544 420164 151600
rect 416773 151542 420164 151544
rect 416773 151539 416839 151542
rect 307293 151466 307359 151469
rect 307293 151464 310040 151466
rect 307293 151408 307298 151464
rect 307354 151408 310040 151464
rect 307293 151406 310040 151408
rect 307293 151403 307359 151406
rect 252277 151194 252343 151197
rect 248952 151192 252343 151194
rect 214005 150922 214071 150925
rect 217182 150922 217242 151164
rect 248952 151136 252282 151192
rect 252338 151136 252343 151192
rect 248952 151134 252343 151136
rect 252277 151131 252343 151134
rect 306925 151058 306991 151061
rect 306925 151056 310040 151058
rect 306925 151000 306930 151056
rect 306986 151000 310040 151056
rect 306925 150998 310040 151000
rect 306925 150995 306991 150998
rect 324313 150922 324379 150925
rect 496813 150922 496879 150925
rect 214005 150920 217242 150922
rect 214005 150864 214010 150920
rect 214066 150864 217242 150920
rect 214005 150862 217242 150864
rect 321908 150920 324379 150922
rect 321908 150864 324318 150920
rect 324374 150864 324379 150920
rect 321908 150862 324379 150864
rect 494316 150920 496879 150922
rect 494316 150864 496818 150920
rect 496874 150864 496879 150920
rect 494316 150862 496879 150864
rect 214005 150859 214071 150862
rect 324313 150859 324379 150862
rect 496813 150859 496879 150862
rect 252369 150786 252435 150789
rect 248952 150784 252435 150786
rect 248952 150728 252374 150784
rect 252430 150728 252435 150784
rect 248952 150726 252435 150728
rect 252369 150723 252435 150726
rect 213913 150650 213979 150653
rect 307661 150650 307727 150653
rect 213913 150648 217242 150650
rect 213913 150592 213918 150648
rect 213974 150592 217242 150648
rect 213913 150590 217242 150592
rect 213913 150587 213979 150590
rect 217182 150484 217242 150590
rect 307661 150648 310040 150650
rect 307661 150592 307666 150648
rect 307722 150592 310040 150648
rect 307661 150590 310040 150592
rect 307661 150587 307727 150590
rect 252461 150242 252527 150245
rect 248952 150240 252527 150242
rect 248952 150184 252466 150240
rect 252522 150184 252527 150240
rect 248952 150182 252527 150184
rect 252461 150179 252527 150182
rect 306557 150242 306623 150245
rect 306557 150240 310040 150242
rect 306557 150184 306562 150240
rect 306618 150184 310040 150240
rect 306557 150182 310040 150184
rect 306557 150179 306623 150182
rect 214005 150106 214071 150109
rect 324313 150106 324379 150109
rect 214005 150104 217242 150106
rect 214005 150048 214010 150104
rect 214066 150048 217242 150104
rect 214005 150046 217242 150048
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 214005 150043 214071 150046
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150046
rect 324313 150043 324379 150046
rect 252277 149834 252343 149837
rect 248952 149832 252343 149834
rect -960 149774 3483 149776
rect 248952 149776 252282 149832
rect 252338 149776 252343 149832
rect 248952 149774 252343 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 252277 149771 252343 149774
rect 306925 149834 306991 149837
rect 416773 149834 416839 149837
rect 496813 149834 496879 149837
rect 306925 149832 310040 149834
rect 306925 149776 306930 149832
rect 306986 149776 310040 149832
rect 306925 149774 310040 149776
rect 416773 149832 420164 149834
rect 416773 149776 416778 149832
rect 416834 149776 420164 149832
rect 416773 149774 420164 149776
rect 494316 149832 496879 149834
rect 494316 149776 496818 149832
rect 496874 149776 496879 149832
rect 494316 149774 496879 149776
rect 306925 149771 306991 149774
rect 416773 149771 416839 149774
rect 496813 149771 496879 149774
rect 251766 149636 251772 149700
rect 251836 149698 251842 149700
rect 286409 149698 286475 149701
rect 251836 149696 286475 149698
rect 251836 149640 286414 149696
rect 286470 149640 286475 149696
rect 251836 149638 286475 149640
rect 251836 149636 251842 149638
rect 286409 149635 286475 149638
rect 324497 149698 324563 149701
rect 326654 149698 326660 149700
rect 324497 149696 326660 149698
rect 324497 149640 324502 149696
rect 324558 149640 326660 149696
rect 324497 149638 326660 149640
rect 324497 149635 324563 149638
rect 326654 149636 326660 149638
rect 326724 149636 326730 149700
rect 214557 149562 214623 149565
rect 214557 149560 217242 149562
rect 214557 149504 214562 149560
rect 214618 149504 217242 149560
rect 214557 149502 217242 149504
rect 214557 149499 214623 149502
rect 217182 149124 217242 149502
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 249149 149290 249215 149293
rect 248952 149288 249215 149290
rect 248952 149232 249154 149288
rect 249210 149232 249215 149288
rect 248952 149230 249215 149232
rect 249149 149227 249215 149230
rect 307293 149290 307359 149293
rect 307293 149288 310040 149290
rect 307293 149232 307298 149288
rect 307354 149232 310040 149288
rect 307293 149230 310040 149232
rect 307293 149227 307359 149230
rect 252369 148882 252435 148885
rect 248952 148880 252435 148882
rect 248952 148824 252374 148880
rect 252430 148824 252435 148880
rect 248952 148822 252435 148824
rect 252369 148819 252435 148822
rect 307477 148882 307543 148885
rect 307477 148880 310040 148882
rect 307477 148824 307482 148880
rect 307538 148824 310040 148880
rect 307477 148822 310040 148824
rect 307477 148819 307543 148822
rect 213913 148746 213979 148749
rect 496813 148746 496879 148749
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 494316 148744 496879 148746
rect 494316 148688 496818 148744
rect 496874 148688 496879 148744
rect 494316 148686 496879 148688
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 496813 148683 496879 148686
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 307569 148474 307635 148477
rect 307569 148472 310040 148474
rect 307569 148416 307574 148472
rect 307630 148416 310040 148472
rect 307569 148414 310040 148416
rect 307569 148411 307635 148414
rect 252461 148338 252527 148341
rect 248952 148336 252527 148338
rect 248952 148280 252466 148336
rect 252522 148280 252527 148336
rect 248952 148278 252527 148280
rect 252461 148275 252527 148278
rect 340086 148276 340092 148340
rect 340156 148338 340162 148340
rect 369853 148338 369919 148341
rect 340156 148336 369919 148338
rect 340156 148280 369858 148336
rect 369914 148280 369919 148336
rect 340156 148278 369919 148280
rect 340156 148276 340162 148278
rect 369853 148275 369919 148278
rect 416773 148202 416839 148205
rect 416773 148200 420164 148202
rect 416773 148144 416778 148200
rect 416834 148144 420164 148200
rect 416773 148142 420164 148144
rect 416773 148139 416839 148142
rect 214557 148066 214623 148069
rect 269062 148066 269068 148068
rect 214557 148064 217242 148066
rect 214557 148008 214562 148064
rect 214618 148008 217242 148064
rect 214557 148006 217242 148008
rect 214557 148003 214623 148006
rect 217182 147900 217242 148006
rect 258030 148006 269068 148066
rect 258030 147930 258090 148006
rect 269062 148004 269068 148006
rect 269132 148004 269138 148068
rect 307661 148066 307727 148069
rect 307661 148064 310040 148066
rect 307661 148008 307666 148064
rect 307722 148008 310040 148064
rect 307661 148006 310040 148008
rect 307661 148003 307727 148006
rect 248952 147870 258090 147930
rect 324405 147794 324471 147797
rect 321908 147792 324471 147794
rect 321908 147736 324410 147792
rect 324466 147736 324471 147792
rect 321908 147734 324471 147736
rect 324405 147731 324471 147734
rect 306925 147658 306991 147661
rect 496813 147658 496879 147661
rect 306925 147656 310040 147658
rect 306925 147600 306930 147656
rect 306986 147600 310040 147656
rect 306925 147598 310040 147600
rect 494316 147656 496879 147658
rect 494316 147600 496818 147656
rect 496874 147600 496879 147656
rect 494316 147598 496879 147600
rect 306925 147595 306991 147598
rect 496813 147595 496879 147598
rect 252461 147522 252527 147525
rect 248952 147520 252527 147522
rect 248952 147464 252466 147520
rect 252522 147464 252527 147520
rect 248952 147462 252527 147464
rect 252461 147459 252527 147462
rect 307477 147250 307543 147253
rect 307477 147248 310040 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 307477 147192 307482 147248
rect 307538 147192 310040 147248
rect 307477 147190 310040 147192
rect 307477 147187 307543 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 252093 146978 252159 146981
rect 248952 146976 252159 146978
rect 248952 146920 252098 146976
rect 252154 146920 252159 146976
rect 248952 146918 252159 146920
rect 252093 146915 252159 146918
rect 307569 146842 307635 146845
rect 307569 146840 310040 146842
rect 307569 146784 307574 146840
rect 307630 146784 310040 146840
rect 307569 146782 310040 146784
rect 307569 146779 307635 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 214005 146643 214071 146646
rect 254526 146570 254532 146572
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 248952 146510 254532 146570
rect 254526 146508 254532 146510
rect 254596 146508 254602 146572
rect 416773 146570 416839 146573
rect 416773 146568 420164 146570
rect 416773 146512 416778 146568
rect 416834 146512 420164 146568
rect 416773 146510 420164 146512
rect 416773 146507 416839 146510
rect 307661 146434 307727 146437
rect 495709 146434 495775 146437
rect 307661 146432 310040 146434
rect 307661 146376 307666 146432
rect 307722 146376 310040 146432
rect 307661 146374 310040 146376
rect 494316 146432 495775 146434
rect 494316 146376 495714 146432
rect 495770 146376 495775 146432
rect 494316 146374 495775 146376
rect 307661 146371 307727 146374
rect 495709 146371 495775 146374
rect 324313 146298 324379 146301
rect 216814 146238 217426 146298
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 252461 146026 252527 146029
rect 248952 146024 252527 146026
rect 248952 145968 252466 146024
rect 252522 145968 252527 146024
rect 248952 145966 252527 145968
rect 252461 145963 252527 145966
rect 307477 145890 307543 145893
rect 307477 145888 310040 145890
rect 217182 145346 217242 145860
rect 307477 145832 307482 145888
rect 307538 145832 310040 145888
rect 307477 145830 310040 145832
rect 307477 145827 307543 145830
rect 252369 145618 252435 145621
rect 248952 145616 252435 145618
rect 248952 145560 252374 145616
rect 252430 145560 252435 145616
rect 248952 145558 252435 145560
rect 252369 145555 252435 145558
rect 306925 145482 306991 145485
rect 324405 145482 324471 145485
rect 306925 145480 310040 145482
rect 306925 145424 306930 145480
rect 306986 145424 310040 145480
rect 306925 145422 310040 145424
rect 321908 145480 324471 145482
rect 321908 145424 324410 145480
rect 324466 145424 324471 145480
rect 321908 145422 324471 145424
rect 306925 145419 306991 145422
rect 324405 145419 324471 145422
rect 496813 145346 496879 145349
rect 200070 145286 217242 145346
rect 494316 145344 496879 145346
rect 494316 145288 496818 145344
rect 496874 145288 496879 145344
rect 494316 145286 496879 145288
rect 168966 144876 168972 144940
rect 169036 144938 169042 144940
rect 200070 144938 200130 145286
rect 496813 145283 496879 145286
rect 169036 144878 200130 144938
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 259494 145074 259500 145076
rect 248952 145014 259500 145074
rect 259494 145012 259500 145014
rect 259564 145012 259570 145076
rect 307385 145074 307451 145077
rect 307385 145072 310040 145074
rect 307385 145016 307390 145072
rect 307446 145016 310040 145072
rect 307385 145014 310040 145016
rect 307385 145011 307451 145014
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 169036 144876 169042 144878
rect 213913 144875 213979 144878
rect 252502 144666 252508 144668
rect 248952 144606 252508 144666
rect 252502 144604 252508 144606
rect 252572 144604 252578 144668
rect 306557 144666 306623 144669
rect 306557 144664 310040 144666
rect 306557 144608 306562 144664
rect 306618 144608 310040 144664
rect 306557 144606 310040 144608
rect 306557 144603 306623 144606
rect 214649 143986 214715 143989
rect 217182 143986 217242 144500
rect 307661 144258 307727 144261
rect 307661 144256 310040 144258
rect 307661 144200 307666 144256
rect 307722 144200 310040 144256
rect 307661 144198 310040 144200
rect 307661 144195 307727 144198
rect 252461 144122 252527 144125
rect 248952 144120 252527 144122
rect 248952 144064 252466 144120
rect 252522 144064 252527 144120
rect 248952 144062 252527 144064
rect 321878 144122 321938 144772
rect 336038 144740 336044 144804
rect 336108 144802 336114 144804
rect 342345 144802 342411 144805
rect 336108 144800 342411 144802
rect 336108 144744 342350 144800
rect 342406 144744 342411 144800
rect 336108 144742 342411 144744
rect 336108 144740 336114 144742
rect 342345 144739 342411 144742
rect 416865 144802 416931 144805
rect 416865 144800 420164 144802
rect 416865 144744 416870 144800
rect 416926 144744 420164 144800
rect 416865 144742 420164 144744
rect 416865 144739 416931 144742
rect 496813 144258 496879 144261
rect 494316 144256 496879 144258
rect 494316 144200 496818 144256
rect 496874 144200 496879 144256
rect 494316 144198 496879 144200
rect 496813 144195 496879 144198
rect 331438 144122 331444 144124
rect 321878 144062 331444 144122
rect 252461 144059 252527 144062
rect 331438 144060 331444 144062
rect 331508 144060 331514 144124
rect 325785 143986 325851 143989
rect 214649 143984 217242 143986
rect 214649 143928 214654 143984
rect 214710 143928 217242 143984
rect 214649 143926 217242 143928
rect 321908 143984 325851 143986
rect 321908 143928 325790 143984
rect 325846 143928 325851 143984
rect 321908 143926 325851 143928
rect 214649 143923 214715 143926
rect 325785 143923 325851 143926
rect 307293 143850 307359 143853
rect 307293 143848 310040 143850
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 307293 143792 307298 143848
rect 307354 143792 310040 143848
rect 307293 143790 310040 143792
rect 307293 143787 307359 143790
rect 252369 143714 252435 143717
rect 248952 143712 252435 143714
rect 248952 143656 252374 143712
rect 252430 143656 252435 143712
rect 248952 143654 252435 143656
rect 252369 143651 252435 143654
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 213913 143515 213979 143518
rect 307569 143442 307635 143445
rect 307569 143440 310040 143442
rect 307569 143384 307574 143440
rect 307630 143384 310040 143440
rect 307569 143382 310040 143384
rect 307569 143379 307635 143382
rect 213913 142762 213979 142765
rect 217182 142762 217242 143276
rect 252461 143170 252527 143173
rect 324313 143170 324379 143173
rect 248952 143168 252527 143170
rect 248952 143112 252466 143168
rect 252522 143112 252527 143168
rect 248952 143110 252527 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 252461 143107 252527 143110
rect 324313 143107 324379 143110
rect 416773 143170 416839 143173
rect 496905 143170 496971 143173
rect 416773 143168 420164 143170
rect 416773 143112 416778 143168
rect 416834 143112 420164 143168
rect 416773 143110 420164 143112
rect 494316 143168 496971 143170
rect 494316 143112 496910 143168
rect 496966 143112 496971 143168
rect 494316 143110 496971 143112
rect 416773 143107 416839 143110
rect 496905 143107 496971 143110
rect 307661 143034 307727 143037
rect 307661 143032 310040 143034
rect 307661 142976 307666 143032
rect 307722 142976 310040 143032
rect 307661 142974 310040 142976
rect 307661 142971 307727 142974
rect 252369 142762 252435 142765
rect 213913 142760 217242 142762
rect 213913 142704 213918 142760
rect 213974 142704 217242 142760
rect 213913 142702 217242 142704
rect 248952 142760 252435 142762
rect 248952 142704 252374 142760
rect 252430 142704 252435 142760
rect 248952 142702 252435 142704
rect 213913 142699 213979 142702
rect 252369 142699 252435 142702
rect 214465 142354 214531 142357
rect 217366 142354 217426 142596
rect 307201 142490 307267 142493
rect 324497 142490 324563 142493
rect 307201 142488 310040 142490
rect 307201 142432 307206 142488
rect 307262 142432 310040 142488
rect 307201 142430 310040 142432
rect 321908 142488 324563 142490
rect 321908 142432 324502 142488
rect 324558 142432 324563 142488
rect 321908 142430 324563 142432
rect 307201 142427 307267 142430
rect 324497 142427 324563 142430
rect 214465 142352 217426 142354
rect 214465 142296 214470 142352
rect 214526 142296 217426 142352
rect 214465 142294 217426 142296
rect 214465 142291 214531 142294
rect 266302 142218 266308 142220
rect 248952 142158 266308 142218
rect 266302 142156 266308 142158
rect 266372 142156 266378 142220
rect 307569 142082 307635 142085
rect 307569 142080 310040 142082
rect 307569 142024 307574 142080
rect 307630 142024 310040 142080
rect 307569 142022 310040 142024
rect 307569 142019 307635 142022
rect 496813 141946 496879 141949
rect 494316 141944 496879 141946
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 494316 141888 496818 141944
rect 496874 141888 496879 141944
rect 494316 141886 496879 141888
rect 496813 141883 496879 141886
rect 253565 141810 253631 141813
rect 248952 141808 253631 141810
rect 248952 141752 253570 141808
rect 253626 141752 253631 141808
rect 248952 141750 253631 141752
rect 253565 141747 253631 141750
rect 306833 141674 306899 141677
rect 324313 141674 324379 141677
rect 306833 141672 310040 141674
rect 306833 141616 306838 141672
rect 306894 141616 310040 141672
rect 306833 141614 310040 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 306833 141611 306899 141614
rect 324313 141611 324379 141614
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 416773 141402 416839 141405
rect 416773 141400 420164 141402
rect 214005 141342 217242 141344
rect 214005 141339 214071 141342
rect 248860 141298 249442 141358
rect 416773 141344 416778 141400
rect 416834 141344 420164 141400
rect 416773 141342 420164 141344
rect 416773 141339 416839 141342
rect 213913 140858 213979 140861
rect 217182 140858 217242 141236
rect 249382 140994 249442 141298
rect 306966 141204 306972 141268
rect 307036 141266 307042 141268
rect 307036 141206 310040 141266
rect 307036 141204 307042 141206
rect 253289 141130 253355 141133
rect 255446 141130 255452 141132
rect 253289 141128 255452 141130
rect 253289 141072 253294 141128
rect 253350 141072 255452 141128
rect 253289 141070 255452 141072
rect 253289 141067 253355 141070
rect 255446 141068 255452 141070
rect 255516 141068 255522 141132
rect 259678 140994 259684 140996
rect 249382 140934 259684 140994
rect 259678 140932 259684 140934
rect 259748 140932 259754 140996
rect 253289 140858 253355 140861
rect 213913 140856 217242 140858
rect 213913 140800 213918 140856
rect 213974 140800 217242 140856
rect 213913 140798 217242 140800
rect 248952 140856 253355 140858
rect 248952 140800 253294 140856
rect 253350 140800 253355 140856
rect 248952 140798 253355 140800
rect 213913 140795 213979 140798
rect 253289 140795 253355 140798
rect 253565 140858 253631 140861
rect 263542 140858 263548 140860
rect 253565 140856 263548 140858
rect 253565 140800 253570 140856
rect 253626 140800 263548 140856
rect 253565 140798 263548 140800
rect 253565 140795 253631 140798
rect 263542 140796 263548 140798
rect 263612 140796 263618 140860
rect 307661 140858 307727 140861
rect 324405 140858 324471 140861
rect 496813 140858 496879 140861
rect 307661 140856 310040 140858
rect 307661 140800 307666 140856
rect 307722 140800 310040 140856
rect 307661 140798 310040 140800
rect 321908 140856 324471 140858
rect 321908 140800 324410 140856
rect 324466 140800 324471 140856
rect 321908 140798 324471 140800
rect 494316 140856 496879 140858
rect 494316 140800 496818 140856
rect 496874 140800 496879 140856
rect 494316 140798 496879 140800
rect 307661 140795 307727 140798
rect 324405 140795 324471 140798
rect 496813 140795 496879 140798
rect 214005 140042 214071 140045
rect 217182 140042 217242 140556
rect 252461 140450 252527 140453
rect 248952 140448 252527 140450
rect 248952 140392 252466 140448
rect 252522 140392 252527 140448
rect 248952 140390 252527 140392
rect 252461 140387 252527 140390
rect 307477 140450 307543 140453
rect 307477 140448 310040 140450
rect 307477 140392 307482 140448
rect 307538 140392 310040 140448
rect 307477 140390 310040 140392
rect 307477 140387 307543 140390
rect 214005 140040 217242 140042
rect 214005 139984 214010 140040
rect 214066 139984 217242 140040
rect 214005 139982 217242 139984
rect 307569 140042 307635 140045
rect 307569 140040 310040 140042
rect 307569 139984 307574 140040
rect 307630 139984 310040 140040
rect 307569 139982 310040 139984
rect 214005 139979 214071 139982
rect 307569 139979 307635 139982
rect 252369 139906 252435 139909
rect 248952 139904 252435 139906
rect 213913 139498 213979 139501
rect 217182 139498 217242 139876
rect 248952 139848 252374 139904
rect 252430 139848 252435 139904
rect 248952 139846 252435 139848
rect 252369 139843 252435 139846
rect 307661 139634 307727 139637
rect 307661 139632 310040 139634
rect 307661 139576 307666 139632
rect 307722 139576 310040 139632
rect 307661 139574 310040 139576
rect 307661 139571 307727 139574
rect 249793 139498 249859 139501
rect 213913 139496 217242 139498
rect 213913 139440 213918 139496
rect 213974 139440 217242 139496
rect 213913 139438 217242 139440
rect 248952 139496 249859 139498
rect 248952 139440 249798 139496
rect 249854 139440 249859 139496
rect 248952 139438 249859 139440
rect 321878 139498 321938 140148
rect 416773 139770 416839 139773
rect 496813 139770 496879 139773
rect 416773 139768 420164 139770
rect 416773 139712 416778 139768
rect 416834 139712 420164 139768
rect 416773 139710 420164 139712
rect 494316 139768 496879 139770
rect 494316 139712 496818 139768
rect 496874 139712 496879 139768
rect 494316 139710 496879 139712
rect 416773 139707 416839 139710
rect 496813 139707 496879 139710
rect 330334 139498 330340 139500
rect 321878 139438 330340 139498
rect 213913 139435 213979 139438
rect 249793 139435 249859 139438
rect 330334 139436 330340 139438
rect 330404 139436 330410 139500
rect 327022 139362 327028 139364
rect 321908 139302 327028 139362
rect 327022 139300 327028 139302
rect 327092 139300 327098 139364
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 214005 138818 214071 138821
rect 217182 138818 217242 139196
rect 309504 138986 310132 139046
rect 248860 138850 249442 138910
rect 214005 138816 217242 138818
rect 214005 138760 214010 138816
rect 214066 138760 217242 138816
rect 214005 138758 217242 138760
rect 214005 138755 214071 138758
rect 249382 138682 249442 138850
rect 213913 138138 213979 138141
rect 217182 138138 217242 138652
rect 249382 138622 253490 138682
rect 252461 138546 252527 138549
rect 248952 138544 252527 138546
rect 248952 138488 252466 138544
rect 252522 138488 252527 138544
rect 248952 138486 252527 138488
rect 252461 138483 252527 138486
rect 253430 138274 253490 138622
rect 253606 138348 253612 138412
rect 253676 138410 253682 138412
rect 309504 138410 309564 138986
rect 309685 138682 309751 138685
rect 496813 138682 496879 138685
rect 309685 138680 310040 138682
rect 309685 138624 309690 138680
rect 309746 138624 310040 138680
rect 309685 138622 310040 138624
rect 494316 138680 496879 138682
rect 494316 138624 496818 138680
rect 496874 138624 496879 138680
rect 494316 138622 496879 138624
rect 309685 138619 309751 138622
rect 496813 138619 496879 138622
rect 324313 138546 324379 138549
rect 321908 138544 324379 138546
rect 321908 138488 324318 138544
rect 324374 138488 324379 138544
rect 321908 138486 324379 138488
rect 324313 138483 324379 138486
rect 253676 138350 309564 138410
rect 253676 138348 253682 138350
rect 262254 138274 262260 138276
rect 253430 138214 262260 138274
rect 262254 138212 262260 138214
rect 262324 138212 262330 138276
rect 307661 138274 307727 138277
rect 307661 138272 310040 138274
rect 307661 138216 307666 138272
rect 307722 138216 310040 138272
rect 307661 138214 310040 138216
rect 307661 138211 307727 138214
rect 213913 138136 217242 138138
rect 213913 138080 213918 138136
rect 213974 138080 217242 138136
rect 213913 138078 217242 138080
rect 307569 138138 307635 138141
rect 309685 138138 309751 138141
rect 307569 138136 309751 138138
rect 307569 138080 307574 138136
rect 307630 138080 309690 138136
rect 309746 138080 309751 138136
rect 307569 138078 309751 138080
rect 213913 138075 213979 138078
rect 307569 138075 307635 138078
rect 309685 138075 309751 138078
rect 252461 138002 252527 138005
rect 248952 138000 252527 138002
rect 213913 137458 213979 137461
rect 217182 137458 217242 137972
rect 248952 137944 252466 138000
rect 252522 137944 252527 138000
rect 248952 137942 252527 137944
rect 252461 137939 252527 137942
rect 416773 138002 416839 138005
rect 416773 138000 420164 138002
rect 416773 137944 416778 138000
rect 416834 137944 420164 138000
rect 416773 137942 420164 137944
rect 416773 137939 416839 137942
rect 307661 137866 307727 137869
rect 324313 137866 324379 137869
rect 307661 137864 310040 137866
rect 307661 137808 307666 137864
rect 307722 137808 310040 137864
rect 307661 137806 310040 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307661 137803 307727 137806
rect 324313 137803 324379 137806
rect 252369 137594 252435 137597
rect 248952 137592 252435 137594
rect 248952 137536 252374 137592
rect 252430 137536 252435 137592
rect 248952 137534 252435 137536
rect 252369 137531 252435 137534
rect 213913 137456 217242 137458
rect 213913 137400 213918 137456
rect 213974 137400 217242 137456
rect 213913 137398 217242 137400
rect 307109 137458 307175 137461
rect 496813 137458 496879 137461
rect 307109 137456 310040 137458
rect 307109 137400 307114 137456
rect 307170 137400 310040 137456
rect 307109 137398 310040 137400
rect 494316 137456 496879 137458
rect 494316 137400 496818 137456
rect 496874 137400 496879 137456
rect 494316 137398 496879 137400
rect 213913 137395 213979 137398
rect 307109 137395 307175 137398
rect 496813 137395 496879 137398
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 170438 136716 170444 136780
rect 170508 136778 170514 136780
rect 217182 136778 217242 137292
rect 249885 137050 249951 137053
rect 248952 137048 249951 137050
rect 248952 136992 249890 137048
rect 249946 136992 249951 137048
rect 248952 136990 249951 136992
rect 249885 136987 249951 136990
rect 307017 137050 307083 137053
rect 324405 137050 324471 137053
rect 307017 137048 310040 137050
rect 307017 136992 307022 137048
rect 307078 136992 310040 137048
rect 307017 136990 310040 136992
rect 321908 137048 324471 137050
rect 321908 136992 324410 137048
rect 324466 136992 324471 137048
rect 321908 136990 324471 136992
rect 307017 136987 307083 136990
rect 324405 136987 324471 136990
rect 170508 136718 217242 136778
rect 170508 136716 170514 136718
rect 252461 136642 252527 136645
rect 248952 136640 252527 136642
rect 170254 136036 170260 136100
rect 170324 136098 170330 136100
rect 214005 136098 214071 136101
rect 217182 136098 217242 136612
rect 248952 136584 252466 136640
rect 252522 136584 252527 136640
rect 248952 136582 252527 136584
rect 252461 136579 252527 136582
rect 307477 136642 307543 136645
rect 307477 136640 310040 136642
rect 307477 136584 307482 136640
rect 307538 136584 310040 136640
rect 307477 136582 310040 136584
rect 307477 136579 307543 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 416773 136370 416839 136373
rect 496813 136370 496879 136373
rect 416773 136368 420164 136370
rect 416773 136312 416778 136368
rect 416834 136312 420164 136368
rect 416773 136310 420164 136312
rect 494316 136368 496879 136370
rect 494316 136312 496818 136368
rect 496874 136312 496879 136368
rect 494316 136310 496879 136312
rect 416773 136307 416839 136310
rect 496813 136307 496879 136310
rect 252369 136234 252435 136237
rect 248952 136232 252435 136234
rect 248952 136176 252374 136232
rect 252430 136176 252435 136232
rect 248952 136174 252435 136176
rect 252369 136171 252435 136174
rect 307109 136234 307175 136237
rect 307109 136232 310040 136234
rect 307109 136176 307114 136232
rect 307170 136176 310040 136232
rect 307109 136174 310040 136176
rect 307109 136171 307175 136174
rect 170324 136038 200130 136098
rect 170324 136036 170330 136038
rect 200070 135554 200130 136038
rect 214005 136096 217242 136098
rect 214005 136040 214010 136096
rect 214066 136040 217242 136096
rect 214005 136038 217242 136040
rect 214005 136035 214071 136038
rect 213913 135690 213979 135693
rect 217182 135690 217242 135932
rect 252185 135690 252251 135693
rect 213913 135688 217242 135690
rect 213913 135632 213918 135688
rect 213974 135632 217242 135688
rect 213913 135630 217242 135632
rect 248952 135688 252251 135690
rect 248952 135632 252190 135688
rect 252246 135632 252251 135688
rect 248952 135630 252251 135632
rect 213913 135627 213979 135630
rect 252185 135627 252251 135630
rect 307569 135690 307635 135693
rect 307569 135688 310040 135690
rect 307569 135632 307574 135688
rect 307630 135632 310040 135688
rect 307569 135630 310040 135632
rect 307569 135627 307635 135630
rect 217317 135554 217383 135557
rect 323301 135554 323367 135557
rect 200070 135552 217383 135554
rect 200070 135496 217322 135552
rect 217378 135496 217383 135552
rect 200070 135494 217383 135496
rect 321908 135552 323367 135554
rect 321908 135496 323306 135552
rect 323362 135496 323367 135552
rect 321908 135494 323367 135496
rect 217317 135491 217383 135494
rect 323301 135491 323367 135494
rect 200070 135358 217242 135418
rect 169150 135220 169156 135284
rect 169220 135282 169226 135284
rect 200070 135282 200130 135358
rect 169220 135222 200130 135282
rect 217182 135252 217242 135358
rect 252277 135282 252343 135285
rect 248952 135280 252343 135282
rect 248952 135224 252282 135280
rect 252338 135224 252343 135280
rect 248952 135222 252343 135224
rect 169220 135220 169226 135222
rect 252277 135219 252343 135222
rect 307661 135282 307727 135285
rect 496905 135282 496971 135285
rect 307661 135280 310040 135282
rect 307661 135224 307666 135280
rect 307722 135224 310040 135280
rect 307661 135222 310040 135224
rect 494316 135280 496971 135282
rect 494316 135224 496910 135280
rect 496966 135224 496971 135280
rect 494316 135222 496971 135224
rect 307661 135219 307727 135222
rect 496905 135219 496971 135222
rect 307569 134874 307635 134877
rect 307569 134872 310040 134874
rect 307569 134816 307574 134872
rect 307630 134816 310040 134872
rect 307569 134814 310040 134816
rect 307569 134811 307635 134814
rect 252461 134738 252527 134741
rect 324313 134738 324379 134741
rect 494145 134738 494211 134741
rect 248952 134736 252527 134738
rect 248952 134680 252466 134736
rect 252522 134680 252527 134736
rect 248952 134678 252527 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 252461 134675 252527 134678
rect 324313 134675 324379 134678
rect 494102 134736 494211 134738
rect 494102 134680 494150 134736
rect 494206 134680 494211 134736
rect 494102 134675 494211 134680
rect 417325 134602 417391 134605
rect 419165 134602 419231 134605
rect 417325 134600 420164 134602
rect 214741 134194 214807 134197
rect 217182 134194 217242 134572
rect 417325 134544 417330 134600
rect 417386 134544 419170 134600
rect 419226 134544 420164 134600
rect 417325 134542 420164 134544
rect 417325 134539 417391 134542
rect 419165 134539 419231 134542
rect 307661 134466 307727 134469
rect 307661 134464 310040 134466
rect 307661 134408 307666 134464
rect 307722 134408 310040 134464
rect 307661 134406 310040 134408
rect 307661 134403 307727 134406
rect 252369 134330 252435 134333
rect 248952 134328 252435 134330
rect 248952 134272 252374 134328
rect 252430 134272 252435 134328
rect 248952 134270 252435 134272
rect 252369 134267 252435 134270
rect 214741 134192 217242 134194
rect 214741 134136 214746 134192
rect 214802 134136 217242 134192
rect 214741 134134 217242 134136
rect 214741 134131 214807 134134
rect 257286 134132 257292 134196
rect 257356 134194 257362 134196
rect 257356 134134 296730 134194
rect 494102 134164 494162 134675
rect 257356 134132 257362 134134
rect 213913 134058 213979 134061
rect 296670 134058 296730 134134
rect 324405 134058 324471 134061
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 296670 133998 310040 134058
rect 321908 134056 324471 134058
rect 321908 134000 324410 134056
rect 324466 134000 324471 134056
rect 321908 133998 324471 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 324405 133995 324471 133998
rect 252461 133786 252527 133789
rect 248952 133784 252527 133786
rect 248952 133728 252466 133784
rect 252522 133728 252527 133784
rect 248952 133726 252527 133728
rect 252461 133723 252527 133726
rect 307569 133650 307635 133653
rect 307569 133648 310040 133650
rect 307569 133592 307574 133648
rect 307630 133592 310040 133648
rect 307569 133590 310040 133592
rect 307569 133587 307635 133590
rect 252369 133378 252435 133381
rect 248952 133376 252435 133378
rect 166390 132772 166396 132836
rect 166460 132834 166466 132836
rect 217182 132834 217242 133348
rect 248952 133320 252374 133376
rect 252430 133320 252435 133376
rect 248952 133318 252435 133320
rect 252369 133315 252435 133318
rect 306925 133242 306991 133245
rect 324313 133242 324379 133245
rect 306925 133240 310040 133242
rect 306925 133184 306930 133240
rect 306986 133184 310040 133240
rect 306925 133182 310040 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 306925 133179 306991 133182
rect 324313 133179 324379 133182
rect 419349 132970 419415 132973
rect 496813 132970 496879 132973
rect 419349 132968 420164 132970
rect 419349 132912 419354 132968
rect 419410 132912 420164 132968
rect 419349 132910 420164 132912
rect 494316 132968 496879 132970
rect 494316 132912 496818 132968
rect 496874 132912 496879 132968
rect 494316 132910 496879 132912
rect 419349 132907 419415 132910
rect 496813 132907 496879 132910
rect 252093 132834 252159 132837
rect 166460 132774 217242 132834
rect 248952 132832 252159 132834
rect 248952 132776 252098 132832
rect 252154 132776 252159 132832
rect 248952 132774 252159 132776
rect 166460 132772 166466 132774
rect 252093 132771 252159 132774
rect 170254 132636 170260 132700
rect 170324 132698 170330 132700
rect 307661 132698 307727 132701
rect 321553 132698 321619 132701
rect 170324 132638 217058 132698
rect 307661 132696 310040 132698
rect 170324 132636 170330 132638
rect 216998 132510 217058 132638
rect 217366 132510 217426 132668
rect 307661 132640 307666 132696
rect 307722 132640 310040 132696
rect 307661 132638 310040 132640
rect 321510 132696 321619 132698
rect 321510 132640 321558 132696
rect 321614 132640 321619 132696
rect 307661 132635 307727 132638
rect 321510 132635 321619 132640
rect 216998 132450 217426 132510
rect 252461 132426 252527 132429
rect 248952 132424 252527 132426
rect 248952 132368 252466 132424
rect 252522 132368 252527 132424
rect 321510 132396 321570 132635
rect 248952 132366 252527 132368
rect 252461 132363 252527 132366
rect 306557 132290 306623 132293
rect 306557 132288 310040 132290
rect 306557 132232 306562 132288
rect 306618 132232 310040 132288
rect 306557 132230 310040 132232
rect 306557 132227 306623 132230
rect 494329 132154 494395 132157
rect 494286 132152 494395 132154
rect 494286 132096 494334 132152
rect 494390 132096 494395 132152
rect 494286 132091 494395 132096
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 252369 131882 252435 131885
rect 248952 131880 252435 131882
rect 248952 131824 252374 131880
rect 252430 131824 252435 131880
rect 248952 131822 252435 131824
rect 252369 131819 252435 131822
rect 307661 131882 307727 131885
rect 307661 131880 310040 131882
rect 307661 131824 307666 131880
rect 307722 131824 310040 131880
rect 494286 131852 494346 132091
rect 307661 131822 310040 131824
rect 307661 131819 307727 131822
rect 252461 131474 252527 131477
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 248952 131472 252527 131474
rect 248952 131416 252466 131472
rect 252522 131416 252527 131472
rect 248952 131414 252527 131416
rect 214005 131411 214071 131414
rect 252461 131411 252527 131414
rect 307569 131474 307635 131477
rect 307569 131472 310040 131474
rect 307569 131416 307574 131472
rect 307630 131416 310040 131472
rect 307569 131414 310040 131416
rect 307569 131411 307635 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 321878 131202 321938 131716
rect 417325 131338 417391 131341
rect 419717 131338 419783 131341
rect 417325 131336 420164 131338
rect 417325 131280 417330 131336
rect 417386 131280 419722 131336
rect 419778 131280 420164 131336
rect 417325 131278 420164 131280
rect 417325 131275 417391 131278
rect 419717 131275 419783 131278
rect 331254 131202 331260 131204
rect 321878 131142 331260 131202
rect 331254 131140 331260 131142
rect 331324 131140 331330 131204
rect 216814 131006 217426 131066
rect 307293 131066 307359 131069
rect 307293 131064 310040 131066
rect 307293 131008 307298 131064
rect 307354 131008 310040 131064
rect 307293 131006 310040 131008
rect 307293 131003 307359 131006
rect 321502 131004 321508 131068
rect 321572 131004 321578 131068
rect 252461 130930 252527 130933
rect 248952 130928 252527 130930
rect 248952 130872 252466 130928
rect 252522 130872 252527 130928
rect 321510 130900 321570 131004
rect 248952 130870 252527 130872
rect 252461 130867 252527 130870
rect 496813 130794 496879 130797
rect 494316 130792 496879 130794
rect 494316 130736 496818 130792
rect 496874 130736 496879 130792
rect 494316 130734 496879 130736
rect 496813 130731 496879 130734
rect 307569 130658 307635 130661
rect 307569 130656 310040 130658
rect 214005 130114 214071 130117
rect 217182 130114 217242 130628
rect 307569 130600 307574 130656
rect 307630 130600 310040 130656
rect 307569 130598 310040 130600
rect 307569 130595 307635 130598
rect 252461 130522 252527 130525
rect 248952 130520 252527 130522
rect 248952 130464 252466 130520
rect 252522 130464 252527 130520
rect 248952 130462 252527 130464
rect 252461 130459 252527 130462
rect 307661 130250 307727 130253
rect 307661 130248 310040 130250
rect 307661 130192 307666 130248
rect 307722 130192 310040 130248
rect 307661 130190 310040 130192
rect 307661 130187 307727 130190
rect 252369 130114 252435 130117
rect 324313 130114 324379 130117
rect 214005 130112 217242 130114
rect 214005 130056 214010 130112
rect 214066 130056 217242 130112
rect 214005 130054 217242 130056
rect 248952 130112 252435 130114
rect 248952 130056 252374 130112
rect 252430 130056 252435 130112
rect 248952 130054 252435 130056
rect 321908 130112 324379 130114
rect 321908 130056 324318 130112
rect 324374 130056 324379 130112
rect 321908 130054 324379 130056
rect 214005 130051 214071 130054
rect 252369 130051 252435 130054
rect 324313 130051 324379 130054
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 305494 129780 305500 129844
rect 305564 129842 305570 129844
rect 305564 129782 310040 129842
rect 305564 129780 305570 129782
rect 216814 129646 217426 129706
rect 321645 129706 321711 129709
rect 496813 129706 496879 129709
rect 321645 129704 321754 129706
rect 321645 129648 321650 129704
rect 321706 129648 321754 129704
rect 321645 129643 321754 129648
rect 494316 129704 496879 129706
rect 494316 129648 496818 129704
rect 496874 129648 496879 129704
rect 494316 129646 496879 129648
rect 496813 129643 496879 129646
rect 251909 129570 251975 129573
rect 248952 129568 251975 129570
rect 248952 129512 251914 129568
rect 251970 129512 251975 129568
rect 248952 129510 251975 129512
rect 251909 129507 251975 129510
rect 321694 129404 321754 129643
rect 419625 129570 419691 129573
rect 419625 129568 420164 129570
rect 419625 129512 419630 129568
rect 419686 129512 420164 129568
rect 419625 129510 420164 129512
rect 419625 129507 419691 129510
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 213453 128890 213519 128893
rect 217182 128890 217242 129268
rect 309550 129194 310132 129254
rect 252369 129162 252435 129165
rect 248952 129160 252435 129162
rect 248952 129104 252374 129160
rect 252430 129104 252435 129160
rect 248952 129102 252435 129104
rect 252369 129099 252435 129102
rect 213453 128888 217242 128890
rect 213453 128832 213458 128888
rect 213514 128832 217242 128888
rect 213453 128830 217242 128832
rect 213453 128827 213519 128830
rect 172094 128556 172100 128620
rect 172164 128618 172170 128620
rect 172164 128558 213746 128618
rect 172164 128556 172170 128558
rect 168230 128420 168236 128484
rect 168300 128482 168306 128484
rect 213453 128482 213519 128485
rect 168300 128480 213519 128482
rect 168300 128424 213458 128480
rect 213514 128424 213519 128480
rect 168300 128422 213519 128424
rect 213686 128482 213746 128558
rect 217366 128482 217426 128724
rect 255814 128692 255820 128756
rect 255884 128754 255890 128756
rect 309550 128754 309610 129194
rect 494053 129026 494119 129029
rect 494053 129024 494162 129026
rect 494053 128968 494058 129024
rect 494114 128968 494162 129024
rect 494053 128963 494162 128968
rect 255884 128694 309610 128754
rect 309734 128786 310132 128846
rect 255884 128692 255890 128694
rect 252461 128618 252527 128621
rect 248952 128616 252527 128618
rect 248952 128560 252466 128616
rect 252522 128560 252527 128616
rect 248952 128558 252527 128560
rect 252461 128555 252527 128558
rect 307569 128618 307635 128621
rect 309734 128618 309794 128786
rect 324313 128618 324379 128621
rect 307569 128616 309794 128618
rect 307569 128560 307574 128616
rect 307630 128560 309794 128616
rect 307569 128558 309794 128560
rect 321908 128616 324379 128618
rect 321908 128560 324318 128616
rect 324374 128560 324379 128616
rect 321908 128558 324379 128560
rect 307569 128555 307635 128558
rect 324313 128555 324379 128558
rect 213686 128422 217426 128482
rect 307661 128482 307727 128485
rect 307661 128480 310040 128482
rect 307661 128424 307666 128480
rect 307722 128424 310040 128480
rect 494102 128452 494162 128963
rect 307661 128422 310040 128424
rect 168300 128420 168306 128422
rect 213453 128419 213519 128422
rect 307661 128419 307727 128422
rect 252461 128210 252527 128213
rect 248952 128208 252527 128210
rect 248952 128152 252466 128208
rect 252522 128152 252527 128208
rect 248952 128150 252527 128152
rect 252461 128147 252527 128150
rect 67357 128074 67423 128077
rect 68142 128074 68816 128080
rect 67357 128072 68816 128074
rect 67357 128016 67362 128072
rect 67418 128020 68816 128072
rect 306557 128074 306623 128077
rect 306557 128072 310040 128074
rect 67418 128016 68202 128020
rect 67357 128014 68202 128016
rect 67357 128011 67423 128014
rect 217182 127530 217242 128044
rect 306557 128016 306562 128072
rect 306618 128016 310040 128072
rect 306557 128014 310040 128016
rect 306557 128011 306623 128014
rect 417601 127938 417667 127941
rect 419257 127938 419323 127941
rect 417601 127936 420164 127938
rect 417601 127880 417606 127936
rect 417662 127880 419262 127936
rect 419318 127880 420164 127936
rect 417601 127878 420164 127880
rect 417601 127875 417667 127878
rect 419257 127875 419323 127878
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252369 127666 252435 127669
rect 248952 127664 252435 127666
rect 248952 127608 252374 127664
rect 252430 127608 252435 127664
rect 248952 127606 252435 127608
rect 252369 127603 252435 127606
rect 307150 127604 307156 127668
rect 307220 127666 307226 127668
rect 307220 127606 310040 127666
rect 307220 127604 307226 127606
rect 200070 127470 217242 127530
rect 166206 127060 166212 127124
rect 166276 127122 166282 127124
rect 200070 127122 200130 127470
rect 496813 127394 496879 127397
rect 494316 127392 496879 127394
rect 166276 127062 200130 127122
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 494316 127336 496818 127392
rect 496874 127336 496879 127392
rect 494316 127334 496879 127336
rect 496813 127331 496879 127334
rect 252277 127258 252343 127261
rect 248952 127256 252343 127258
rect 248952 127200 252282 127256
rect 252338 127200 252343 127256
rect 248952 127198 252343 127200
rect 252277 127195 252343 127198
rect 307661 127258 307727 127261
rect 307661 127256 310040 127258
rect 307661 127200 307666 127256
rect 307722 127200 310040 127256
rect 307661 127198 310040 127200
rect 307661 127195 307727 127198
rect 324405 127122 324471 127125
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 213913 127062 217242 127064
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 166276 127060 166282 127062
rect 213913 127059 213979 127062
rect 324405 127059 324471 127062
rect 306557 126850 306623 126853
rect 306557 126848 310040 126850
rect 306557 126792 306562 126848
rect 306618 126792 310040 126848
rect 306557 126790 310040 126792
rect 306557 126787 306623 126790
rect 252461 126714 252527 126717
rect 248952 126712 252527 126714
rect 65149 126306 65215 126309
rect 68142 126306 68816 126312
rect 65149 126304 68816 126306
rect 65149 126248 65154 126304
rect 65210 126252 68816 126304
rect 65210 126248 68202 126252
rect 65149 126246 68202 126248
rect 65149 126243 65215 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 248952 126656 252466 126712
rect 252522 126656 252527 126712
rect 248952 126654 252527 126656
rect 252461 126651 252527 126654
rect 307569 126442 307635 126445
rect 307569 126440 310040 126442
rect 307569 126384 307574 126440
rect 307630 126384 310040 126440
rect 307569 126382 310040 126384
rect 307569 126379 307635 126382
rect 252185 126306 252251 126309
rect 496813 126306 496879 126309
rect 248952 126304 252251 126306
rect 248952 126248 252190 126304
rect 252246 126248 252251 126304
rect 494316 126304 496879 126306
rect 248952 126246 252251 126248
rect 252185 126243 252251 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 307661 125898 307727 125901
rect 307661 125896 310040 125898
rect 307661 125840 307666 125896
rect 307722 125840 310040 125896
rect 307661 125838 310040 125840
rect 307661 125835 307727 125838
rect 251909 125762 251975 125765
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 248952 125760 251975 125762
rect 248952 125704 251914 125760
rect 251970 125704 251975 125760
rect 248952 125702 251975 125704
rect 213913 125699 213979 125702
rect 251909 125699 251975 125702
rect 321878 125626 321938 126276
rect 494316 126248 496818 126304
rect 496874 126248 496879 126304
rect 494316 126246 496879 126248
rect 496813 126243 496879 126246
rect 419441 126170 419507 126173
rect 419441 126168 420164 126170
rect 419441 126112 419446 126168
rect 419502 126112 420164 126168
rect 419441 126110 420164 126112
rect 419441 126107 419507 126110
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 328494 125626 328500 125628
rect 321878 125566 328500 125626
rect 328494 125564 328500 125566
rect 328564 125564 328570 125628
rect 307293 125490 307359 125493
rect 324313 125490 324379 125493
rect 307293 125488 310040 125490
rect 307293 125432 307298 125488
rect 307354 125432 310040 125488
rect 307293 125430 310040 125432
rect 321908 125488 324379 125490
rect 321908 125432 324318 125488
rect 324374 125432 324379 125488
rect 321908 125430 324379 125432
rect 307293 125427 307359 125430
rect 324313 125427 324379 125430
rect 252369 125354 252435 125357
rect 248952 125352 252435 125354
rect 67449 125218 67515 125221
rect 68142 125218 68816 125224
rect 67449 125216 68816 125218
rect 67449 125160 67454 125216
rect 67510 125164 68816 125216
rect 67510 125160 68202 125164
rect 67449 125158 68202 125160
rect 67449 125155 67515 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 248952 125296 252374 125352
rect 252430 125296 252435 125352
rect 248952 125294 252435 125296
rect 252369 125291 252435 125294
rect 496813 125218 496879 125221
rect 494316 125216 496879 125218
rect 494316 125160 496818 125216
rect 496874 125160 496879 125216
rect 494316 125158 496879 125160
rect 496813 125155 496879 125158
rect 307569 125082 307635 125085
rect 307569 125080 310040 125082
rect 307569 125024 307574 125080
rect 307630 125024 310040 125080
rect 307569 125022 310040 125024
rect 307569 125019 307635 125022
rect 252461 124810 252527 124813
rect 324405 124810 324471 124813
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 248952 124808 252527 124810
rect 248952 124752 252466 124808
rect 252522 124752 252527 124808
rect 248952 124750 252527 124752
rect 321908 124808 324471 124810
rect 321908 124752 324410 124808
rect 324466 124752 324471 124808
rect 321908 124750 324471 124752
rect 214005 124747 214071 124750
rect 252461 124747 252527 124750
rect 324405 124747 324471 124750
rect 307661 124674 307727 124677
rect 307661 124672 310040 124674
rect 213913 124266 213979 124269
rect 217182 124266 217242 124644
rect 307661 124616 307666 124672
rect 307722 124616 310040 124672
rect 307661 124614 310040 124616
rect 307661 124611 307727 124614
rect 419533 124538 419599 124541
rect 419533 124536 420164 124538
rect 419533 124480 419538 124536
rect 419594 124480 420164 124536
rect 419533 124478 420164 124480
rect 419533 124475 419599 124478
rect 252277 124402 252343 124405
rect 248952 124400 252343 124402
rect 248952 124344 252282 124400
rect 252338 124344 252343 124400
rect 248952 124342 252343 124344
rect 252277 124339 252343 124342
rect 213913 124264 217242 124266
rect 213913 124208 213918 124264
rect 213974 124208 217242 124264
rect 213913 124206 217242 124208
rect 307201 124266 307267 124269
rect 307201 124264 310040 124266
rect 307201 124208 307206 124264
rect 307262 124208 310040 124264
rect 307201 124206 310040 124208
rect 213913 124203 213979 124206
rect 307201 124203 307267 124206
rect 496813 124130 496879 124133
rect 494316 124128 496879 124130
rect -960 123572 480 123812
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 494316 124072 496818 124128
rect 496874 124072 496879 124128
rect 494316 124070 496879 124072
rect 496813 124067 496879 124070
rect 252369 123994 252435 123997
rect 324313 123994 324379 123997
rect 248952 123992 252435 123994
rect 248952 123936 252374 123992
rect 252430 123936 252435 123992
rect 248952 123934 252435 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252369 123931 252435 123934
rect 324313 123931 324379 123934
rect 307569 123858 307635 123861
rect 307569 123856 310040 123858
rect 307569 123800 307574 123856
rect 307630 123800 310040 123856
rect 307569 123798 310040 123800
rect 307569 123795 307635 123798
rect 214005 123584 217242 123586
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 66069 123523 66135 123526
rect 214005 123523 214071 123526
rect 252461 123450 252527 123453
rect 308397 123450 308463 123453
rect 248952 123448 252527 123450
rect 213913 122906 213979 122909
rect 217182 122906 217242 123420
rect 248952 123392 252466 123448
rect 252522 123392 252527 123448
rect 248952 123390 252527 123392
rect 252461 123387 252527 123390
rect 258030 123448 308463 123450
rect 258030 123392 308402 123448
rect 308458 123392 308463 123448
rect 258030 123390 308463 123392
rect 251950 123252 251956 123316
rect 252020 123314 252026 123316
rect 258030 123314 258090 123390
rect 308397 123387 308463 123390
rect 309550 123346 310132 123406
rect 252020 123254 258090 123314
rect 305821 123314 305887 123317
rect 309550 123314 309610 123346
rect 305821 123312 309610 123314
rect 305821 123256 305826 123312
rect 305882 123256 309610 123312
rect 305821 123254 309610 123256
rect 252020 123252 252026 123254
rect 305821 123251 305887 123254
rect 324405 123178 324471 123181
rect 321908 123176 324471 123178
rect 321908 123120 324410 123176
rect 324466 123120 324471 123176
rect 321908 123118 324471 123120
rect 324405 123115 324471 123118
rect 251766 123042 251772 123044
rect 248952 122982 251772 123042
rect 251766 122980 251772 122982
rect 251836 122980 251842 123044
rect 307661 123042 307727 123045
rect 307661 123040 310040 123042
rect 307661 122984 307666 123040
rect 307722 122984 310040 123040
rect 307661 122982 310040 122984
rect 307661 122979 307727 122982
rect 496905 122906 496971 122909
rect 213913 122904 217242 122906
rect 213913 122848 213918 122904
rect 213974 122848 217242 122904
rect 213913 122846 217242 122848
rect 494316 122904 496971 122906
rect 494316 122848 496910 122904
rect 496966 122848 496971 122904
rect 494316 122846 496971 122848
rect 213913 122843 213979 122846
rect 496905 122843 496971 122846
rect 416773 122770 416839 122773
rect 416773 122768 420164 122770
rect 67265 122634 67331 122637
rect 68142 122634 68816 122640
rect 67265 122632 68816 122634
rect 67265 122576 67270 122632
rect 67326 122580 68816 122632
rect 67326 122576 68202 122580
rect 67265 122574 68202 122576
rect 67265 122571 67331 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 416773 122712 416778 122768
rect 416834 122712 420164 122768
rect 416773 122710 420164 122712
rect 416773 122707 416839 122710
rect 252461 122498 252527 122501
rect 248952 122496 252527 122498
rect 248952 122440 252466 122496
rect 252522 122440 252527 122496
rect 248952 122438 252527 122440
rect 252461 122435 252527 122438
rect 307569 122498 307635 122501
rect 324313 122498 324379 122501
rect 307569 122496 310040 122498
rect 307569 122440 307574 122496
rect 307630 122440 310040 122496
rect 307569 122438 310040 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307569 122435 307635 122438
rect 324313 122435 324379 122438
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 214005 122163 214071 122166
rect 252369 122090 252435 122093
rect 248952 122088 252435 122090
rect 213913 121818 213979 121821
rect 217182 121818 217242 122060
rect 248952 122032 252374 122088
rect 252430 122032 252435 122088
rect 248952 122030 252435 122032
rect 252369 122027 252435 122030
rect 307017 122090 307083 122093
rect 307017 122088 310040 122090
rect 307017 122032 307022 122088
rect 307078 122032 310040 122088
rect 307017 122030 310040 122032
rect 307017 122027 307083 122030
rect 496813 121818 496879 121821
rect 213913 121816 217242 121818
rect 213913 121760 213918 121816
rect 213974 121760 217242 121816
rect 213913 121758 217242 121760
rect 494316 121816 496879 121818
rect 494316 121760 496818 121816
rect 496874 121760 496879 121816
rect 494316 121758 496879 121760
rect 213913 121755 213979 121758
rect 496813 121755 496879 121758
rect 307661 121682 307727 121685
rect 324405 121682 324471 121685
rect 307661 121680 310040 121682
rect 307661 121624 307666 121680
rect 307722 121624 310040 121680
rect 307661 121622 310040 121624
rect 321908 121680 324471 121682
rect 321908 121624 324410 121680
rect 324466 121624 324471 121680
rect 321908 121622 324471 121624
rect 307661 121619 307727 121622
rect 324405 121619 324471 121622
rect 252277 121546 252343 121549
rect 248952 121544 252343 121546
rect 248952 121488 252282 121544
rect 252338 121488 252343 121544
rect 248952 121486 252343 121488
rect 252277 121483 252343 121486
rect 67633 120866 67699 120869
rect 68142 120866 68816 120872
rect 67633 120864 68816 120866
rect 67633 120808 67638 120864
rect 67694 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 307477 121274 307543 121277
rect 307477 121272 310040 121274
rect 307477 121216 307482 121272
rect 307538 121216 310040 121272
rect 307477 121214 310040 121216
rect 307477 121211 307543 121214
rect 252277 121138 252343 121141
rect 248952 121136 252343 121138
rect 248952 121080 252282 121136
rect 252338 121080 252343 121136
rect 248952 121078 252343 121080
rect 252277 121075 252343 121078
rect 416773 121138 416839 121141
rect 416773 121136 420164 121138
rect 416773 121080 416778 121136
rect 416834 121080 420164 121136
rect 416773 121078 420164 121080
rect 416773 121075 416839 121078
rect 214005 120864 217242 120866
rect 67694 120808 68202 120812
rect 67633 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310040 120866
rect 307569 120808 307574 120864
rect 307630 120808 310040 120864
rect 307569 120806 310040 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 67633 120803 67699 120806
rect 214005 120803 214071 120806
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 498377 120730 498443 120733
rect 494316 120728 498443 120730
rect 213913 120458 213979 120461
rect 217182 120458 217242 120700
rect 494316 120672 498382 120728
rect 498438 120672 498443 120728
rect 494316 120670 498443 120672
rect 498377 120667 498443 120670
rect 252461 120594 252527 120597
rect 248952 120592 252527 120594
rect 248952 120536 252466 120592
rect 252522 120536 252527 120592
rect 248952 120534 252527 120536
rect 252461 120531 252527 120534
rect 213913 120456 217242 120458
rect 213913 120400 213918 120456
rect 213974 120400 217242 120456
rect 213913 120398 217242 120400
rect 307661 120458 307727 120461
rect 307661 120456 310040 120458
rect 307661 120400 307666 120456
rect 307722 120400 310040 120456
rect 307661 120398 310040 120400
rect 213913 120395 213979 120398
rect 307661 120395 307727 120398
rect 252369 120186 252435 120189
rect 324405 120186 324471 120189
rect 248952 120184 252435 120186
rect 248952 120128 252374 120184
rect 252430 120128 252435 120184
rect 248952 120126 252435 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 252369 120123 252435 120126
rect 324405 120123 324471 120126
rect 307569 120050 307635 120053
rect 307569 120048 310040 120050
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 307569 119992 307574 120048
rect 307630 119992 310040 120048
rect 307569 119990 310040 119992
rect 307569 119987 307635 119990
rect 252461 119642 252527 119645
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 248952 119640 252527 119642
rect 248952 119584 252466 119640
rect 252522 119584 252527 119640
rect 248952 119582 252527 119584
rect 214005 119579 214071 119582
rect 252461 119579 252527 119582
rect 307661 119642 307727 119645
rect 496813 119642 496879 119645
rect 307661 119640 310040 119642
rect 307661 119584 307666 119640
rect 307722 119584 310040 119640
rect 307661 119582 310040 119584
rect 494316 119640 496879 119642
rect 494316 119584 496818 119640
rect 496874 119584 496879 119640
rect 494316 119582 496879 119584
rect 307661 119579 307727 119582
rect 496813 119579 496879 119582
rect 213453 119098 213519 119101
rect 217182 119098 217242 119476
rect 254945 119370 255011 119373
rect 306966 119370 306972 119372
rect 254945 119368 306972 119370
rect 254945 119312 254950 119368
rect 255006 119312 306972 119368
rect 254945 119310 306972 119312
rect 254945 119307 255011 119310
rect 306966 119308 306972 119310
rect 307036 119308 307042 119372
rect 325877 119370 325943 119373
rect 321908 119368 325943 119370
rect 321908 119312 325882 119368
rect 325938 119312 325943 119368
rect 321908 119310 325943 119312
rect 325877 119307 325943 119310
rect 417417 119370 417483 119373
rect 417417 119368 420164 119370
rect 417417 119312 417422 119368
rect 417478 119312 420164 119368
rect 417417 119310 420164 119312
rect 417417 119307 417483 119310
rect 252369 119234 252435 119237
rect 248952 119232 252435 119234
rect 248952 119176 252374 119232
rect 252430 119176 252435 119232
rect 248952 119174 252435 119176
rect 252369 119171 252435 119174
rect 213453 119096 217242 119098
rect 213453 119040 213458 119096
rect 213514 119040 217242 119096
rect 213453 119038 217242 119040
rect 307293 119098 307359 119101
rect 307293 119096 310040 119098
rect 307293 119040 307298 119096
rect 307354 119040 310040 119096
rect 307293 119038 310040 119040
rect 213453 119035 213519 119038
rect 307293 119035 307359 119038
rect 213913 118962 213979 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 252001 118826 252067 118829
rect 248952 118824 252067 118826
rect 248952 118768 252006 118824
rect 252062 118768 252067 118824
rect 248952 118766 252067 118768
rect 252001 118763 252067 118766
rect 307477 118690 307543 118693
rect 307477 118688 310040 118690
rect 307477 118632 307482 118688
rect 307538 118632 310040 118688
rect 307477 118630 310040 118632
rect 307477 118627 307543 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 496813 118418 496879 118421
rect 494316 118416 496879 118418
rect 494316 118360 496818 118416
rect 496874 118360 496879 118416
rect 494316 118358 496879 118360
rect 496813 118355 496879 118358
rect 252461 118282 252527 118285
rect 248952 118280 252527 118282
rect 248952 118224 252466 118280
rect 252522 118224 252527 118280
rect 248952 118222 252527 118224
rect 252461 118219 252527 118222
rect 307569 118282 307635 118285
rect 307569 118280 310040 118282
rect 307569 118224 307574 118280
rect 307630 118224 310040 118280
rect 307569 118222 310040 118224
rect 307569 118219 307635 118222
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 252369 117874 252435 117877
rect 248952 117872 252435 117874
rect 248952 117816 252374 117872
rect 252430 117816 252435 117872
rect 248952 117814 252435 117816
rect 252369 117811 252435 117814
rect 306741 117874 306807 117877
rect 324405 117874 324471 117877
rect 306741 117872 310040 117874
rect 306741 117816 306746 117872
rect 306802 117816 310040 117872
rect 306741 117814 310040 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 306741 117811 306807 117814
rect 324405 117811 324471 117814
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 214005 117539 214071 117542
rect 307661 117466 307727 117469
rect 307661 117464 310040 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 307661 117408 307666 117464
rect 307722 117408 310040 117464
rect 307661 117406 310040 117408
rect 307661 117403 307727 117406
rect 251817 117330 251883 117333
rect 248952 117328 251883 117330
rect 248952 117272 251822 117328
rect 251878 117272 251883 117328
rect 248952 117270 251883 117272
rect 251817 117267 251883 117270
rect 334566 117268 334572 117332
rect 334636 117330 334642 117332
rect 420134 117330 420194 117708
rect 496813 117330 496879 117333
rect 334636 117270 420194 117330
rect 494316 117328 496879 117330
rect 494316 117272 496818 117328
rect 496874 117272 496879 117328
rect 494316 117270 496879 117272
rect 334636 117268 334642 117270
rect 496813 117267 496879 117270
rect 216814 117134 217426 117194
rect 307477 117058 307543 117061
rect 324313 117058 324379 117061
rect 307477 117056 310040 117058
rect 307477 117000 307482 117056
rect 307538 117000 310040 117056
rect 307477 116998 310040 117000
rect 321908 117056 324379 117058
rect 321908 117000 324318 117056
rect 324374 117000 324379 117056
rect 321908 116998 324379 117000
rect 307477 116995 307543 116998
rect 324313 116995 324379 116998
rect 252461 116922 252527 116925
rect 248952 116920 252527 116922
rect 248952 116864 252466 116920
rect 252522 116864 252527 116920
rect 248952 116862 252527 116864
rect 252461 116859 252527 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 307569 116650 307635 116653
rect 307569 116648 310040 116650
rect 307569 116592 307574 116648
rect 307630 116592 310040 116648
rect 307569 116590 310040 116592
rect 307569 116587 307635 116590
rect 252277 116378 252343 116381
rect 324405 116378 324471 116381
rect 248952 116376 252343 116378
rect 248952 116320 252282 116376
rect 252338 116320 252343 116376
rect 248952 116318 252343 116320
rect 321908 116376 324471 116378
rect 321908 116320 324410 116376
rect 324466 116320 324471 116376
rect 321908 116318 324471 116320
rect 252277 116315 252343 116318
rect 324405 116315 324471 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 307661 116242 307727 116245
rect 496905 116242 496971 116245
rect 307661 116240 310040 116242
rect 307661 116184 307666 116240
rect 307722 116184 310040 116240
rect 307661 116182 310040 116184
rect 494316 116240 496971 116242
rect 494316 116184 496910 116240
rect 496966 116184 496971 116240
rect 494316 116182 496971 116184
rect 214005 116179 214071 116182
rect 307661 116179 307727 116182
rect 496905 116179 496971 116182
rect 416773 116106 416839 116109
rect 416773 116104 420164 116106
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 416773 116048 416778 116104
rect 416834 116048 420164 116104
rect 416773 116046 420164 116048
rect 416773 116043 416839 116046
rect 252369 115970 252435 115973
rect 248952 115968 252435 115970
rect 248952 115912 252374 115968
rect 252430 115912 252435 115968
rect 248952 115910 252435 115912
rect 252369 115907 252435 115910
rect 216814 115774 217426 115834
rect 307569 115698 307635 115701
rect 307569 115696 310040 115698
rect 307569 115640 307574 115696
rect 307630 115640 310040 115696
rect 307569 115638 310040 115640
rect 307569 115635 307635 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 252461 115426 252527 115429
rect 248952 115424 252527 115426
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 248952 115368 252466 115424
rect 252522 115368 252527 115424
rect 248952 115366 252527 115368
rect 252461 115363 252527 115366
rect 307661 115290 307727 115293
rect 307661 115288 310040 115290
rect 307661 115232 307666 115288
rect 307722 115232 310040 115288
rect 307661 115230 310040 115232
rect 307661 115227 307727 115230
rect 498285 115154 498351 115157
rect 494316 115152 498351 115154
rect 494316 115096 498290 115152
rect 498346 115096 498351 115152
rect 494316 115094 498351 115096
rect 498285 115091 498351 115094
rect 252369 115018 252435 115021
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 248952 115016 252435 115018
rect 248952 114960 252374 115016
rect 252430 114960 252435 115016
rect 248952 114958 252435 114960
rect 214005 114955 214071 114958
rect 252369 114955 252435 114958
rect 213913 114610 213979 114613
rect 217182 114610 217242 114852
rect 249558 114820 249564 114884
rect 249628 114882 249634 114884
rect 249628 114822 310040 114882
rect 249628 114820 249634 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 213913 114608 217242 114610
rect 213913 114552 213918 114608
rect 213974 114552 217242 114608
rect 213913 114550 217242 114552
rect 213913 114547 213979 114550
rect 252461 114474 252527 114477
rect 248952 114472 252527 114474
rect 248952 114416 252466 114472
rect 252522 114416 252527 114472
rect 248952 114414 252527 114416
rect 252461 114411 252527 114414
rect 309550 114370 310132 114430
rect 302734 114276 302740 114340
rect 302804 114338 302810 114340
rect 309550 114338 309610 114370
rect 302804 114278 309610 114338
rect 302804 114276 302810 114278
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 252369 114066 252435 114069
rect 248952 114064 252435 114066
rect 248952 114008 252374 114064
rect 252430 114008 252435 114064
rect 248952 114006 252435 114008
rect 252369 114003 252435 114006
rect 307569 114066 307635 114069
rect 324313 114066 324379 114069
rect 307569 114064 310040 114066
rect 307569 114008 307574 114064
rect 307630 114008 310040 114064
rect 307569 114006 310040 114008
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307569 114003 307635 114006
rect 324313 114003 324379 114006
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 307661 113658 307727 113661
rect 307661 113656 310040 113658
rect 307661 113600 307666 113656
rect 307722 113600 310040 113656
rect 307661 113598 310040 113600
rect 214005 113595 214071 113598
rect 307661 113595 307727 113598
rect 252277 113522 252343 113525
rect 248952 113520 252343 113522
rect 213913 113250 213979 113253
rect 217366 113250 217426 113492
rect 248952 113464 252282 113520
rect 252338 113464 252343 113520
rect 248952 113462 252343 113464
rect 252277 113459 252343 113462
rect 213913 113248 217426 113250
rect 213913 113192 213918 113248
rect 213974 113192 217426 113248
rect 213913 113190 217426 113192
rect 306741 113250 306807 113253
rect 324405 113250 324471 113253
rect 306741 113248 310040 113250
rect 306741 113192 306746 113248
rect 306802 113192 310040 113248
rect 306741 113190 310040 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 213913 113187 213979 113190
rect 306741 113187 306807 113190
rect 324405 113187 324471 113190
rect 345606 113188 345612 113252
rect 345676 113250 345682 113252
rect 420134 113250 420194 114308
rect 495433 113930 495499 113933
rect 494316 113928 495499 113930
rect 494316 113872 495438 113928
rect 495494 113872 495499 113928
rect 494316 113870 495499 113872
rect 495433 113867 495499 113870
rect 345676 113190 420194 113250
rect 345676 113188 345682 113190
rect 252461 113114 252527 113117
rect 248952 113112 252527 113114
rect 248952 113056 252466 113112
rect 252522 113056 252527 113112
rect 248952 113054 252527 113056
rect 252461 113051 252527 113054
rect 496905 112842 496971 112845
rect 494316 112840 496971 112842
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 494316 112784 496910 112840
rect 496966 112784 496971 112840
rect 494316 112782 496971 112784
rect 496905 112779 496971 112782
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 252461 112706 252527 112709
rect 248952 112704 252527 112706
rect 248952 112648 252466 112704
rect 252522 112648 252527 112704
rect 248952 112646 252527 112648
rect 252461 112643 252527 112646
rect 307569 112706 307635 112709
rect 416773 112706 416839 112709
rect 307569 112704 310040 112706
rect 307569 112648 307574 112704
rect 307630 112648 310040 112704
rect 307569 112646 310040 112648
rect 416773 112704 420164 112706
rect 416773 112648 416778 112704
rect 416834 112648 420164 112704
rect 583520 112692 584960 112782
rect 416773 112646 420164 112648
rect 307569 112643 307635 112646
rect 416773 112643 416839 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 214005 112235 214071 112238
rect 309550 112194 310132 112254
rect 252369 112162 252435 112165
rect 248952 112160 252435 112162
rect 213913 111890 213979 111893
rect 217366 111890 217426 112132
rect 248952 112104 252374 112160
rect 252430 112104 252435 112160
rect 248952 112102 252435 112104
rect 252369 112099 252435 112102
rect 305913 112026 305979 112029
rect 309550 112026 309610 112194
rect 305913 112024 309610 112026
rect 305913 111968 305918 112024
rect 305974 111968 309610 112024
rect 305913 111966 309610 111968
rect 305913 111963 305979 111966
rect 213913 111888 217426 111890
rect 213913 111832 213918 111888
rect 213974 111832 217426 111888
rect 213913 111830 217426 111832
rect 307661 111890 307727 111893
rect 307661 111888 310040 111890
rect 307661 111832 307666 111888
rect 307722 111832 310040 111888
rect 307661 111830 310040 111832
rect 213913 111827 213979 111830
rect 307661 111827 307727 111830
rect 167913 111754 167979 111757
rect 252461 111754 252527 111757
rect 323025 111754 323091 111757
rect 496813 111754 496879 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 248952 111752 252527 111754
rect 248952 111696 252466 111752
rect 252522 111696 252527 111752
rect 248952 111694 252527 111696
rect 321908 111752 323091 111754
rect 321908 111696 323030 111752
rect 323086 111696 323091 111752
rect 321908 111694 323091 111696
rect 494316 111752 496879 111754
rect 494316 111696 496818 111752
rect 496874 111696 496879 111752
rect 494316 111694 496879 111696
rect 167913 111691 167979 111694
rect 252461 111691 252527 111694
rect 323025 111691 323091 111694
rect 496813 111691 496879 111694
rect 307477 111482 307543 111485
rect 307477 111480 310040 111482
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 307477 111424 307482 111480
rect 307538 111424 310040 111480
rect 307477 111422 310040 111424
rect 307477 111419 307543 111422
rect 252369 111210 252435 111213
rect 248952 111208 252435 111210
rect 248952 111152 252374 111208
rect 252430 111152 252435 111208
rect 248952 111150 252435 111152
rect 252369 111147 252435 111150
rect 307569 111074 307635 111077
rect 307569 111072 310040 111074
rect 307569 111016 307574 111072
rect 307630 111016 310040 111072
rect 307569 111014 310040 111016
rect 307569 111011 307635 111014
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 416773 110938 416839 110941
rect 416773 110936 420164 110938
rect 214005 110878 217242 110880
rect 214005 110875 214071 110878
rect 252461 110802 252527 110805
rect 248952 110800 252527 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217366 110530 217426 110772
rect 248952 110744 252466 110800
rect 252522 110744 252527 110800
rect 248952 110742 252527 110744
rect 252461 110739 252527 110742
rect 307661 110666 307727 110669
rect 307661 110664 310040 110666
rect 307661 110608 307666 110664
rect 307722 110608 310040 110664
rect 307661 110606 310040 110608
rect 307661 110603 307727 110606
rect 321878 110533 321938 110908
rect 416773 110880 416778 110936
rect 416834 110880 420164 110936
rect 416773 110878 420164 110880
rect 416773 110875 416839 110878
rect 213913 110528 217426 110530
rect 213913 110472 213918 110528
rect 213974 110472 217426 110528
rect 213913 110470 217426 110472
rect 321829 110528 321938 110533
rect 321829 110472 321834 110528
rect 321890 110472 321938 110528
rect 321829 110470 321938 110472
rect 494286 110530 494346 110636
rect 502374 110530 502380 110532
rect 494286 110470 502380 110530
rect 213913 110467 213979 110470
rect 321829 110467 321895 110470
rect 502374 110468 502380 110470
rect 502444 110468 502450 110532
rect 252461 110258 252527 110261
rect 248952 110256 252527 110258
rect 168005 110122 168071 110125
rect 164694 110120 168071 110122
rect 164694 110064 168010 110120
rect 168066 110064 168071 110120
rect 164694 110062 168071 110064
rect 168005 110059 168071 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 248952 110200 252466 110256
rect 252522 110200 252527 110256
rect 248952 110198 252527 110200
rect 252461 110195 252527 110198
rect 307569 110258 307635 110261
rect 307569 110256 310040 110258
rect 307569 110200 307574 110256
rect 307630 110200 310040 110256
rect 307569 110198 310040 110200
rect 307569 110195 307635 110198
rect 252369 109850 252435 109853
rect 248952 109848 252435 109850
rect 248952 109792 252374 109848
rect 252430 109792 252435 109848
rect 248952 109790 252435 109792
rect 252369 109787 252435 109790
rect 306741 109850 306807 109853
rect 306741 109848 310040 109850
rect 306741 109792 306746 109848
rect 306802 109792 310040 109848
rect 306741 109790 310040 109792
rect 306741 109787 306807 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 214005 109651 214071 109654
rect 321510 109580 321570 110092
rect 213913 109170 213979 109173
rect 217182 109170 217242 109548
rect 321502 109516 321508 109580
rect 321572 109516 321578 109580
rect 324313 109442 324379 109445
rect 496813 109442 496879 109445
rect 321908 109440 324379 109442
rect 321908 109384 324318 109440
rect 324374 109384 324379 109440
rect 321908 109382 324379 109384
rect 494316 109440 496879 109442
rect 494316 109384 496818 109440
rect 496874 109384 496879 109440
rect 494316 109382 496879 109384
rect 324313 109379 324379 109382
rect 496813 109379 496879 109382
rect 252277 109306 252343 109309
rect 248952 109304 252343 109306
rect 248952 109248 252282 109304
rect 252338 109248 252343 109304
rect 248952 109246 252343 109248
rect 252277 109243 252343 109246
rect 307661 109306 307727 109309
rect 416773 109306 416839 109309
rect 307661 109304 310040 109306
rect 307661 109248 307666 109304
rect 307722 109248 310040 109304
rect 307661 109246 310040 109248
rect 416773 109304 420164 109306
rect 416773 109248 416778 109304
rect 416834 109248 420164 109304
rect 416773 109246 420164 109248
rect 307661 109243 307727 109246
rect 416773 109243 416839 109246
rect 213913 109168 217242 109170
rect 213913 109112 213918 109168
rect 213974 109112 217242 109168
rect 213913 109110 217242 109112
rect 213913 109107 213979 109110
rect 252461 108898 252527 108901
rect 248952 108896 252527 108898
rect 169017 108762 169083 108765
rect 164694 108760 169083 108762
rect 164694 108704 169022 108760
rect 169078 108704 169083 108760
rect 164694 108702 169083 108704
rect 169017 108699 169083 108702
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 248952 108840 252466 108896
rect 252522 108840 252527 108896
rect 248952 108838 252527 108840
rect 252461 108835 252527 108838
rect 306925 108898 306991 108901
rect 306925 108896 310040 108898
rect 306925 108840 306930 108896
rect 306986 108840 310040 108896
rect 306925 108838 310040 108840
rect 306925 108835 306991 108838
rect 324681 108626 324747 108629
rect 321908 108624 324747 108626
rect 321908 108568 324686 108624
rect 324742 108568 324747 108624
rect 321908 108566 324747 108568
rect 324681 108563 324747 108566
rect 307569 108490 307635 108493
rect 307569 108488 310040 108490
rect 307569 108432 307574 108488
rect 307630 108432 310040 108488
rect 307569 108430 310040 108432
rect 307569 108427 307635 108430
rect 252277 108354 252343 108357
rect 497089 108354 497155 108357
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 248952 108352 252343 108354
rect 248952 108296 252282 108352
rect 252338 108296 252343 108352
rect 248952 108294 252343 108296
rect 494316 108352 497155 108354
rect 494316 108296 497094 108352
rect 497150 108296 497155 108352
rect 494316 108294 497155 108296
rect 214005 108291 214071 108294
rect 252277 108291 252343 108294
rect 497089 108291 497155 108294
rect 213913 107810 213979 107813
rect 217182 107810 217242 108188
rect 307661 108082 307727 108085
rect 307661 108080 310040 108082
rect 307661 108024 307666 108080
rect 307722 108024 310040 108080
rect 307661 108022 310040 108024
rect 307661 108019 307727 108022
rect 252369 107946 252435 107949
rect 248952 107944 252435 107946
rect 248952 107888 252374 107944
rect 252430 107888 252435 107944
rect 248952 107886 252435 107888
rect 252369 107883 252435 107886
rect 213913 107808 217242 107810
rect 213913 107752 213918 107808
rect 213974 107752 217242 107808
rect 213913 107750 217242 107752
rect 305729 107810 305795 107813
rect 307569 107810 307635 107813
rect 324313 107810 324379 107813
rect 305729 107808 307635 107810
rect 305729 107752 305734 107808
rect 305790 107752 307574 107808
rect 307630 107752 307635 107808
rect 305729 107750 307635 107752
rect 321908 107808 324379 107810
rect 321908 107752 324318 107808
rect 324374 107752 324379 107808
rect 321908 107750 324379 107752
rect 213913 107747 213979 107750
rect 305729 107747 305795 107750
rect 307569 107747 307635 107750
rect 324313 107747 324379 107750
rect 307477 107674 307543 107677
rect 307477 107672 310040 107674
rect 307477 107616 307482 107672
rect 307538 107616 310040 107672
rect 307477 107614 310040 107616
rect 307477 107611 307543 107614
rect 252461 107538 252527 107541
rect 248952 107536 252527 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 248952 107480 252466 107536
rect 252522 107480 252527 107536
rect 248952 107478 252527 107480
rect 252461 107475 252527 107478
rect 416773 107538 416839 107541
rect 416773 107536 420164 107538
rect 416773 107480 416778 107536
rect 416834 107480 420164 107536
rect 416773 107478 420164 107480
rect 416773 107475 416839 107478
rect 307569 107266 307635 107269
rect 496997 107266 497063 107269
rect 307569 107264 310040 107266
rect 307569 107208 307574 107264
rect 307630 107208 310040 107264
rect 307569 107206 310040 107208
rect 494316 107264 497063 107266
rect 494316 107208 497002 107264
rect 497058 107208 497063 107264
rect 494316 107206 497063 107208
rect 307569 107203 307635 107206
rect 496997 107203 497063 107206
rect 324313 107130 324379 107133
rect 321908 107128 324379 107130
rect 321908 107072 324318 107128
rect 324374 107072 324379 107128
rect 321908 107070 324379 107072
rect 324313 107067 324379 107070
rect 252369 106994 252435 106997
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 248952 106992 252435 106994
rect 248952 106936 252374 106992
rect 252430 106936 252435 106992
rect 248952 106934 252435 106936
rect 214005 106931 214071 106934
rect 252369 106931 252435 106934
rect 307477 106858 307543 106861
rect 307477 106856 310040 106858
rect 213913 106450 213979 106453
rect 217182 106450 217242 106828
rect 307477 106800 307482 106856
rect 307538 106800 310040 106856
rect 307477 106798 310040 106800
rect 307477 106795 307543 106798
rect 252093 106586 252159 106589
rect 248952 106584 252159 106586
rect 248952 106528 252098 106584
rect 252154 106528 252159 106584
rect 248952 106526 252159 106528
rect 252093 106523 252159 106526
rect 213913 106448 217242 106450
rect 213913 106392 213918 106448
rect 213974 106392 217242 106448
rect 213913 106390 217242 106392
rect 307661 106450 307727 106453
rect 307661 106448 310040 106450
rect 307661 106392 307666 106448
rect 307722 106392 310040 106448
rect 307661 106390 310040 106392
rect 213913 106387 213979 106390
rect 307661 106387 307727 106390
rect 323117 106314 323183 106317
rect 321908 106312 323183 106314
rect 321908 106256 323122 106312
rect 323178 106256 323183 106312
rect 321908 106254 323183 106256
rect 323117 106251 323183 106254
rect 496905 106178 496971 106181
rect 494316 106176 496971 106178
rect 213913 105770 213979 105773
rect 217182 105770 217242 106148
rect 494316 106120 496910 106176
rect 496966 106120 496971 106176
rect 494316 106118 496971 106120
rect 496905 106115 496971 106118
rect 252461 106042 252527 106045
rect 248952 106040 252527 106042
rect 248952 105984 252466 106040
rect 252522 105984 252527 106040
rect 248952 105982 252527 105984
rect 252461 105979 252527 105982
rect 307477 105906 307543 105909
rect 416773 105906 416839 105909
rect 307477 105904 310040 105906
rect 307477 105848 307482 105904
rect 307538 105848 310040 105904
rect 307477 105846 310040 105848
rect 416773 105904 420164 105906
rect 416773 105848 416778 105904
rect 416834 105848 420164 105904
rect 416773 105846 420164 105848
rect 307477 105843 307543 105846
rect 416773 105843 416839 105846
rect 213913 105768 217242 105770
rect 213913 105712 213918 105768
rect 213974 105712 217242 105768
rect 213913 105710 217242 105712
rect 213913 105707 213979 105710
rect 251817 105634 251883 105637
rect 248952 105632 251883 105634
rect 216121 105362 216187 105365
rect 217182 105362 217242 105604
rect 248952 105576 251822 105632
rect 251878 105576 251883 105632
rect 248952 105574 251883 105576
rect 251817 105571 251883 105574
rect 307569 105498 307635 105501
rect 323209 105498 323275 105501
rect 307569 105496 310040 105498
rect 307569 105440 307574 105496
rect 307630 105440 310040 105496
rect 307569 105438 310040 105440
rect 321908 105496 323275 105498
rect 321908 105440 323214 105496
rect 323270 105440 323275 105496
rect 321908 105438 323275 105440
rect 307569 105435 307635 105438
rect 323209 105435 323275 105438
rect 216121 105360 217242 105362
rect 216121 105304 216126 105360
rect 216182 105304 217242 105360
rect 216121 105302 217242 105304
rect 216121 105299 216187 105302
rect 214598 105164 214604 105228
rect 214668 105226 214674 105228
rect 214668 105166 217426 105226
rect 214668 105164 214674 105166
rect 217366 104924 217426 105166
rect 252001 105090 252067 105093
rect 248952 105088 252067 105090
rect 248952 105032 252006 105088
rect 252062 105032 252067 105088
rect 248952 105030 252067 105032
rect 252001 105027 252067 105030
rect 307661 105090 307727 105093
rect 307661 105088 310040 105090
rect 307661 105032 307666 105088
rect 307722 105032 310040 105088
rect 307661 105030 310040 105032
rect 307661 105027 307727 105030
rect 496813 104954 496879 104957
rect 494316 104952 496879 104954
rect 494316 104896 496818 104952
rect 496874 104896 496879 104952
rect 494316 104894 496879 104896
rect 496813 104891 496879 104894
rect 324405 104818 324471 104821
rect 321908 104816 324471 104818
rect 321908 104760 324410 104816
rect 324466 104760 324471 104816
rect 321908 104758 324471 104760
rect 324405 104755 324471 104758
rect 252461 104682 252527 104685
rect 248952 104680 252527 104682
rect 248952 104624 252466 104680
rect 252522 104624 252527 104680
rect 248952 104622 252527 104624
rect 252461 104619 252527 104622
rect 307569 104682 307635 104685
rect 307569 104680 310040 104682
rect 307569 104624 307574 104680
rect 307630 104624 310040 104680
rect 307569 104622 310040 104624
rect 307569 104619 307635 104622
rect 306741 104274 306807 104277
rect 306741 104272 310040 104274
rect 213913 103730 213979 103733
rect 217182 103730 217242 104244
rect 306741 104216 306746 104272
rect 306802 104216 310040 104272
rect 306741 104214 310040 104216
rect 306741 104211 306807 104214
rect 252369 104138 252435 104141
rect 248952 104136 252435 104138
rect 248952 104080 252374 104136
rect 252430 104080 252435 104136
rect 248952 104078 252435 104080
rect 252369 104075 252435 104078
rect 416773 104138 416839 104141
rect 416773 104136 420164 104138
rect 416773 104080 416778 104136
rect 416834 104080 420164 104136
rect 416773 104078 420164 104080
rect 416773 104075 416839 104078
rect 325601 104002 325667 104005
rect 321908 104000 325667 104002
rect 321908 103944 325606 104000
rect 325662 103944 325667 104000
rect 321908 103942 325667 103944
rect 325601 103939 325667 103942
rect 307661 103866 307727 103869
rect 307661 103864 310040 103866
rect 307661 103808 307666 103864
rect 307722 103808 310040 103864
rect 307661 103806 310040 103808
rect 307661 103803 307727 103806
rect 494286 103733 494346 103836
rect 252277 103730 252343 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 248952 103728 252343 103730
rect 248952 103672 252282 103728
rect 252338 103672 252343 103728
rect 248952 103670 252343 103672
rect 494286 103728 494395 103733
rect 494286 103672 494334 103728
rect 494390 103672 494395 103728
rect 494286 103670 494395 103672
rect 213913 103667 213979 103670
rect 252277 103667 252343 103670
rect 494329 103667 494395 103670
rect 214414 103532 214420 103596
rect 214484 103594 214490 103596
rect 214484 103534 217058 103594
rect 214484 103532 214490 103534
rect 216998 103530 217058 103534
rect 217182 103530 217242 103564
rect 216998 103470 217242 103530
rect 307569 103458 307635 103461
rect 307569 103456 310040 103458
rect 307569 103400 307574 103456
rect 307630 103400 310040 103456
rect 307569 103398 310040 103400
rect 307569 103395 307635 103398
rect 252461 103186 252527 103189
rect 248952 103184 252527 103186
rect 248952 103128 252466 103184
rect 252522 103128 252527 103184
rect 248952 103126 252527 103128
rect 252461 103123 252527 103126
rect 306741 103050 306807 103053
rect 306741 103048 310040 103050
rect 306741 102992 306746 103048
rect 306802 102992 310040 103048
rect 306741 102990 310040 102992
rect 306741 102987 306807 102990
rect 214005 102506 214071 102509
rect 217182 102506 217242 102884
rect 321694 102781 321754 103156
rect 252369 102778 252435 102781
rect 248952 102776 252435 102778
rect 248952 102720 252374 102776
rect 252430 102720 252435 102776
rect 248952 102718 252435 102720
rect 252369 102715 252435 102718
rect 321645 102776 321754 102781
rect 321645 102720 321650 102776
rect 321706 102720 321754 102776
rect 321645 102718 321754 102720
rect 321645 102715 321711 102718
rect 214005 102504 217242 102506
rect 214005 102448 214010 102504
rect 214066 102448 217242 102504
rect 214005 102446 217242 102448
rect 307661 102506 307727 102509
rect 416773 102506 416839 102509
rect 307661 102504 310040 102506
rect 307661 102448 307666 102504
rect 307722 102448 310040 102504
rect 416773 102504 420164 102506
rect 307661 102446 310040 102448
rect 214005 102443 214071 102446
rect 307661 102443 307727 102446
rect 66069 102370 66135 102373
rect 68142 102370 68816 102376
rect 66069 102368 68816 102370
rect 66069 102312 66074 102368
rect 66130 102316 68816 102368
rect 213913 102370 213979 102373
rect 213913 102368 217242 102370
rect 66130 102312 68202 102316
rect 66069 102310 68202 102312
rect 213913 102312 213918 102368
rect 213974 102312 217242 102368
rect 213913 102310 217242 102312
rect 66069 102307 66135 102310
rect 213913 102307 213979 102310
rect 217182 102204 217242 102310
rect 321694 102237 321754 102476
rect 416773 102448 416778 102504
rect 416834 102448 420164 102504
rect 416773 102446 420164 102448
rect 416773 102443 416839 102446
rect 251173 102234 251239 102237
rect 248952 102232 251239 102234
rect 248952 102176 251178 102232
rect 251234 102176 251239 102232
rect 248952 102174 251239 102176
rect 321694 102232 321803 102237
rect 493918 102236 493978 102748
rect 321694 102176 321742 102232
rect 321798 102176 321803 102232
rect 321694 102174 321803 102176
rect 251173 102171 251239 102174
rect 321737 102171 321803 102174
rect 493910 102172 493916 102236
rect 493980 102172 493986 102236
rect 307569 102098 307635 102101
rect 307569 102096 310040 102098
rect 307569 102040 307574 102096
rect 307630 102040 310040 102096
rect 307569 102038 310040 102040
rect 307569 102035 307635 102038
rect 252461 101826 252527 101829
rect 248952 101824 252527 101826
rect 248952 101768 252466 101824
rect 252522 101768 252527 101824
rect 248952 101766 252527 101768
rect 252461 101763 252527 101766
rect 324497 101690 324563 101693
rect 321908 101688 324563 101690
rect 309550 101586 310132 101646
rect 321908 101632 324502 101688
rect 324558 101632 324563 101688
rect 321908 101630 324563 101632
rect 324497 101627 324563 101630
rect 167729 101418 167795 101421
rect 173934 101418 173940 101420
rect 167729 101416 173940 101418
rect 167729 101360 167734 101416
rect 167790 101360 173940 101416
rect 167729 101358 173940 101360
rect 167729 101355 167795 101358
rect 173934 101356 173940 101358
rect 174004 101356 174010 101420
rect 214005 101282 214071 101285
rect 217182 101282 217242 101524
rect 253197 101418 253263 101421
rect 248952 101416 253263 101418
rect 248952 101360 253202 101416
rect 253258 101360 253263 101416
rect 248952 101358 253263 101360
rect 253197 101355 253263 101358
rect 214005 101280 217242 101282
rect 214005 101224 214010 101280
rect 214066 101224 217242 101280
rect 214005 101222 217242 101224
rect 214005 101219 214071 101222
rect 213913 101146 213979 101149
rect 213913 101144 217242 101146
rect 213913 101088 213918 101144
rect 213974 101088 217242 101144
rect 213913 101086 217242 101088
rect 213913 101083 213979 101086
rect 217182 100980 217242 101086
rect 304206 101084 304212 101148
rect 304276 101146 304282 101148
rect 309550 101146 309610 101586
rect 304276 101086 309610 101146
rect 309734 101178 310132 101238
rect 304276 101084 304282 101086
rect 307661 101010 307727 101013
rect 309734 101010 309794 101178
rect 493961 101146 494027 101149
rect 494102 101146 494162 101660
rect 493961 101144 494162 101146
rect 493961 101088 493966 101144
rect 494022 101088 494162 101144
rect 493961 101086 494162 101088
rect 493961 101083 494027 101086
rect 307661 101008 309794 101010
rect 307661 100952 307666 101008
rect 307722 100952 309794 101008
rect 307661 100950 309794 100952
rect 307661 100947 307727 100950
rect 252277 100874 252343 100877
rect 248952 100872 252343 100874
rect 248952 100816 252282 100872
rect 252338 100816 252343 100872
rect 248952 100814 252343 100816
rect 252277 100811 252343 100814
rect 306925 100874 306991 100877
rect 324589 100874 324655 100877
rect 306925 100872 310040 100874
rect 306925 100816 306930 100872
rect 306986 100816 310040 100872
rect 306925 100814 310040 100816
rect 321908 100872 324655 100874
rect 321908 100816 324594 100872
rect 324650 100816 324655 100872
rect 321908 100814 324655 100816
rect 306925 100811 306991 100814
rect 324589 100811 324655 100814
rect 417509 100874 417575 100877
rect 417509 100872 420164 100874
rect 417509 100816 417514 100872
rect 417570 100816 420164 100872
rect 417509 100814 420164 100816
rect 417509 100811 417575 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 67725 100675 67791 100678
rect 494102 100469 494162 100572
rect 252461 100466 252527 100469
rect 248952 100464 252527 100466
rect 248952 100408 252466 100464
rect 252522 100408 252527 100464
rect 248952 100406 252527 100408
rect 252461 100403 252527 100406
rect 307569 100466 307635 100469
rect 307569 100464 310040 100466
rect 307569 100408 307574 100464
rect 307630 100408 310040 100464
rect 307569 100406 310040 100408
rect 494053 100464 494162 100469
rect 494053 100408 494058 100464
rect 494114 100408 494162 100464
rect 494053 100406 494162 100408
rect 307569 100403 307635 100406
rect 494053 100403 494119 100406
rect 213913 99786 213979 99789
rect 217182 99786 217242 100300
rect 309550 99954 310132 100014
rect 252369 99922 252435 99925
rect 248952 99920 252435 99922
rect 248952 99864 252374 99920
rect 252430 99864 252435 99920
rect 248952 99862 252435 99864
rect 252369 99859 252435 99862
rect 213913 99784 217242 99786
rect 213913 99728 213918 99784
rect 213974 99728 217242 99784
rect 213913 99726 217242 99728
rect 213913 99723 213979 99726
rect 305637 99650 305703 99653
rect 309550 99650 309610 99954
rect 305637 99648 309610 99650
rect 214005 99514 214071 99517
rect 214005 99512 216874 99514
rect 214005 99456 214010 99512
rect 214066 99456 216874 99512
rect 214005 99454 216874 99456
rect 214005 99451 214071 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 305637 99592 305642 99648
rect 305698 99592 309610 99648
rect 321510 99653 321570 100164
rect 321510 99648 321619 99653
rect 305637 99590 309610 99592
rect 305637 99587 305703 99590
rect 309734 99546 310132 99606
rect 321510 99592 321558 99648
rect 321614 99592 321619 99648
rect 321510 99590 321619 99592
rect 321553 99587 321619 99590
rect 252277 99514 252343 99517
rect 248952 99512 252343 99514
rect 248952 99456 252282 99512
rect 252338 99456 252343 99512
rect 248952 99454 252343 99456
rect 252277 99451 252343 99454
rect 307661 99514 307727 99517
rect 309734 99514 309794 99546
rect 307661 99512 309794 99514
rect 307661 99456 307666 99512
rect 307722 99456 309794 99512
rect 307661 99454 309794 99456
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 307661 99451 307727 99454
rect 580165 99451 580231 99454
rect 216814 99318 217426 99378
rect 583520 99364 584960 99454
rect 307661 99106 307727 99109
rect 307661 99104 310040 99106
rect 307661 99048 307666 99104
rect 307722 99048 310040 99104
rect 307661 99046 310040 99048
rect 307661 99043 307727 99046
rect 252461 98970 252527 98973
rect 248952 98968 252527 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 248952 98912 252466 98968
rect 252522 98912 252527 98968
rect 248952 98910 252527 98912
rect 252461 98907 252527 98910
rect 321369 98834 321435 98837
rect 321510 98834 321570 99348
rect 321369 98832 321570 98834
rect 321369 98776 321374 98832
rect 321430 98776 321570 98832
rect 321369 98774 321570 98776
rect 321369 98771 321435 98774
rect 306741 98698 306807 98701
rect 494145 98698 494211 98701
rect 494462 98698 494468 98700
rect 306741 98696 310040 98698
rect 306741 98640 306746 98696
rect 306802 98640 310040 98696
rect 306741 98638 310040 98640
rect 494145 98696 494468 98698
rect 494145 98640 494150 98696
rect 494206 98640 494468 98696
rect 494145 98638 494468 98640
rect 306741 98635 306807 98638
rect 494145 98635 494211 98638
rect 494462 98636 494468 98638
rect 494532 98636 494538 98700
rect 251909 98562 251975 98565
rect 324262 98562 324268 98564
rect 248952 98560 251975 98562
rect 248952 98504 251914 98560
rect 251970 98504 251975 98560
rect 248952 98502 251975 98504
rect 321908 98502 324268 98562
rect 251909 98499 251975 98502
rect 324262 98500 324268 98502
rect 324332 98500 324338 98564
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 214005 98363 214071 98366
rect 249374 98364 249380 98428
rect 249444 98426 249450 98428
rect 249444 98366 296730 98426
rect 249444 98364 249450 98366
rect 296670 98290 296730 98366
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 296670 98230 310040 98290
rect 251817 98018 251883 98021
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 248952 98016 251883 98018
rect 248952 97960 251822 98016
rect 251878 97960 251883 98016
rect 248952 97958 251883 97960
rect 213913 97955 213979 97958
rect 251817 97955 251883 97958
rect 306925 97882 306991 97885
rect 324405 97882 324471 97885
rect 306925 97880 310040 97882
rect 306925 97824 306930 97880
rect 306986 97824 310040 97880
rect 306925 97822 310040 97824
rect 321908 97880 324471 97882
rect 321908 97824 324410 97880
rect 324466 97824 324471 97880
rect 321908 97822 324471 97824
rect 306925 97819 306991 97822
rect 324405 97819 324471 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect 252185 97610 252251 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 248952 97608 252251 97610
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 214557 97066 214623 97069
rect 217182 97066 217242 97580
rect 248952 97552 252190 97608
rect 252246 97552 252251 97608
rect 248952 97550 252251 97552
rect 252185 97547 252251 97550
rect 307569 97474 307635 97477
rect 307569 97472 310040 97474
rect 307569 97416 307574 97472
rect 307630 97416 310040 97472
rect 307569 97414 310040 97416
rect 307569 97411 307635 97414
rect 251357 97066 251423 97069
rect 251950 97066 251956 97068
rect 214557 97064 217242 97066
rect 214557 97008 214562 97064
rect 214618 97008 217242 97064
rect 214557 97006 217242 97008
rect 248952 97064 251956 97066
rect 248952 97008 251362 97064
rect 251418 97008 251956 97064
rect 248952 97006 251956 97008
rect 214557 97003 214623 97006
rect 251357 97003 251423 97006
rect 251950 97004 251956 97006
rect 252020 97004 252026 97068
rect 306966 97004 306972 97068
rect 307036 97066 307042 97068
rect 324313 97066 324379 97069
rect 307036 97006 310040 97066
rect 321908 97064 324379 97066
rect 321908 97008 324318 97064
rect 324374 97008 324379 97064
rect 321908 97006 324379 97008
rect 307036 97004 307042 97006
rect 324313 97003 324379 97006
rect 214833 96658 214899 96661
rect 217182 96658 217242 96900
rect 249149 96658 249215 96661
rect 252001 96658 252067 96661
rect 214833 96656 217242 96658
rect 214833 96600 214838 96656
rect 214894 96600 217242 96656
rect 214833 96598 217242 96600
rect 248952 96656 252067 96658
rect 248952 96600 249154 96656
rect 249210 96600 252006 96656
rect 252062 96600 252067 96656
rect 248952 96598 252067 96600
rect 214833 96595 214899 96598
rect 249149 96595 249215 96598
rect 252001 96595 252067 96598
rect 307661 96658 307727 96661
rect 321461 96658 321527 96661
rect 307661 96656 310040 96658
rect 307661 96600 307666 96656
rect 307722 96600 310040 96656
rect 307661 96598 310040 96600
rect 321461 96656 321570 96658
rect 321461 96600 321466 96656
rect 321522 96600 321570 96656
rect 307661 96595 307727 96598
rect 321461 96595 321570 96600
rect 321510 96356 321570 96595
rect 396717 96522 396783 96525
rect 493910 96522 493916 96524
rect 396717 96520 493916 96522
rect 396717 96464 396722 96520
rect 396778 96464 493916 96520
rect 396717 96462 493916 96464
rect 396717 96459 396783 96462
rect 493910 96460 493916 96462
rect 493980 96460 493986 96524
rect 213913 95842 213979 95845
rect 217182 95842 217242 96356
rect 251265 96250 251331 96253
rect 248860 96248 251331 96250
rect 248860 96192 251270 96248
rect 251326 96192 251331 96248
rect 248860 96190 251331 96192
rect 251265 96187 251331 96190
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 213913 95840 217242 95842
rect 213913 95784 213918 95840
rect 213974 95784 217242 95840
rect 213913 95782 217242 95784
rect 213913 95779 213979 95782
rect 188981 95162 189047 95165
rect 321502 95162 321508 95164
rect 188981 95160 321508 95162
rect 188981 95104 188986 95160
rect 189042 95104 321508 95160
rect 188981 95102 321508 95104
rect 188981 95099 189047 95102
rect 321502 95100 321508 95102
rect 321572 95100 321578 95164
rect 66161 94890 66227 94893
rect 216121 94890 216187 94893
rect 66161 94888 216187 94890
rect 66161 94832 66166 94888
rect 66222 94832 216126 94888
rect 216182 94832 216187 94888
rect 66161 94830 216187 94832
rect 66161 94827 66227 94830
rect 216121 94827 216187 94830
rect 85573 94756 85639 94757
rect 112345 94756 112411 94757
rect 122833 94756 122899 94757
rect 124489 94756 124555 94757
rect 85528 94692 85534 94756
rect 85598 94754 85639 94756
rect 85598 94752 85690 94754
rect 85634 94696 85690 94752
rect 85598 94694 85690 94696
rect 85598 94692 85639 94694
rect 112320 94692 112326 94756
rect 112390 94754 112411 94756
rect 112390 94752 112482 94754
rect 112406 94696 112482 94752
rect 112390 94694 112482 94696
rect 112390 94692 112411 94694
rect 122792 94692 122798 94756
rect 122862 94754 122899 94756
rect 122862 94752 122954 94754
rect 122894 94696 122954 94752
rect 122862 94694 122954 94696
rect 122862 94692 122899 94694
rect 124424 94692 124430 94756
rect 124494 94754 124555 94756
rect 124494 94752 124586 94754
rect 124550 94696 124586 94752
rect 124494 94694 124586 94696
rect 124494 94692 124555 94694
rect 151486 94692 151492 94756
rect 151556 94754 151562 94756
rect 151760 94754 151766 94756
rect 151556 94694 151766 94754
rect 151556 94692 151562 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 85573 94691 85639 94692
rect 112345 94691 112411 94692
rect 122833 94691 122899 94692
rect 124489 94691 124555 94692
rect 67357 93802 67423 93805
rect 214598 93802 214604 93804
rect 67357 93800 214604 93802
rect 67357 93744 67362 93800
rect 67418 93744 214604 93800
rect 67357 93742 214604 93744
rect 67357 93739 67423 93742
rect 214598 93740 214604 93742
rect 214668 93740 214674 93804
rect 151721 93668 151787 93669
rect 151670 93666 151676 93668
rect 151630 93606 151676 93666
rect 151740 93664 151787 93668
rect 151782 93608 151787 93664
rect 151670 93604 151676 93606
rect 151740 93604 151787 93608
rect 151721 93603 151787 93604
rect 200757 93666 200823 93669
rect 324262 93666 324268 93668
rect 200757 93664 324268 93666
rect 200757 93608 200762 93664
rect 200818 93608 324268 93664
rect 200757 93606 324268 93608
rect 200757 93603 200823 93606
rect 324262 93604 324268 93606
rect 324332 93604 324338 93668
rect 123201 93532 123267 93533
rect 123150 93530 123156 93532
rect 123110 93470 123156 93530
rect 123220 93528 123267 93532
rect 123262 93472 123267 93528
rect 123150 93468 123156 93470
rect 123220 93468 123267 93472
rect 123201 93467 123267 93468
rect 100569 93260 100635 93261
rect 110137 93260 110203 93261
rect 100518 93196 100524 93260
rect 100588 93258 100635 93260
rect 110086 93258 110092 93260
rect 100588 93256 100680 93258
rect 100630 93200 100680 93256
rect 100588 93198 100680 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 100588 93196 100635 93198
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 100569 93195 100635 93196
rect 110137 93195 110203 93196
rect 74809 92444 74875 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 84326 92380 84332 92444
rect 84396 92442 84402 92444
rect 84837 92442 84903 92445
rect 86769 92444 86835 92445
rect 88057 92444 88123 92445
rect 86718 92442 86724 92444
rect 84396 92440 84903 92442
rect 84396 92384 84842 92440
rect 84898 92384 84903 92440
rect 84396 92382 84903 92384
rect 86678 92382 86724 92442
rect 86788 92440 86835 92444
rect 88006 92442 88012 92444
rect 86830 92384 86835 92440
rect 84396 92380 84402 92382
rect 74809 92379 74875 92380
rect 84837 92379 84903 92382
rect 86718 92380 86724 92382
rect 86788 92380 86835 92384
rect 87966 92382 88012 92442
rect 88076 92440 88123 92444
rect 88118 92384 88123 92440
rect 88006 92380 88012 92382
rect 88076 92380 88123 92384
rect 99966 92380 99972 92444
rect 100036 92442 100042 92444
rect 100109 92442 100175 92445
rect 101949 92444 102015 92445
rect 101949 92442 101996 92444
rect 100036 92440 100175 92442
rect 100036 92384 100114 92440
rect 100170 92384 100175 92440
rect 100036 92382 100175 92384
rect 101904 92440 101996 92442
rect 101904 92384 101954 92440
rect 101904 92382 101996 92384
rect 100036 92380 100042 92382
rect 86769 92379 86835 92380
rect 88057 92379 88123 92380
rect 100109 92379 100175 92382
rect 101949 92380 101996 92382
rect 102060 92380 102066 92444
rect 102726 92380 102732 92444
rect 102796 92442 102802 92444
rect 103421 92442 103487 92445
rect 104433 92444 104499 92445
rect 105721 92444 105787 92445
rect 102796 92440 103487 92442
rect 102796 92384 103426 92440
rect 103482 92384 103487 92440
rect 102796 92382 103487 92384
rect 102796 92380 102802 92382
rect 101949 92379 102015 92380
rect 103421 92379 103487 92382
rect 104382 92380 104388 92444
rect 104452 92442 104499 92444
rect 104452 92440 104544 92442
rect 104494 92384 104544 92440
rect 104452 92382 104544 92384
rect 104452 92380 104499 92382
rect 105670 92380 105676 92444
rect 105740 92442 105787 92444
rect 105740 92440 105832 92442
rect 105782 92384 105832 92440
rect 105740 92382 105832 92384
rect 105740 92380 105787 92382
rect 106590 92380 106596 92444
rect 106660 92442 106666 92444
rect 107561 92442 107627 92445
rect 106660 92440 107627 92442
rect 106660 92384 107566 92440
rect 107622 92384 107627 92440
rect 106660 92382 107627 92384
rect 106660 92380 106666 92382
rect 104433 92379 104499 92380
rect 105721 92379 105787 92380
rect 107561 92379 107627 92382
rect 107694 92380 107700 92444
rect 107764 92442 107770 92444
rect 107929 92442 107995 92445
rect 107764 92440 107995 92442
rect 107764 92384 107934 92440
rect 107990 92384 107995 92440
rect 107764 92382 107995 92384
rect 107764 92380 107770 92382
rect 107929 92379 107995 92382
rect 108062 92380 108068 92444
rect 108132 92442 108138 92444
rect 108297 92442 108363 92445
rect 108132 92440 108363 92442
rect 108132 92384 108302 92440
rect 108358 92384 108363 92440
rect 108132 92382 108363 92384
rect 108132 92380 108138 92382
rect 108297 92379 108363 92382
rect 109166 92380 109172 92444
rect 109236 92442 109242 92444
rect 110045 92442 110111 92445
rect 110689 92444 110755 92445
rect 110638 92442 110644 92444
rect 109236 92440 110111 92442
rect 109236 92384 110050 92440
rect 110106 92384 110111 92440
rect 109236 92382 110111 92384
rect 110598 92382 110644 92442
rect 110708 92440 110755 92444
rect 110750 92384 110755 92440
rect 109236 92380 109242 92382
rect 110045 92379 110111 92382
rect 110638 92380 110644 92382
rect 110708 92380 110755 92384
rect 113214 92380 113220 92444
rect 113284 92442 113290 92444
rect 113817 92442 113883 92445
rect 119337 92444 119403 92445
rect 119286 92442 119292 92444
rect 113284 92440 113883 92442
rect 113284 92384 113822 92440
rect 113878 92384 113883 92440
rect 113284 92382 113883 92384
rect 119246 92382 119292 92442
rect 119356 92440 119403 92444
rect 119398 92384 119403 92440
rect 113284 92380 113290 92382
rect 110689 92379 110755 92380
rect 113817 92379 113883 92382
rect 119286 92380 119292 92382
rect 119356 92380 119403 92384
rect 119654 92380 119660 92444
rect 119724 92442 119730 92444
rect 119889 92442 119955 92445
rect 129457 92444 129523 92445
rect 133137 92444 133203 92445
rect 136081 92444 136147 92445
rect 151537 92444 151603 92445
rect 152089 92444 152155 92445
rect 129406 92442 129412 92444
rect 119724 92440 119955 92442
rect 119724 92384 119894 92440
rect 119950 92384 119955 92440
rect 119724 92382 119955 92384
rect 129366 92382 129412 92442
rect 129476 92440 129523 92444
rect 133086 92442 133092 92444
rect 129518 92384 129523 92440
rect 119724 92380 119730 92382
rect 119337 92379 119403 92380
rect 119889 92379 119955 92382
rect 129406 92380 129412 92382
rect 129476 92380 129523 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 136030 92442 136036 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 151486 92442 151492 92444
rect 136142 92384 136147 92440
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 152038 92442 152044 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 129457 92379 129523 92380
rect 133137 92379 133203 92380
rect 136081 92379 136147 92380
rect 151537 92379 151603 92380
rect 152089 92379 152155 92380
rect 100702 92244 100708 92308
rect 100772 92306 100778 92308
rect 101857 92306 101923 92309
rect 100772 92304 101923 92306
rect 100772 92248 101862 92304
rect 101918 92248 101923 92304
rect 100772 92246 101923 92248
rect 100772 92244 100778 92246
rect 101857 92243 101923 92246
rect 102542 92244 102548 92308
rect 102612 92306 102618 92308
rect 103329 92306 103395 92309
rect 104617 92308 104683 92309
rect 102612 92304 103395 92306
rect 102612 92248 103334 92304
rect 103390 92248 103395 92304
rect 102612 92246 103395 92248
rect 102612 92244 102618 92246
rect 103329 92243 103395 92246
rect 104566 92244 104572 92308
rect 104636 92306 104683 92308
rect 104636 92304 104728 92306
rect 104678 92248 104728 92304
rect 104636 92246 104728 92248
rect 104636 92244 104683 92246
rect 105486 92244 105492 92308
rect 105556 92306 105562 92308
rect 106181 92306 106247 92309
rect 105556 92304 106247 92306
rect 105556 92248 106186 92304
rect 106242 92248 106247 92304
rect 105556 92246 106247 92248
rect 105556 92244 105562 92246
rect 104617 92243 104683 92244
rect 106181 92243 106247 92246
rect 106406 92244 106412 92308
rect 106476 92306 106482 92308
rect 107469 92306 107535 92309
rect 106476 92304 107535 92306
rect 106476 92248 107474 92304
rect 107530 92248 107535 92304
rect 106476 92246 107535 92248
rect 106476 92244 106482 92246
rect 107469 92243 107535 92246
rect 116710 92244 116716 92308
rect 116780 92306 116786 92308
rect 198181 92306 198247 92309
rect 116780 92304 198247 92306
rect 116780 92248 198186 92304
rect 198242 92248 198247 92304
rect 116780 92246 198247 92248
rect 116780 92244 116786 92246
rect 198181 92243 198247 92246
rect 101806 92108 101812 92172
rect 101876 92170 101882 92172
rect 102041 92170 102107 92173
rect 117129 92172 117195 92173
rect 117078 92170 117084 92172
rect 101876 92168 102107 92170
rect 101876 92112 102046 92168
rect 102102 92112 102107 92168
rect 101876 92110 102107 92112
rect 117038 92110 117084 92170
rect 117148 92168 117195 92172
rect 117190 92112 117195 92168
rect 101876 92108 101882 92110
rect 102041 92107 102107 92110
rect 117078 92108 117084 92110
rect 117148 92108 117195 92112
rect 117129 92107 117195 92108
rect 88977 91764 89043 91765
rect 88926 91762 88932 91764
rect 88886 91702 88932 91762
rect 88996 91760 89043 91764
rect 89038 91704 89043 91760
rect 88926 91700 88932 91702
rect 88996 91700 89043 91704
rect 111190 91700 111196 91764
rect 111260 91762 111266 91764
rect 111609 91762 111675 91765
rect 111260 91760 111675 91762
rect 111260 91704 111614 91760
rect 111670 91704 111675 91760
rect 111260 91702 111675 91704
rect 111260 91700 111266 91702
rect 88977 91699 89043 91700
rect 111609 91699 111675 91702
rect 114502 91700 114508 91764
rect 114572 91762 114578 91764
rect 114572 91702 122850 91762
rect 114572 91700 114578 91702
rect 118049 91628 118115 91629
rect 117998 91626 118004 91628
rect 117958 91566 118004 91626
rect 118068 91624 118115 91628
rect 118110 91568 118115 91624
rect 117998 91564 118004 91566
rect 118068 91564 118115 91568
rect 120574 91564 120580 91628
rect 120644 91626 120650 91628
rect 120901 91626 120967 91629
rect 120644 91624 120967 91626
rect 120644 91568 120906 91624
rect 120962 91568 120967 91624
rect 120644 91566 120967 91568
rect 122790 91626 122850 91702
rect 134374 91700 134380 91764
rect 134444 91762 134450 91764
rect 134885 91762 134951 91765
rect 134444 91760 134951 91762
rect 134444 91704 134890 91760
rect 134946 91704 134951 91760
rect 134444 91702 134951 91704
rect 134444 91700 134450 91702
rect 134885 91699 134951 91702
rect 207749 91626 207815 91629
rect 122790 91624 207815 91626
rect 122790 91568 207754 91624
rect 207810 91568 207815 91624
rect 122790 91566 207815 91568
rect 120644 91564 120650 91566
rect 118049 91563 118115 91564
rect 120901 91563 120967 91566
rect 207749 91563 207815 91566
rect 97206 91428 97212 91492
rect 97276 91490 97282 91492
rect 97441 91490 97507 91493
rect 97276 91488 97507 91490
rect 97276 91432 97446 91488
rect 97502 91432 97507 91488
rect 97276 91430 97507 91432
rect 97276 91428 97282 91430
rect 97441 91427 97507 91430
rect 98126 91428 98132 91492
rect 98196 91490 98202 91492
rect 99189 91490 99255 91493
rect 98196 91488 99255 91490
rect 98196 91432 99194 91488
rect 99250 91432 99255 91488
rect 98196 91430 99255 91432
rect 98196 91428 98202 91430
rect 99189 91427 99255 91430
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99281 91354 99347 91357
rect 98564 91352 99347 91354
rect 98564 91296 99286 91352
rect 99342 91296 99347 91352
rect 98564 91294 99347 91296
rect 98564 91292 98570 91294
rect 99281 91291 99347 91294
rect 115749 91356 115815 91357
rect 122097 91356 122163 91357
rect 126697 91356 126763 91357
rect 115749 91352 115796 91356
rect 115860 91354 115866 91356
rect 122046 91354 122052 91356
rect 115749 91296 115754 91352
rect 115749 91292 115796 91296
rect 115860 91294 115906 91354
rect 122006 91294 122052 91354
rect 122116 91352 122163 91356
rect 126646 91354 126652 91356
rect 122158 91296 122163 91352
rect 115860 91292 115866 91294
rect 122046 91292 122052 91294
rect 122116 91292 122163 91296
rect 126606 91294 126652 91354
rect 126716 91352 126763 91356
rect 126758 91296 126763 91352
rect 126646 91292 126652 91294
rect 126716 91292 126763 91296
rect 115749 91291 115815 91292
rect 122097 91291 122163 91292
rect 126697 91291 126763 91292
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90633 91218 90699 91221
rect 90284 91216 90699 91218
rect 90284 91160 90638 91216
rect 90694 91160 90699 91216
rect 90284 91158 90699 91160
rect 90284 91156 90290 91158
rect 90633 91155 90699 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97073 91218 97139 91221
rect 99097 91220 99163 91221
rect 99046 91218 99052 91220
rect 96724 91216 97139 91218
rect 96724 91160 97078 91216
rect 97134 91160 97139 91216
rect 96724 91158 97139 91160
rect 99006 91158 99052 91218
rect 99116 91216 99163 91220
rect 99158 91160 99163 91216
rect 96724 91156 96730 91158
rect 97073 91155 97139 91158
rect 99046 91156 99052 91158
rect 99116 91156 99163 91160
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 99097 91155 99163 91156
rect 110321 91155 110387 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 114369 91220 114435 91221
rect 114318 91218 114324 91220
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 114278 91158 114324 91218
rect 114388 91216 114435 91220
rect 114430 91160 114435 91216
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 114318 91156 114324 91158
rect 114388 91156 114435 91160
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115289 91218 115355 91221
rect 114940 91216 115355 91218
rect 114940 91160 115294 91216
rect 115350 91160 115355 91216
rect 114940 91158 115355 91160
rect 114940 91156 114946 91158
rect 114369 91155 114435 91156
rect 115289 91155 115355 91158
rect 115422 91156 115428 91220
rect 115492 91218 115498 91220
rect 115841 91218 115907 91221
rect 115492 91216 115907 91218
rect 115492 91160 115846 91216
rect 115902 91160 115907 91216
rect 115492 91158 115907 91160
rect 115492 91156 115498 91158
rect 115841 91155 115907 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 118601 91155 118667 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 122741 91218 122807 91221
rect 124121 91220 124187 91221
rect 124070 91218 124076 91220
rect 121748 91216 122807 91218
rect 121748 91160 122746 91216
rect 122802 91160 122807 91216
rect 121748 91158 122807 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 124182 91160 124187 91216
rect 121748 91156 121754 91158
rect 122741 91155 122807 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 124121 91155 124187 91156
rect 125501 91155 125567 91158
rect 125726 91156 125732 91220
rect 125796 91218 125802 91220
rect 126053 91218 126119 91221
rect 125796 91216 126119 91218
rect 125796 91160 126058 91216
rect 126114 91160 126119 91216
rect 125796 91158 126119 91160
rect 125796 91156 125802 91158
rect 126053 91155 126119 91158
rect 126462 91156 126468 91220
rect 126532 91218 126538 91220
rect 126881 91218 126947 91221
rect 126532 91216 126947 91218
rect 126532 91160 126886 91216
rect 126942 91160 126947 91216
rect 126532 91158 126947 91160
rect 126532 91156 126538 91158
rect 126881 91155 126947 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 127636 91156 127642 91158
rect 128261 91155 128327 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 151302 91156 151308 91220
rect 151372 91218 151378 91220
rect 151629 91218 151695 91221
rect 151372 91216 151695 91218
rect 151372 91160 151634 91216
rect 151690 91160 151695 91216
rect 151372 91158 151695 91160
rect 151372 91156 151378 91158
rect 151629 91155 151695 91158
rect 67449 91082 67515 91085
rect 214414 91082 214420 91084
rect 67449 91080 214420 91082
rect 67449 91024 67454 91080
rect 67510 91024 214420 91080
rect 67449 91022 214420 91024
rect 67449 91019 67515 91022
rect 214414 91020 214420 91022
rect 214484 91020 214490 91084
rect 132350 90884 132356 90948
rect 132420 90946 132426 90948
rect 168966 90946 168972 90948
rect 132420 90886 168972 90946
rect 132420 90884 132426 90886
rect 168966 90884 168972 90886
rect 169036 90884 169042 90948
rect 67265 89722 67331 89725
rect 207841 89722 207907 89725
rect 67265 89720 207907 89722
rect 67265 89664 67270 89720
rect 67326 89664 207846 89720
rect 207902 89664 207907 89720
rect 67265 89662 207907 89664
rect 67265 89659 67331 89662
rect 207841 89659 207907 89662
rect 105721 88226 105787 88229
rect 180241 88226 180307 88229
rect 105721 88224 180307 88226
rect 105721 88168 105726 88224
rect 105782 88168 180246 88224
rect 180302 88168 180307 88224
rect 105721 88166 180307 88168
rect 105721 88163 105787 88166
rect 180241 88163 180307 88166
rect 191230 87484 191236 87548
rect 191300 87546 191306 87548
rect 255313 87546 255379 87549
rect 334750 87546 334756 87548
rect 191300 87544 334756 87546
rect 191300 87488 255318 87544
rect 255374 87488 334756 87544
rect 191300 87486 334756 87488
rect 191300 87484 191306 87486
rect 255313 87483 255379 87486
rect 334750 87484 334756 87486
rect 334820 87484 334826 87548
rect 108297 86866 108363 86869
rect 166390 86866 166396 86868
rect 108297 86864 166396 86866
rect 108297 86808 108302 86864
rect 108358 86808 166396 86864
rect 108297 86806 166396 86808
rect 108297 86803 108363 86806
rect 166390 86804 166396 86806
rect 166460 86804 166466 86868
rect 193806 86124 193812 86188
rect 193876 86186 193882 86188
rect 331949 86186 332015 86189
rect 193876 86184 332015 86186
rect 193876 86128 331954 86184
rect 332010 86128 332015 86184
rect 193876 86126 332015 86128
rect 193876 86124 193882 86126
rect 331949 86123 332015 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 242157 84962 242223 84965
rect 342846 84962 342852 84964
rect 242157 84960 342852 84962
rect 242157 84904 242162 84960
rect 242218 84904 342852 84960
rect 242157 84902 342852 84904
rect 242157 84899 242223 84902
rect 342846 84900 342852 84902
rect 342916 84900 342922 84964
rect 178677 84826 178743 84829
rect 307150 84826 307156 84828
rect 178677 84824 307156 84826
rect -960 84690 480 84780
rect 178677 84768 178682 84824
rect 178738 84768 307156 84824
rect 178677 84766 307156 84768
rect 178677 84763 178743 84766
rect 307150 84764 307156 84766
rect 307220 84764 307226 84828
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 113081 84146 113147 84149
rect 169150 84146 169156 84148
rect 113081 84144 169156 84146
rect 113081 84088 113086 84144
rect 113142 84088 169156 84144
rect 113081 84086 169156 84088
rect 113081 84083 113147 84086
rect 169150 84084 169156 84086
rect 169220 84084 169226 84148
rect 173014 83404 173020 83468
rect 173084 83466 173090 83468
rect 261661 83466 261727 83469
rect 173084 83464 261727 83466
rect 173084 83408 261666 83464
rect 261722 83408 261727 83464
rect 173084 83406 261727 83408
rect 173084 83404 173090 83406
rect 261661 83403 261727 83406
rect 274081 83466 274147 83469
rect 340270 83466 340276 83468
rect 274081 83464 340276 83466
rect 274081 83408 274086 83464
rect 274142 83408 340276 83464
rect 274081 83406 340276 83408
rect 274081 83403 274147 83406
rect 340270 83404 340276 83406
rect 340340 83404 340346 83468
rect 115841 82786 115907 82789
rect 170438 82786 170444 82788
rect 115841 82784 170444 82786
rect 115841 82728 115846 82784
rect 115902 82728 170444 82784
rect 115841 82726 170444 82728
rect 115841 82723 115907 82726
rect 170438 82724 170444 82726
rect 170508 82724 170514 82788
rect 195094 82044 195100 82108
rect 195164 82106 195170 82108
rect 324313 82106 324379 82109
rect 195164 82104 324379 82106
rect 195164 82048 324318 82104
rect 324374 82048 324379 82104
rect 195164 82046 324379 82048
rect 195164 82044 195170 82046
rect 324313 82043 324379 82046
rect 99097 81426 99163 81429
rect 172094 81426 172100 81428
rect 99097 81424 172100 81426
rect 99097 81368 99102 81424
rect 99158 81368 172100 81424
rect 99097 81366 172100 81368
rect 99097 81363 99163 81366
rect 172094 81364 172100 81366
rect 172164 81364 172170 81428
rect 217317 80746 217383 80749
rect 251173 80746 251239 80749
rect 332910 80746 332916 80748
rect 217317 80744 332916 80746
rect 217317 80688 217322 80744
rect 217378 80688 251178 80744
rect 251234 80688 332916 80744
rect 217317 80686 332916 80688
rect 217317 80683 217383 80686
rect 251173 80683 251239 80686
rect 332910 80684 332916 80686
rect 332980 80684 332986 80748
rect 99189 80066 99255 80069
rect 166206 80066 166212 80068
rect 99189 80064 166212 80066
rect 99189 80008 99194 80064
rect 99250 80008 166212 80064
rect 99189 80006 166212 80008
rect 99189 80003 99255 80006
rect 166206 80004 166212 80006
rect 166276 80004 166282 80068
rect 260281 79386 260347 79389
rect 335854 79386 335860 79388
rect 260281 79384 335860 79386
rect 260281 79328 260286 79384
rect 260342 79328 335860 79384
rect 260281 79326 335860 79328
rect 260281 79323 260347 79326
rect 335854 79324 335860 79326
rect 335924 79324 335930 79388
rect 101857 78570 101923 78573
rect 168230 78570 168236 78572
rect 101857 78568 168236 78570
rect 101857 78512 101862 78568
rect 101918 78512 168236 78568
rect 101857 78510 168236 78512
rect 101857 78507 101923 78510
rect 168230 78508 168236 78510
rect 168300 78508 168306 78572
rect 338246 78508 338252 78572
rect 338316 78570 338322 78572
rect 339401 78570 339467 78573
rect 338316 78568 339467 78570
rect 338316 78512 339406 78568
rect 339462 78512 339467 78568
rect 338316 78510 339467 78512
rect 338316 78508 338322 78510
rect 339401 78507 339467 78510
rect 107561 78434 107627 78437
rect 170254 78434 170260 78436
rect 107561 78432 170260 78434
rect 107561 78376 107566 78432
rect 107622 78376 170260 78432
rect 107561 78374 170260 78376
rect 107561 78371 107627 78374
rect 170254 78372 170260 78374
rect 170324 78372 170330 78436
rect 300710 76468 300716 76532
rect 300780 76530 300786 76532
rect 473353 76530 473419 76533
rect 300780 76528 473419 76530
rect 300780 76472 473358 76528
rect 473414 76472 473419 76528
rect 300780 76470 473419 76472
rect 300780 76468 300786 76470
rect 473353 76467 473419 76470
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 258574 67492 258580 67556
rect 258644 67554 258650 67556
rect 262213 67554 262279 67557
rect 258644 67552 262279 67554
rect 258644 67496 262218 67552
rect 262274 67496 262279 67552
rect 258644 67494 262279 67496
rect 258644 67492 258650 67494
rect 262213 67491 262279 67494
rect 61694 62868 61700 62932
rect 61764 62930 61770 62932
rect 243537 62930 243603 62933
rect 61764 62928 243603 62930
rect 61764 62872 243542 62928
rect 243598 62872 243603 62928
rect 61764 62870 243603 62872
rect 61764 62868 61770 62870
rect 243537 62867 243603 62870
rect 62982 62732 62988 62796
rect 63052 62794 63058 62796
rect 280889 62794 280955 62797
rect 63052 62792 280955 62794
rect 63052 62736 280894 62792
rect 280950 62736 280955 62792
rect 63052 62734 280955 62736
rect 63052 62732 63058 62734
rect 280889 62731 280955 62734
rect 66110 59876 66116 59940
rect 66180 59938 66186 59940
rect 308397 59938 308463 59941
rect 66180 59936 308463 59938
rect 66180 59880 308402 59936
rect 308458 59880 308463 59936
rect 66180 59878 308463 59880
rect 66180 59876 66186 59878
rect 308397 59875 308463 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 77293 51778 77359 51781
rect 257286 51778 257292 51780
rect 77293 51776 257292 51778
rect 77293 51720 77298 51776
rect 77354 51720 257292 51776
rect 77293 51718 257292 51720
rect 77293 51715 77359 51718
rect 257286 51716 257292 51718
rect 257356 51716 257362 51780
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 189942 46140 189948 46204
rect 190012 46202 190018 46204
rect 278037 46202 278103 46205
rect 340873 46204 340939 46205
rect 190012 46200 278103 46202
rect 190012 46144 278042 46200
rect 278098 46144 278103 46200
rect 190012 46142 278103 46144
rect 190012 46140 190018 46142
rect 278037 46139 278103 46142
rect 340822 46140 340828 46204
rect 340892 46202 340939 46204
rect 340892 46200 340984 46202
rect 340934 46144 340984 46200
rect 583520 46188 584960 46278
rect 340892 46142 340984 46144
rect 340892 46140 340939 46142
rect 340873 46139 340939 46140
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 280889 45522 280955 45525
rect 338614 45522 338620 45524
rect 280889 45520 338620 45522
rect 280889 45464 280894 45520
rect 280950 45464 338620 45520
rect 280889 45462 338620 45464
rect 280889 45459 280955 45462
rect 338614 45460 338620 45462
rect 338684 45460 338690 45524
rect 280153 44298 280219 44301
rect 280889 44298 280955 44301
rect 280153 44296 280955 44298
rect 280153 44240 280158 44296
rect 280214 44240 280894 44296
rect 280950 44240 280955 44296
rect 280153 44238 280955 44240
rect 280153 44235 280219 44238
rect 280889 44235 280955 44238
rect 186814 43420 186820 43484
rect 186884 43482 186890 43484
rect 316677 43482 316743 43485
rect 317321 43482 317387 43485
rect 186884 43480 317387 43482
rect 186884 43424 316682 43480
rect 316738 43424 317326 43480
rect 317382 43424 317387 43480
rect 186884 43422 317387 43424
rect 186884 43420 186890 43422
rect 316677 43419 316743 43422
rect 317321 43419 317387 43422
rect 64454 42196 64460 42260
rect 64524 42258 64530 42260
rect 289169 42258 289235 42261
rect 64524 42256 289235 42258
rect 64524 42200 289174 42256
rect 289230 42200 289235 42256
rect 64524 42198 289235 42200
rect 64524 42196 64530 42198
rect 289169 42195 289235 42198
rect 33133 42122 33199 42125
rect 304206 42122 304212 42124
rect 33133 42120 304212 42122
rect 33133 42064 33138 42120
rect 33194 42064 304212 42120
rect 33133 42062 304212 42064
rect 33133 42059 33199 42062
rect 304206 42060 304212 42062
rect 304276 42060 304282 42124
rect 184054 40564 184060 40628
rect 184124 40626 184130 40628
rect 308489 40626 308555 40629
rect 184124 40624 308555 40626
rect 184124 40568 308494 40624
rect 308550 40568 308555 40624
rect 184124 40566 308555 40568
rect 184124 40564 184130 40566
rect 308489 40563 308555 40566
rect 300669 39540 300735 39541
rect 300669 39538 300716 39540
rect 300624 39536 300716 39538
rect 300624 39480 300674 39536
rect 300624 39478 300716 39480
rect 300669 39476 300716 39478
rect 300780 39476 300786 39540
rect 300669 39475 300735 39476
rect 120073 37906 120139 37909
rect 253054 37906 253060 37908
rect 120073 37904 253060 37906
rect 120073 37848 120078 37904
rect 120134 37848 253060 37904
rect 120073 37846 253060 37848
rect 120073 37843 120139 37846
rect 253054 37844 253060 37846
rect 253124 37844 253130 37908
rect 268326 35124 268332 35188
rect 268396 35186 268402 35188
rect 295425 35186 295491 35189
rect 268396 35184 295491 35186
rect 268396 35128 295430 35184
rect 295486 35128 295491 35184
rect 268396 35126 295491 35128
rect 268396 35124 268402 35126
rect 295425 35123 295491 35126
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 191046 28188 191052 28252
rect 191116 28250 191122 28252
rect 276841 28250 276907 28253
rect 278221 28250 278287 28253
rect 191116 28248 278287 28250
rect 191116 28192 276846 28248
rect 276902 28192 278226 28248
rect 278282 28192 278287 28248
rect 191116 28190 278287 28192
rect 191116 28188 191122 28190
rect 276841 28187 276907 28190
rect 278221 28187 278287 28190
rect 58934 26148 58940 26212
rect 59004 26210 59010 26212
rect 260281 26210 260347 26213
rect 59004 26208 260347 26210
rect 59004 26152 260286 26208
rect 260342 26152 260347 26208
rect 59004 26150 260347 26152
rect 59004 26148 59010 26150
rect 260281 26147 260347 26150
rect 259453 24986 259519 24989
rect 260281 24986 260347 24989
rect 259453 24984 260347 24986
rect 259453 24928 259458 24984
rect 259514 24928 260286 24984
rect 260342 24928 260347 24984
rect 259453 24926 260347 24928
rect 259453 24923 259519 24926
rect 260281 24923 260347 24926
rect 61878 19892 61884 19956
rect 61948 19954 61954 19956
rect 249057 19954 249123 19957
rect 61948 19952 249123 19954
rect 61948 19896 249062 19952
rect 249118 19896 249123 19952
rect 61948 19894 249123 19896
rect 61948 19892 61954 19894
rect 249057 19891 249123 19894
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 17217 18594 17283 18597
rect 306966 18594 306972 18596
rect 17217 18592 306972 18594
rect 17217 18536 17222 18592
rect 17278 18536 306972 18592
rect 17217 18534 306972 18536
rect 17217 18531 17283 18534
rect 306966 18532 306972 18534
rect 307036 18532 307042 18596
rect 42793 17234 42859 17237
rect 305494 17234 305500 17236
rect 42793 17232 305500 17234
rect 42793 17176 42798 17232
rect 42854 17176 305500 17232
rect 42793 17174 305500 17176
rect 42793 17171 42859 17174
rect 305494 17172 305500 17174
rect 305564 17172 305570 17236
rect 337009 15194 337075 15197
rect 494094 15194 494100 15196
rect 337009 15192 494100 15194
rect 337009 15136 337014 15192
rect 337070 15136 494100 15192
rect 337009 15134 494100 15136
rect 337009 15131 337075 15134
rect 494094 15132 494100 15134
rect 494164 15132 494170 15196
rect 39113 14514 39179 14517
rect 255814 14514 255820 14516
rect 39113 14512 255820 14514
rect 39113 14456 39118 14512
rect 39174 14456 255820 14512
rect 39113 14454 255820 14456
rect 39113 14451 39179 14454
rect 255814 14452 255820 14454
rect 255884 14452 255890 14516
rect 340822 11732 340828 11796
rect 340892 11794 340898 11796
rect 342161 11794 342227 11797
rect 340892 11792 342227 11794
rect 340892 11736 342166 11792
rect 342222 11736 342227 11792
rect 340892 11734 342227 11736
rect 340892 11732 340898 11734
rect 342161 11731 342227 11734
rect 30833 11658 30899 11661
rect 249190 11658 249196 11660
rect 30833 11656 249196 11658
rect 30833 11600 30838 11656
rect 30894 11600 249196 11656
rect 30833 11598 249196 11600
rect 30833 11595 30899 11598
rect 249190 11596 249196 11598
rect 249260 11596 249266 11660
rect 20161 10298 20227 10301
rect 249374 10298 249380 10300
rect 20161 10296 249380 10298
rect 20161 10240 20166 10296
rect 20222 10240 249380 10296
rect 20161 10238 249380 10240
rect 20161 10235 20227 10238
rect 249374 10236 249380 10238
rect 249444 10236 249450 10300
rect 354765 8258 354831 8261
rect 499798 8258 499804 8260
rect 354765 8256 499804 8258
rect 354765 8200 354770 8256
rect 354826 8200 499804 8256
rect 354765 8198 499804 8200
rect 354765 8195 354831 8198
rect 499798 8196 499804 8198
rect 499868 8196 499874 8260
rect 340965 7578 341031 7581
rect 354765 7578 354831 7581
rect 340965 7576 354831 7578
rect 340965 7520 340970 7576
rect 341026 7520 354770 7576
rect 354826 7520 354831 7576
rect 340965 7518 354831 7520
rect 340965 7515 341031 7518
rect 354765 7515 354831 7518
rect 188286 6836 188292 6900
rect 188356 6898 188362 6900
rect 268561 6898 268627 6901
rect 188356 6896 268627 6898
rect 188356 6840 268566 6896
rect 268622 6840 268627 6896
rect 188356 6838 268627 6840
rect 188356 6836 188362 6838
rect 268561 6835 268627 6838
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3325 6490 3391 6493
rect -960 6488 3391 6490
rect -960 6432 3330 6488
rect 3386 6432 3391 6488
rect 583520 6476 584960 6566
rect -960 6430 3391 6432
rect -960 6340 480 6430
rect 3325 6427 3391 6430
rect 27705 4858 27771 4861
rect 302734 4858 302740 4860
rect 27705 4856 302740 4858
rect 27705 4800 27710 4856
rect 27766 4800 302740 4856
rect 27705 4798 302740 4800
rect 27705 4795 27771 4798
rect 302734 4796 302740 4798
rect 302804 4796 302810 4860
rect 348417 4042 348483 4045
rect 496854 4042 496860 4044
rect 348417 4040 496860 4042
rect 348417 3984 348422 4040
rect 348478 3984 496860 4040
rect 348417 3982 496860 3984
rect 348417 3979 348483 3982
rect 496854 3980 496860 3982
rect 496924 3980 496930 4044
rect 299565 3634 299631 3637
rect 300761 3634 300827 3637
rect 299565 3632 300827 3634
rect 299565 3576 299570 3632
rect 299626 3576 300766 3632
rect 300822 3576 300827 3632
rect 299565 3574 300827 3576
rect 299565 3571 299631 3574
rect 300761 3571 300827 3574
rect 125869 3362 125935 3365
rect 173934 3362 173940 3364
rect 125869 3360 173940 3362
rect 125869 3304 125874 3360
rect 125930 3304 173940 3360
rect 125869 3302 173940 3304
rect 125869 3299 125935 3302
rect 173934 3300 173940 3302
rect 174004 3300 174010 3364
<< via3 >>
rect 115980 585108 116044 585172
rect 52316 583884 52380 583948
rect 111748 582524 111812 582588
rect 39804 582388 39868 582452
rect 124260 582388 124324 582452
rect 69796 581360 69860 581364
rect 69796 581304 69846 581360
rect 69846 581304 69860 581360
rect 69796 581300 69860 581304
rect 107700 578716 107764 578780
rect 66116 577764 66180 577828
rect 110644 577492 110708 577556
rect 64644 575044 64708 575108
rect 114508 573140 114572 573204
rect 55076 571916 55140 571980
rect 62988 570148 63052 570212
rect 59124 563212 59188 563276
rect 105492 562940 105556 563004
rect 69980 557364 70044 557428
rect 106412 556276 106476 556340
rect 68876 553964 68940 554028
rect 61884 549476 61948 549540
rect 107884 542676 107948 542740
rect 107700 537372 107764 537436
rect 69612 536828 69676 536892
rect 101260 536828 101324 536892
rect 101996 536828 102060 536892
rect 115980 534652 116044 534716
rect 110828 529076 110892 529140
rect 44036 526356 44100 526420
rect 143580 499564 143644 499628
rect 115980 497388 116044 497452
rect 111748 496028 111812 496092
rect 50844 493308 50908 493372
rect 52316 493308 52380 493372
rect 111748 492764 111812 492828
rect 124260 491812 124324 491876
rect 99236 491676 99300 491740
rect 103836 490588 103900 490652
rect 57836 490452 57900 490516
rect 108988 490452 109052 490516
rect 53604 489092 53668 489156
rect 52316 487188 52380 487252
rect 69060 486644 69124 486708
rect 110644 486372 110708 486436
rect 122052 486372 122116 486436
rect 39804 485692 39868 485756
rect 69796 485888 69860 485892
rect 69796 485832 69846 485888
rect 69846 485832 69860 485888
rect 69796 485828 69860 485832
rect 113036 485012 113100 485076
rect 65932 484604 65996 484668
rect 70348 484604 70412 484668
rect 99420 484468 99484 484532
rect 124076 483108 124140 483172
rect 114508 482352 114572 482356
rect 114508 482296 114558 482352
rect 114558 482296 114572 482352
rect 114508 482292 114572 482296
rect 113036 480796 113100 480860
rect 66116 478892 66180 478956
rect 64644 477396 64708 477460
rect 68692 477048 68756 477052
rect 68692 476992 68742 477048
rect 68742 476992 68756 477048
rect 68692 476988 68756 476992
rect 104940 474676 105004 474740
rect 105492 474676 105556 474740
rect 110828 474676 110892 474740
rect 66116 474268 66180 474332
rect 55076 473180 55140 473244
rect 62988 471548 63052 471612
rect 61700 471276 61764 471340
rect 62988 471276 63052 471340
rect 62988 467876 63052 467940
rect 59124 463796 59188 463860
rect 106412 464204 106476 464268
rect 60596 463524 60660 463588
rect 60596 462844 60660 462908
rect 106780 462844 106844 462908
rect 146524 462300 146588 462364
rect 111748 459640 111812 459644
rect 111748 459584 111762 459640
rect 111762 459584 111812 459640
rect 111748 459580 111812 459584
rect 68508 454004 68572 454068
rect 68876 454004 68940 454068
rect 126836 453868 126900 453932
rect 107884 451284 107948 451348
rect 61884 449788 61948 449852
rect 141924 449924 141988 449988
rect 61884 448564 61948 448628
rect 64644 447748 64708 447812
rect 101996 446524 102060 446588
rect 61884 445768 61948 445772
rect 61884 445712 61934 445768
rect 61934 445712 61948 445768
rect 61884 445708 61948 445712
rect 99420 442988 99484 443052
rect 101260 442308 101324 442372
rect 101260 441900 101324 441964
rect 69612 440676 69676 440740
rect 70164 439996 70228 440060
rect 106780 439044 106844 439108
rect 103836 438908 103900 438972
rect 44036 438636 44100 438700
rect 115980 437412 116044 437476
rect 105492 437276 105556 437340
rect 65932 436732 65996 436796
rect 99052 435916 99116 435980
rect 53604 435780 53668 435844
rect 69060 435236 69124 435300
rect 57836 434556 57900 434620
rect 120028 407764 120092 407828
rect 338252 407084 338316 407148
rect 122604 405044 122668 405108
rect 340092 404364 340156 404428
rect 168972 403004 169036 403068
rect 160692 401644 160756 401708
rect 68692 401372 68756 401436
rect 68876 400284 68940 400348
rect 118004 399604 118068 399668
rect 128676 399468 128740 399532
rect 124260 397972 124324 398036
rect 68876 396204 68940 396268
rect 53788 395932 53852 395996
rect 133828 394844 133892 394908
rect 114692 392532 114756 392596
rect 129780 391172 129844 391236
rect 52316 390688 52380 390692
rect 52316 390632 52330 390688
rect 52330 390632 52380 390688
rect 52316 390628 52380 390632
rect 68692 390628 68756 390692
rect 115980 389812 116044 389876
rect 170260 389812 170324 389876
rect 57836 389192 57900 389196
rect 57836 389136 57886 389192
rect 57886 389136 57900 389192
rect 57836 389132 57900 389136
rect 143580 388996 143644 389060
rect 108988 388860 109052 388924
rect 191236 387772 191300 387836
rect 50844 387636 50908 387700
rect 118740 387636 118804 387700
rect 118740 386956 118804 387020
rect 58940 386276 59004 386340
rect 121684 385732 121748 385796
rect 340828 385596 340892 385660
rect 69796 385324 69860 385388
rect 69980 383148 70044 383212
rect 61700 382196 61764 382260
rect 61516 381032 61580 381036
rect 61516 380976 61530 381032
rect 61530 380976 61580 381032
rect 61516 380972 61580 380976
rect 122052 380156 122116 380220
rect 140820 380156 140884 380220
rect 66116 379672 66180 379676
rect 66116 379616 66166 379672
rect 66166 379616 66180 379672
rect 66116 379612 66180 379616
rect 124076 378720 124140 378724
rect 124076 378664 124126 378720
rect 124126 378664 124140 378720
rect 124076 378660 124140 378664
rect 128676 378660 128740 378724
rect 115980 378524 116044 378588
rect 115428 377300 115492 377364
rect 122052 376756 122116 376820
rect 115428 376408 115492 376412
rect 115428 376352 115478 376408
rect 115478 376352 115492 376408
rect 115428 376348 115492 376352
rect 321508 375396 321572 375460
rect 188292 374580 188356 374644
rect 118004 372736 118068 372740
rect 118004 372680 118054 372736
rect 118054 372680 118068 372736
rect 118004 372676 118068 372680
rect 62988 371316 63052 371380
rect 65932 371860 65996 371924
rect 69796 369820 69860 369884
rect 332916 369820 332980 369884
rect 59124 368384 59188 368388
rect 59124 368328 59174 368384
rect 59174 368328 59188 368384
rect 59124 368324 59188 368328
rect 60596 366964 60660 367028
rect 62988 366964 63052 367028
rect 62988 365740 63052 365804
rect 66116 365664 66180 365668
rect 66116 365608 66130 365664
rect 66130 365608 66180 365664
rect 66116 365604 66180 365608
rect 66116 364652 66180 364716
rect 330340 364380 330404 364444
rect 184060 363564 184124 363628
rect 320220 363156 320284 363220
rect 345612 361932 345676 361996
rect 320036 361796 320100 361860
rect 200620 361660 200684 361724
rect 146524 360360 146588 360364
rect 146524 360304 146538 360360
rect 146538 360304 146588 360360
rect 146524 360300 146588 360304
rect 334572 360300 334636 360364
rect 199332 360164 199396 360228
rect 173020 359348 173084 359412
rect 120028 358668 120092 358732
rect 197860 358260 197924 358324
rect 331260 357988 331324 358052
rect 68692 356900 68756 356964
rect 195100 356628 195164 356692
rect 53788 355404 53852 355468
rect 320036 355268 320100 355332
rect 327028 354180 327092 354244
rect 137140 353908 137204 353972
rect 199332 353908 199396 353972
rect 66668 353228 66732 353292
rect 321508 352140 321572 352204
rect 191052 351052 191116 351116
rect 68876 350100 68940 350164
rect 64460 349888 64524 349892
rect 64460 349832 64474 349888
rect 64474 349832 64524 349888
rect 64460 349828 64524 349832
rect 64644 349752 64708 349756
rect 64644 349696 64658 349752
rect 64658 349696 64708 349752
rect 64644 349692 64708 349696
rect 186820 348332 186884 348396
rect 61884 346564 61948 346628
rect 200620 346292 200684 346356
rect 189948 345612 190012 345676
rect 126836 343632 126900 343636
rect 126836 343576 126850 343632
rect 126850 343576 126900 343632
rect 126836 343572 126900 343576
rect 133092 342892 133156 342956
rect 193812 342892 193876 342956
rect 120028 342076 120092 342140
rect 70532 341668 70596 341732
rect 69612 340036 69676 340100
rect 124260 339356 124324 339420
rect 66668 338676 66732 338740
rect 122604 337996 122668 338060
rect 142292 338056 142356 338060
rect 142292 338000 142306 338056
rect 142306 338000 142356 338056
rect 142292 337996 142356 338000
rect 121684 337860 121748 337924
rect 197860 333236 197924 333300
rect 70900 332556 70964 332620
rect 122052 331740 122116 331804
rect 124812 331740 124876 331804
rect 133828 331740 133892 331804
rect 128860 331060 128924 331124
rect 326660 331060 326724 331124
rect 69060 324940 69124 325004
rect 71084 322084 71148 322148
rect 178540 320724 178604 320788
rect 321508 318820 321572 318884
rect 128676 318744 128740 318748
rect 128676 318688 128690 318744
rect 128690 318688 128740 318744
rect 128676 318684 128740 318688
rect 125732 309224 125796 309228
rect 125732 309168 125782 309224
rect 125782 309168 125796 309224
rect 125732 309164 125796 309168
rect 69244 307804 69308 307868
rect 71084 302228 71148 302292
rect 123340 292572 123404 292636
rect 70532 289444 70596 289508
rect 128860 288356 128924 288420
rect 70532 284004 70596 284068
rect 69060 276252 69124 276316
rect 69244 269452 69308 269516
rect 123340 267004 123404 267068
rect 133092 256668 133156 256732
rect 128860 255852 128924 255916
rect 197124 252452 197188 252516
rect 192340 251228 192404 251292
rect 119292 247692 119356 247756
rect 70164 246332 70228 246396
rect 120028 245244 120092 245308
rect 140820 242796 140884 242860
rect 70532 242388 70596 242452
rect 196572 242116 196636 242180
rect 70532 241572 70596 241636
rect 120028 241164 120092 241228
rect 70348 240892 70412 240956
rect 69060 240212 69124 240276
rect 320036 240348 320100 240412
rect 200620 240212 200684 240276
rect 70164 239804 70228 239868
rect 124812 239668 124876 239732
rect 70348 238580 70412 238644
rect 129780 238580 129844 238644
rect 320036 238444 320100 238508
rect 71084 237220 71148 237284
rect 125732 237084 125796 237148
rect 321508 236540 321572 236604
rect 196572 235996 196636 236060
rect 57836 235860 57900 235924
rect 129780 233140 129844 233204
rect 137140 233004 137204 233068
rect 328500 232460 328564 232524
rect 255268 231100 255332 231164
rect 69060 228924 69124 228988
rect 192340 228244 192404 228308
rect 321508 224436 321572 224500
rect 178540 221444 178604 221508
rect 120028 217228 120092 217292
rect 160692 215868 160756 215932
rect 268332 215868 268396 215932
rect 263548 206212 263612 206276
rect 258580 204852 258644 204916
rect 259500 200636 259564 200700
rect 254532 198052 254596 198116
rect 336044 197916 336108 197980
rect 266308 195332 266372 195396
rect 65932 195196 65996 195260
rect 258396 191116 258460 191180
rect 259684 190980 259748 191044
rect 262260 189620 262324 189684
rect 502380 189620 502444 189684
rect 263732 187036 263796 187100
rect 249196 186900 249260 186964
rect 200620 185540 200684 185604
rect 256740 184316 256804 184380
rect 70900 184180 70964 184244
rect 166212 183636 166276 183700
rect 168972 181460 169036 181524
rect 321324 181460 321388 181524
rect 252508 181324 252572 181388
rect 166396 180780 166460 180844
rect 255452 180236 255516 180300
rect 262444 180100 262508 180164
rect 197124 179964 197188 180028
rect 269068 178740 269132 178804
rect 249380 178604 249444 178668
rect 331444 178604 331508 178668
rect 342852 178060 342916 178124
rect 100708 177652 100772 177716
rect 105676 177712 105740 177716
rect 105676 177656 105726 177712
rect 105726 177656 105740 177712
rect 105676 177652 105740 177656
rect 106964 177652 107028 177716
rect 110644 177712 110708 177716
rect 110644 177656 110694 177712
rect 110694 177656 110708 177712
rect 110644 177652 110708 177656
rect 112116 177652 112180 177716
rect 118372 177712 118436 177716
rect 118372 177656 118422 177712
rect 118422 177656 118436 177712
rect 118372 177652 118436 177656
rect 119476 177712 119540 177716
rect 119476 177656 119526 177712
rect 119526 177656 119540 177712
rect 119476 177652 119540 177656
rect 123156 177652 123220 177716
rect 124444 177652 124508 177716
rect 129412 177712 129476 177716
rect 129412 177656 129462 177712
rect 129462 177656 129476 177712
rect 129412 177652 129476 177656
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 494100 177244 494164 177308
rect 97028 176972 97092 177036
rect 115796 177032 115860 177036
rect 115796 176976 115846 177032
rect 115846 176976 115860 177032
rect 115796 176972 115860 176976
rect 125732 176972 125796 177036
rect 134380 176972 134444 177036
rect 114324 176836 114388 176900
rect 214420 176836 214484 176900
rect 98316 176700 98380 176764
rect 104572 176760 104636 176764
rect 104572 176704 104622 176760
rect 104622 176704 104636 176760
rect 104572 176700 104636 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 113220 176700 113284 176764
rect 127020 176760 127084 176764
rect 127020 176704 127070 176760
rect 127070 176704 127084 176760
rect 127020 176700 127084 176704
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 499804 176700 499868 176764
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176488 128188 176492
rect 128124 176432 128174 176488
rect 128174 176432 128188 176488
rect 128124 176428 128188 176432
rect 321692 176156 321756 176220
rect 320220 175748 320284 175812
rect 101996 175400 102060 175404
rect 101996 175344 102046 175400
rect 102046 175344 102060 175400
rect 101996 175340 102060 175344
rect 116900 175400 116964 175404
rect 116900 175344 116950 175400
rect 116950 175344 116964 175400
rect 116900 175340 116964 175344
rect 120764 175400 120828 175404
rect 120764 175344 120814 175400
rect 120814 175344 120828 175400
rect 120764 175340 120828 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 130700 175400 130764 175404
rect 130700 175344 130750 175400
rect 130750 175344 130764 175400
rect 130700 175340 130764 175344
rect 332916 175204 332980 175268
rect 249380 174660 249444 174724
rect 496860 174388 496924 174452
rect 249196 174252 249260 174316
rect 332916 172484 332980 172548
rect 334756 171124 334820 171188
rect 494468 171396 494532 171460
rect 256740 170852 256804 170916
rect 321324 170580 321388 170644
rect 335860 169764 335924 169828
rect 214420 164732 214484 164796
rect 263732 163100 263796 163164
rect 340276 162828 340340 162892
rect 258396 160924 258460 160988
rect 166396 158748 166460 158812
rect 338620 158748 338684 158812
rect 166212 156028 166276 156092
rect 255268 156300 255332 156364
rect 321692 155212 321756 155276
rect 262444 154532 262508 154596
rect 251772 149636 251836 149700
rect 326660 149636 326724 149700
rect 340092 148276 340156 148340
rect 269068 148004 269132 148068
rect 254532 146508 254596 146572
rect 168972 144876 169036 144940
rect 259500 145012 259564 145076
rect 252508 144604 252572 144668
rect 336044 144740 336108 144804
rect 331444 144060 331508 144124
rect 266308 142156 266372 142220
rect 306972 141204 307036 141268
rect 255452 141068 255516 141132
rect 259684 140932 259748 140996
rect 263548 140796 263612 140860
rect 330340 139436 330404 139500
rect 327028 139300 327092 139364
rect 253612 138348 253676 138412
rect 262260 138212 262324 138276
rect 170444 136716 170508 136780
rect 170260 136036 170324 136100
rect 169156 135220 169220 135284
rect 257292 134132 257356 134196
rect 166396 132772 166460 132836
rect 170260 132636 170324 132700
rect 331260 131140 331324 131204
rect 321508 131004 321572 131068
rect 305500 129780 305564 129844
rect 172100 128556 172164 128620
rect 168236 128420 168300 128484
rect 255820 128692 255884 128756
rect 307156 127604 307220 127668
rect 166212 127060 166276 127124
rect 328500 125564 328564 125628
rect 251956 123252 252020 123316
rect 251772 122980 251836 123044
rect 306972 119308 307036 119372
rect 334572 117268 334636 117332
rect 249564 114820 249628 114884
rect 302740 114276 302804 114340
rect 345612 113188 345676 113252
rect 502380 110468 502444 110532
rect 321508 109516 321572 109580
rect 214604 105164 214668 105228
rect 214420 103532 214484 103596
rect 493916 102172 493980 102236
rect 173940 101356 174004 101420
rect 304212 101084 304276 101148
rect 494468 98636 494532 98700
rect 324268 98500 324332 98564
rect 249380 98364 249444 98428
rect 251956 97004 252020 97068
rect 306972 97004 307036 97068
rect 493916 96460 493980 96524
rect 321508 95100 321572 95164
rect 85534 94752 85598 94756
rect 85534 94696 85578 94752
rect 85578 94696 85598 94752
rect 85534 94692 85598 94696
rect 112326 94752 112390 94756
rect 112326 94696 112350 94752
rect 112350 94696 112390 94752
rect 112326 94692 112390 94696
rect 122798 94752 122862 94756
rect 122798 94696 122838 94752
rect 122838 94696 122862 94752
rect 122798 94692 122862 94696
rect 124430 94692 124494 94756
rect 151492 94692 151556 94756
rect 151766 94692 151830 94756
rect 214604 93740 214668 93804
rect 151676 93664 151740 93668
rect 151676 93608 151726 93664
rect 151726 93608 151740 93664
rect 151676 93604 151740 93608
rect 324268 93604 324332 93668
rect 123156 93528 123220 93532
rect 123156 93472 123206 93528
rect 123206 93472 123220 93528
rect 123156 93468 123220 93472
rect 100524 93256 100588 93260
rect 100524 93200 100574 93256
rect 100574 93200 100588 93256
rect 100524 93196 100588 93200
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 84332 92380 84396 92444
rect 86724 92440 86788 92444
rect 86724 92384 86774 92440
rect 86774 92384 86788 92440
rect 86724 92380 86788 92384
rect 88012 92440 88076 92444
rect 88012 92384 88062 92440
rect 88062 92384 88076 92440
rect 88012 92380 88076 92384
rect 99972 92380 100036 92444
rect 101996 92440 102060 92444
rect 101996 92384 102010 92440
rect 102010 92384 102060 92440
rect 101996 92380 102060 92384
rect 102732 92380 102796 92444
rect 104388 92440 104452 92444
rect 104388 92384 104438 92440
rect 104438 92384 104452 92440
rect 104388 92380 104452 92384
rect 105676 92440 105740 92444
rect 105676 92384 105726 92440
rect 105726 92384 105740 92440
rect 105676 92380 105740 92384
rect 106596 92380 106660 92444
rect 107700 92380 107764 92444
rect 108068 92380 108132 92444
rect 109172 92380 109236 92444
rect 110644 92440 110708 92444
rect 110644 92384 110694 92440
rect 110694 92384 110708 92440
rect 110644 92380 110708 92384
rect 113220 92380 113284 92444
rect 119292 92440 119356 92444
rect 119292 92384 119342 92440
rect 119342 92384 119356 92440
rect 119292 92380 119356 92384
rect 119660 92380 119724 92444
rect 129412 92440 129476 92444
rect 129412 92384 129462 92440
rect 129462 92384 129476 92440
rect 129412 92380 129476 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 100708 92244 100772 92308
rect 102548 92244 102612 92308
rect 104572 92304 104636 92308
rect 104572 92248 104622 92304
rect 104622 92248 104636 92304
rect 104572 92244 104636 92248
rect 105492 92244 105556 92308
rect 106412 92244 106476 92308
rect 116716 92244 116780 92308
rect 101812 92108 101876 92172
rect 117084 92168 117148 92172
rect 117084 92112 117134 92168
rect 117134 92112 117148 92168
rect 117084 92108 117148 92112
rect 88932 91760 88996 91764
rect 88932 91704 88982 91760
rect 88982 91704 88996 91760
rect 88932 91700 88996 91704
rect 111196 91700 111260 91764
rect 114508 91700 114572 91764
rect 118004 91624 118068 91628
rect 118004 91568 118054 91624
rect 118054 91568 118068 91624
rect 118004 91564 118068 91568
rect 120580 91564 120644 91628
rect 134380 91700 134444 91764
rect 97212 91428 97276 91492
rect 98132 91428 98196 91492
rect 93900 91292 93964 91356
rect 98500 91292 98564 91356
rect 115796 91352 115860 91356
rect 115796 91296 115810 91352
rect 115810 91296 115860 91352
rect 115796 91292 115860 91296
rect 122052 91352 122116 91356
rect 122052 91296 122102 91352
rect 122102 91296 122116 91352
rect 122052 91292 122116 91296
rect 126652 91352 126716 91356
rect 126652 91296 126702 91352
rect 126702 91296 126716 91352
rect 126652 91292 126716 91296
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96292 91156 96356 91220
rect 96660 91156 96724 91220
rect 99052 91216 99116 91220
rect 99052 91160 99102 91216
rect 99102 91160 99116 91216
rect 99052 91156 99116 91160
rect 109540 91156 109604 91220
rect 111932 91156 111996 91220
rect 114324 91216 114388 91220
rect 114324 91160 114374 91216
rect 114374 91160 114388 91216
rect 114324 91156 114388 91160
rect 114876 91156 114940 91220
rect 115428 91156 115492 91220
rect 118188 91156 118252 91220
rect 120212 91156 120276 91220
rect 121684 91156 121748 91220
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 125364 91156 125428 91220
rect 125732 91156 125796 91220
rect 126468 91156 126532 91220
rect 127572 91156 127636 91220
rect 130700 91156 130764 91220
rect 151308 91156 151372 91220
rect 214420 91020 214484 91084
rect 132356 90884 132420 90948
rect 168972 90884 169036 90948
rect 191236 87484 191300 87548
rect 334756 87484 334820 87548
rect 166396 86804 166460 86868
rect 193812 86124 193876 86188
rect 342852 84900 342916 84964
rect 307156 84764 307220 84828
rect 169156 84084 169220 84148
rect 173020 83404 173084 83468
rect 340276 83404 340340 83468
rect 170444 82724 170508 82788
rect 195100 82044 195164 82108
rect 172100 81364 172164 81428
rect 332916 80684 332980 80748
rect 166212 80004 166276 80068
rect 335860 79324 335924 79388
rect 168236 78508 168300 78572
rect 338252 78508 338316 78572
rect 170260 78372 170324 78436
rect 300716 76468 300780 76532
rect 258580 67492 258644 67556
rect 61700 62868 61764 62932
rect 62988 62732 63052 62796
rect 66116 59876 66180 59940
rect 257292 51716 257356 51780
rect 189948 46140 190012 46204
rect 340828 46200 340892 46204
rect 340828 46144 340878 46200
rect 340878 46144 340892 46200
rect 340828 46140 340892 46144
rect 338620 45460 338684 45524
rect 186820 43420 186884 43484
rect 64460 42196 64524 42260
rect 304212 42060 304276 42124
rect 184060 40564 184124 40628
rect 300716 39536 300780 39540
rect 300716 39480 300730 39536
rect 300730 39480 300780 39536
rect 300716 39476 300780 39480
rect 253060 37844 253124 37908
rect 268332 35124 268396 35188
rect 191052 28188 191116 28252
rect 58940 26148 59004 26212
rect 61884 19892 61948 19956
rect 306972 18532 307036 18596
rect 305500 17172 305564 17236
rect 494100 15132 494164 15196
rect 255820 14452 255884 14516
rect 340828 11732 340892 11796
rect 249196 11596 249260 11660
rect 249380 10236 249444 10300
rect 499804 8196 499868 8260
rect 188292 6836 188356 6900
rect 302740 4796 302804 4860
rect 496860 3980 496924 4044
rect 173940 3300 174004 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 39803 582452 39869 582453
rect 39803 582388 39804 582452
rect 39868 582388 39869 582452
rect 39803 582387 39869 582388
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 39806 485757 39866 582387
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 44035 526420 44101 526421
rect 44035 526356 44036 526420
rect 44100 526356 44101 526420
rect 44035 526355 44101 526356
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 39803 485756 39869 485757
rect 39803 485692 39804 485756
rect 39868 485692 39869 485756
rect 39803 485691 39869 485692
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 44038 438701 44098 526355
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 44035 438700 44101 438701
rect 44035 438636 44036 438700
rect 44100 438636 44101 438700
rect 44035 438635 44101 438636
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 52315 583948 52381 583949
rect 52315 583884 52316 583948
rect 52380 583884 52381 583948
rect 52315 583883 52381 583884
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 52318 493373 52378 583883
rect 55075 571980 55141 571981
rect 55075 571916 55076 571980
rect 55140 571916 55141 571980
rect 55075 571915 55141 571916
rect 50843 493372 50909 493373
rect 50843 493308 50844 493372
rect 50908 493308 50909 493372
rect 50843 493307 50909 493308
rect 52315 493372 52381 493373
rect 52315 493308 52316 493372
rect 52380 493308 52381 493372
rect 52315 493307 52381 493308
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 50846 387701 50906 493307
rect 53603 489156 53669 489157
rect 53603 489092 53604 489156
rect 53668 489092 53669 489156
rect 53603 489091 53669 489092
rect 52315 487252 52381 487253
rect 52315 487188 52316 487252
rect 52380 487188 52381 487252
rect 52315 487187 52381 487188
rect 52318 390693 52378 487187
rect 53606 435845 53666 489091
rect 55078 473245 55138 571915
rect 55794 561454 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 62987 570212 63053 570213
rect 62987 570148 62988 570212
rect 63052 570148 63053 570212
rect 62987 570147 63053 570148
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59123 563276 59189 563277
rect 59123 563212 59124 563276
rect 59188 563212 59189 563276
rect 59123 563211 59189 563212
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 57835 490516 57901 490517
rect 57835 490452 57836 490516
rect 57900 490452 57901 490516
rect 57835 490451 57901 490452
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55075 473244 55141 473245
rect 55075 473180 55076 473244
rect 55140 473180 55141 473244
rect 55075 473179 55141 473180
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 53603 435844 53669 435845
rect 53603 435780 53604 435844
rect 53668 435780 53669 435844
rect 53603 435779 53669 435780
rect 55794 417454 56414 452898
rect 57838 434621 57898 490451
rect 59126 463861 59186 563211
rect 59514 529174 60134 564618
rect 61883 549540 61949 549541
rect 61883 549476 61884 549540
rect 61948 549476 61949 549540
rect 61883 549475 61949 549476
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59123 463860 59189 463861
rect 59123 463796 59124 463860
rect 59188 463796 59189 463860
rect 59123 463795 59189 463796
rect 57835 434620 57901 434621
rect 57835 434556 57836 434620
rect 57900 434556 57901 434620
rect 57835 434555 57901 434556
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 53787 395996 53853 395997
rect 53787 395932 53788 395996
rect 53852 395932 53853 395996
rect 53787 395931 53853 395932
rect 52315 390692 52381 390693
rect 52315 390628 52316 390692
rect 52380 390628 52381 390692
rect 52315 390627 52381 390628
rect 50843 387700 50909 387701
rect 50843 387636 50844 387700
rect 50908 387636 50909 387700
rect 50843 387635 50909 387636
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 53790 355469 53850 395931
rect 55794 381454 56414 416898
rect 57835 389196 57901 389197
rect 57835 389132 57836 389196
rect 57900 389132 57901 389196
rect 57835 389131 57901 389132
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 53787 355468 53853 355469
rect 53787 355404 53788 355468
rect 53852 355404 53853 355468
rect 53787 355403 53853 355404
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 57838 235925 57898 389131
rect 58939 386340 59005 386341
rect 58939 386276 58940 386340
rect 59004 386276 59005 386340
rect 58939 386275 59005 386276
rect 57835 235924 57901 235925
rect 57835 235860 57836 235924
rect 57900 235860 57901 235924
rect 57835 235859 57901 235860
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 58942 26213 59002 386275
rect 59126 368389 59186 463795
rect 59514 457174 60134 492618
rect 61699 471340 61765 471341
rect 61699 471276 61700 471340
rect 61764 471276 61765 471340
rect 61699 471275 61765 471276
rect 60595 463588 60661 463589
rect 60595 463524 60596 463588
rect 60660 463524 60661 463588
rect 60595 463523 60661 463524
rect 60598 462909 60658 463523
rect 60595 462908 60661 462909
rect 60595 462844 60596 462908
rect 60660 462844 60661 462908
rect 60595 462843 60661 462844
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59123 368388 59189 368389
rect 59123 368324 59124 368388
rect 59188 368324 59189 368388
rect 59123 368323 59189 368324
rect 59514 349174 60134 384618
rect 60598 367029 60658 462843
rect 61702 383670 61762 471275
rect 61886 449853 61946 549475
rect 62990 471613 63050 570147
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66115 577828 66181 577829
rect 66115 577764 66116 577828
rect 66180 577764 66181 577828
rect 66115 577763 66181 577764
rect 64643 575108 64709 575109
rect 64643 575044 64644 575108
rect 64708 575044 64709 575108
rect 64643 575043 64709 575044
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 62987 471612 63053 471613
rect 62987 471548 62988 471612
rect 63052 471548 63053 471612
rect 62987 471547 63053 471548
rect 62990 471341 63050 471547
rect 62987 471340 63053 471341
rect 62987 471276 62988 471340
rect 63052 471276 63053 471340
rect 62987 471275 63053 471276
rect 62987 467940 63053 467941
rect 62987 467876 62988 467940
rect 63052 467876 63053 467940
rect 62987 467875 63053 467876
rect 61883 449852 61949 449853
rect 61883 449788 61884 449852
rect 61948 449788 61949 449852
rect 61883 449787 61949 449788
rect 61886 448629 61946 449787
rect 61883 448628 61949 448629
rect 61883 448564 61884 448628
rect 61948 448564 61949 448628
rect 61883 448563 61949 448564
rect 61883 445772 61949 445773
rect 61883 445708 61884 445772
rect 61948 445708 61949 445772
rect 61883 445707 61949 445708
rect 61518 383610 61762 383670
rect 61518 381037 61578 383610
rect 61699 382260 61765 382261
rect 61699 382196 61700 382260
rect 61764 382196 61765 382260
rect 61699 382195 61765 382196
rect 61515 381036 61581 381037
rect 61515 380972 61516 381036
rect 61580 380972 61581 381036
rect 61515 380971 61581 380972
rect 60595 367028 60661 367029
rect 60595 366964 60596 367028
rect 60660 366964 60661 367028
rect 60595 366963 60661 366964
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 61702 62933 61762 382195
rect 61886 346629 61946 445707
rect 62990 371381 63050 467875
rect 63234 460894 63854 496338
rect 64646 477461 64706 575043
rect 65931 484668 65997 484669
rect 65931 484604 65932 484668
rect 65996 484604 65997 484668
rect 65931 484603 65997 484604
rect 64643 477460 64709 477461
rect 64643 477396 64644 477460
rect 64708 477396 64709 477460
rect 64643 477395 64709 477396
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 64643 447812 64709 447813
rect 64643 447748 64644 447812
rect 64708 447748 64709 447812
rect 64643 447747 64709 447748
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 62987 371380 63053 371381
rect 62987 371316 62988 371380
rect 63052 371316 63053 371380
rect 62987 371315 63053 371316
rect 62987 367028 63053 367029
rect 62987 366964 62988 367028
rect 63052 366964 63053 367028
rect 62987 366963 63053 366964
rect 62990 365805 63050 366963
rect 62987 365804 63053 365805
rect 62987 365740 62988 365804
rect 63052 365740 63053 365804
rect 62987 365739 63053 365740
rect 61883 346628 61949 346629
rect 61883 346564 61884 346628
rect 61948 346564 61949 346628
rect 61883 346563 61949 346564
rect 61699 62932 61765 62933
rect 61699 62868 61700 62932
rect 61764 62868 61765 62932
rect 61699 62867 61765 62868
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 58939 26212 59005 26213
rect 58939 26148 58940 26212
rect 59004 26148 59005 26212
rect 58939 26147 59005 26148
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 61886 19957 61946 346563
rect 62990 62797 63050 365739
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 64459 349892 64525 349893
rect 64459 349828 64460 349892
rect 64524 349828 64525 349892
rect 64459 349827 64525 349828
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 62987 62796 63053 62797
rect 62987 62732 62988 62796
rect 63052 62732 63053 62796
rect 62987 62731 63053 62732
rect 63234 28894 63854 64338
rect 64462 42261 64522 349827
rect 64646 349757 64706 447747
rect 65934 436797 65994 484603
rect 66118 478957 66178 577763
rect 66954 572614 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 584000 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 584000 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 584000 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 584000 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 584000 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 584000 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 584000 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 584000 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 69795 581364 69861 581365
rect 69795 581300 69796 581364
rect 69860 581300 69861 581364
rect 69795 581299 69861 581300
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 68875 554028 68941 554029
rect 68875 553964 68876 554028
rect 68940 553964 68941 554028
rect 68875 553963 68941 553964
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66115 478956 66181 478957
rect 66115 478892 66116 478956
rect 66180 478892 66181 478956
rect 66115 478891 66181 478892
rect 66115 474332 66181 474333
rect 66115 474268 66116 474332
rect 66180 474268 66181 474332
rect 66115 474267 66181 474268
rect 65931 436796 65997 436797
rect 65931 436732 65932 436796
rect 65996 436732 65997 436796
rect 65931 436731 65997 436732
rect 66118 379677 66178 474267
rect 66954 464614 67574 500058
rect 68691 477052 68757 477053
rect 68691 476988 68692 477052
rect 68756 476988 68757 477052
rect 68691 476987 68757 476988
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 68507 454068 68573 454069
rect 68507 454004 68508 454068
rect 68572 454004 68573 454068
rect 68507 454003 68573 454004
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 68510 393330 68570 454003
rect 68694 401437 68754 476987
rect 68878 454069 68938 553963
rect 69611 536892 69677 536893
rect 69611 536828 69612 536892
rect 69676 536828 69677 536892
rect 69611 536827 69677 536828
rect 69059 486708 69125 486709
rect 69059 486644 69060 486708
rect 69124 486644 69125 486708
rect 69059 486643 69125 486644
rect 68875 454068 68941 454069
rect 68875 454004 68876 454068
rect 68940 454004 68941 454068
rect 68875 454003 68941 454004
rect 69062 435301 69122 486643
rect 69614 440741 69674 536827
rect 69798 485893 69858 581299
rect 76576 579454 76896 579486
rect 76576 579218 76618 579454
rect 76854 579218 76896 579454
rect 76576 579134 76896 579218
rect 76576 578898 76618 579134
rect 76854 578898 76896 579134
rect 76576 578866 76896 578898
rect 87840 579454 88160 579486
rect 87840 579218 87882 579454
rect 88118 579218 88160 579454
rect 87840 579134 88160 579218
rect 87840 578898 87882 579134
rect 88118 578898 88160 579134
rect 87840 578866 88160 578898
rect 99104 579454 99424 579486
rect 99104 579218 99146 579454
rect 99382 579218 99424 579454
rect 99104 579134 99424 579218
rect 99104 578898 99146 579134
rect 99382 578898 99424 579134
rect 99104 578866 99424 578898
rect 109794 579454 110414 614898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 115979 585172 116045 585173
rect 115979 585108 115980 585172
rect 116044 585108 116045 585172
rect 115979 585107 116045 585108
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111747 582588 111813 582589
rect 111747 582524 111748 582588
rect 111812 582524 111813 582588
rect 111747 582523 111813 582524
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 107699 578780 107765 578781
rect 107699 578716 107700 578780
rect 107764 578716 107765 578780
rect 107699 578715 107765 578716
rect 105491 563004 105557 563005
rect 105491 562940 105492 563004
rect 105556 562940 105557 563004
rect 105491 562939 105557 562940
rect 82208 561454 82528 561486
rect 82208 561218 82250 561454
rect 82486 561218 82528 561454
rect 82208 561134 82528 561218
rect 82208 560898 82250 561134
rect 82486 560898 82528 561134
rect 82208 560866 82528 560898
rect 93472 561454 93792 561486
rect 93472 561218 93514 561454
rect 93750 561218 93792 561454
rect 93472 561134 93792 561218
rect 93472 560898 93514 561134
rect 93750 560898 93792 561134
rect 93472 560866 93792 560898
rect 69979 557428 70045 557429
rect 69979 557364 69980 557428
rect 70044 557364 70045 557428
rect 69979 557363 70045 557364
rect 69982 557290 70042 557363
rect 69982 557230 70410 557290
rect 69795 485892 69861 485893
rect 69795 485828 69796 485892
rect 69860 485828 69861 485892
rect 69795 485827 69861 485828
rect 70350 484669 70410 557230
rect 105494 547890 105554 562939
rect 106411 556340 106477 556341
rect 106411 556276 106412 556340
rect 106476 556276 106477 556340
rect 106411 556275 106477 556276
rect 104942 547830 105554 547890
rect 76576 543454 76896 543486
rect 76576 543218 76618 543454
rect 76854 543218 76896 543454
rect 76576 543134 76896 543218
rect 76576 542898 76618 543134
rect 76854 542898 76896 543134
rect 76576 542866 76896 542898
rect 87840 543454 88160 543486
rect 87840 543218 87882 543454
rect 88118 543218 88160 543454
rect 87840 543134 88160 543218
rect 87840 542898 87882 543134
rect 88118 542898 88160 543134
rect 87840 542866 88160 542898
rect 99104 543454 99424 543486
rect 99104 543218 99146 543454
rect 99382 543218 99424 543454
rect 99104 543134 99424 543218
rect 99104 542898 99146 543134
rect 99382 542898 99424 543134
rect 99104 542866 99424 542898
rect 73794 507454 74414 538000
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 492000 74414 506898
rect 77514 511174 78134 538000
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 492000 78134 510618
rect 81234 514894 81854 538000
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 492000 81854 514338
rect 84954 518614 85574 538000
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 492000 85574 518058
rect 91794 525454 92414 538000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 492000 92414 524898
rect 95514 529174 96134 538000
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 492000 96134 492618
rect 99234 532894 99854 538000
rect 101259 536892 101325 536893
rect 101259 536828 101260 536892
rect 101324 536828 101325 536892
rect 101259 536827 101325 536828
rect 101995 536892 102061 536893
rect 101995 536828 101996 536892
rect 102060 536828 102061 536892
rect 101995 536827 102061 536828
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 492000 99854 496338
rect 99235 491740 99301 491741
rect 99235 491676 99236 491740
rect 99300 491676 99301 491740
rect 99235 491675 99301 491676
rect 70347 484668 70413 484669
rect 70347 484604 70348 484668
rect 70412 484604 70413 484668
rect 70347 484603 70413 484604
rect 99238 484530 99298 491675
rect 99419 484532 99485 484533
rect 99419 484530 99420 484532
rect 99238 484470 99420 484530
rect 99419 484468 99420 484470
rect 99484 484468 99485 484532
rect 99419 484467 99485 484468
rect 75576 471454 75896 471486
rect 75576 471218 75618 471454
rect 75854 471218 75896 471454
rect 75576 471134 75896 471218
rect 75576 470898 75618 471134
rect 75854 470898 75896 471134
rect 75576 470866 75896 470898
rect 84840 471454 85160 471486
rect 84840 471218 84882 471454
rect 85118 471218 85160 471454
rect 84840 471134 85160 471218
rect 84840 470898 84882 471134
rect 85118 470898 85160 471134
rect 84840 470866 85160 470898
rect 94104 471454 94424 471486
rect 94104 471218 94146 471454
rect 94382 471218 94424 471454
rect 94104 471134 94424 471218
rect 94104 470898 94146 471134
rect 94382 470898 94424 471134
rect 94104 470866 94424 470898
rect 80208 453454 80528 453486
rect 80208 453218 80250 453454
rect 80486 453218 80528 453454
rect 80208 453134 80528 453218
rect 80208 452898 80250 453134
rect 80486 452898 80528 453134
rect 80208 452866 80528 452898
rect 89472 453454 89792 453486
rect 89472 453218 89514 453454
rect 89750 453218 89792 453454
rect 89472 453134 89792 453218
rect 89472 452898 89514 453134
rect 89750 452898 89792 453134
rect 89472 452866 89792 452898
rect 99419 443052 99485 443053
rect 99419 443050 99420 443052
rect 99054 442990 99420 443050
rect 69611 440740 69677 440741
rect 69611 440676 69612 440740
rect 69676 440676 69677 440740
rect 69611 440675 69677 440676
rect 69059 435300 69125 435301
rect 69059 435236 69060 435300
rect 69124 435236 69125 435300
rect 69059 435235 69125 435236
rect 68691 401436 68757 401437
rect 68691 401372 68692 401436
rect 68756 401372 68757 401436
rect 68691 401371 68757 401372
rect 68875 400348 68941 400349
rect 68875 400284 68876 400348
rect 68940 400284 68941 400348
rect 68875 400283 68941 400284
rect 68878 396269 68938 400283
rect 68875 396268 68941 396269
rect 68875 396204 68876 396268
rect 68940 396204 68941 396268
rect 68875 396203 68941 396204
rect 68510 393270 68754 393330
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66115 379676 66181 379677
rect 66115 379612 66116 379676
rect 66180 379612 66181 379676
rect 66115 379611 66181 379612
rect 65931 371924 65997 371925
rect 65931 371860 65932 371924
rect 65996 371860 65997 371924
rect 65931 371859 65997 371860
rect 64643 349756 64709 349757
rect 64643 349692 64644 349756
rect 64708 349692 64709 349756
rect 64643 349691 64709 349692
rect 65934 195261 65994 371859
rect 66115 365668 66181 365669
rect 66115 365604 66116 365668
rect 66180 365604 66181 365668
rect 66115 365603 66181 365604
rect 66118 364717 66178 365603
rect 66115 364716 66181 364717
rect 66115 364652 66116 364716
rect 66180 364652 66181 364716
rect 66115 364651 66181 364652
rect 65931 195260 65997 195261
rect 65931 195196 65932 195260
rect 65996 195196 65997 195260
rect 65931 195195 65997 195196
rect 66118 59941 66178 364651
rect 66954 356614 67574 392058
rect 68694 390693 68754 393270
rect 68691 390692 68757 390693
rect 68691 390628 68692 390692
rect 68756 390628 68757 390692
rect 68691 390627 68757 390628
rect 68694 356965 68754 390627
rect 68691 356964 68757 356965
rect 68691 356900 68692 356964
rect 68756 356900 68757 356964
rect 68691 356899 68757 356900
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 353292 66733 353293
rect 66667 353228 66668 353292
rect 66732 353228 66733 353292
rect 66667 353227 66733 353228
rect 66670 338741 66730 353227
rect 66667 338740 66733 338741
rect 66667 338676 66668 338740
rect 66732 338676 66733 338740
rect 66667 338675 66733 338676
rect 66954 320614 67574 356058
rect 68878 350165 68938 396203
rect 68875 350164 68941 350165
rect 68875 350100 68876 350164
rect 68940 350100 68941 350164
rect 68875 350099 68941 350100
rect 69614 340101 69674 440675
rect 70163 440060 70229 440061
rect 70163 439996 70164 440060
rect 70228 439996 70229 440060
rect 70163 439995 70229 439996
rect 70166 437490 70226 439995
rect 70166 437430 70410 437490
rect 69795 385388 69861 385389
rect 69795 385324 69796 385388
rect 69860 385324 69861 385388
rect 69795 385323 69861 385324
rect 69798 369885 69858 385323
rect 69979 383212 70045 383213
rect 69979 383148 69980 383212
rect 70044 383210 70045 383212
rect 70350 383210 70410 437430
rect 73794 435454 74414 438000
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 388000 74414 398898
rect 77514 403174 78134 438000
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 388000 78134 402618
rect 81234 406894 81854 438000
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 388000 81854 406338
rect 84954 410614 85574 438000
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 388000 85574 410058
rect 91794 417454 92414 438000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 388000 92414 416898
rect 95514 421174 96134 438000
rect 99054 435981 99114 442990
rect 99419 442988 99420 442990
rect 99484 442988 99485 443052
rect 99419 442987 99485 442988
rect 101262 442373 101322 536827
rect 101998 446589 102058 536827
rect 102954 536614 103574 538000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 103835 490652 103901 490653
rect 103835 490650 103836 490652
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 101995 446588 102061 446589
rect 101995 446524 101996 446588
rect 102060 446524 102061 446588
rect 101995 446523 102061 446524
rect 101259 442372 101325 442373
rect 101259 442308 101260 442372
rect 101324 442308 101325 442372
rect 101259 442307 101325 442308
rect 101262 441965 101322 442307
rect 101259 441964 101325 441965
rect 101259 441900 101260 441964
rect 101324 441900 101325 441964
rect 101259 441899 101325 441900
rect 99051 435980 99117 435981
rect 99051 435916 99052 435980
rect 99116 435916 99117 435980
rect 99051 435915 99117 435916
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 388000 96134 420618
rect 99234 424894 99854 438000
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 388000 99854 388338
rect 102954 428614 103574 464058
rect 103654 490590 103836 490650
rect 103654 438970 103714 490590
rect 103835 490588 103836 490590
rect 103900 490588 103901 490652
rect 103835 490587 103901 490588
rect 104942 474741 105002 547830
rect 104939 474740 105005 474741
rect 104939 474676 104940 474740
rect 105004 474676 105005 474740
rect 104939 474675 105005 474676
rect 105491 474740 105557 474741
rect 105491 474676 105492 474740
rect 105556 474676 105557 474740
rect 105491 474675 105557 474676
rect 103835 438972 103901 438973
rect 103835 438970 103836 438972
rect 103654 438910 103836 438970
rect 103835 438908 103836 438910
rect 103900 438908 103901 438972
rect 103835 438907 103901 438908
rect 105494 437341 105554 474675
rect 106414 464269 106474 556275
rect 107702 537437 107762 578715
rect 109794 543454 110414 578898
rect 110643 577556 110709 577557
rect 110643 577492 110644 577556
rect 110708 577492 110709 577556
rect 110643 577491 110709 577492
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 107883 542740 107949 542741
rect 107883 542676 107884 542740
rect 107948 542676 107949 542740
rect 107883 542675 107949 542676
rect 107699 537436 107765 537437
rect 107699 537372 107700 537436
rect 107764 537372 107765 537436
rect 107699 537371 107765 537372
rect 106411 464268 106477 464269
rect 106411 464204 106412 464268
rect 106476 464204 106477 464268
rect 106411 464203 106477 464204
rect 106779 462908 106845 462909
rect 106779 462844 106780 462908
rect 106844 462844 106845 462908
rect 106779 462843 106845 462844
rect 106782 439109 106842 462843
rect 107886 451349 107946 542675
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 108987 490516 109053 490517
rect 108987 490452 108988 490516
rect 109052 490452 109053 490516
rect 108987 490451 109053 490452
rect 108990 485790 109050 490451
rect 108806 485730 109050 485790
rect 108806 476130 108866 485730
rect 108806 476070 109050 476130
rect 107883 451348 107949 451349
rect 107883 451284 107884 451348
rect 107948 451284 107949 451348
rect 107883 451283 107949 451284
rect 106779 439108 106845 439109
rect 106779 439044 106780 439108
rect 106844 439044 106845 439108
rect 106779 439043 106845 439044
rect 105491 437340 105557 437341
rect 105491 437276 105492 437340
rect 105556 437276 105557 437340
rect 105491 437275 105557 437276
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 388000 103574 392058
rect 108990 388925 109050 476070
rect 109794 471454 110414 506898
rect 110646 486437 110706 577491
rect 110827 529140 110893 529141
rect 110827 529076 110828 529140
rect 110892 529076 110893 529140
rect 110827 529075 110893 529076
rect 110643 486436 110709 486437
rect 110643 486372 110644 486436
rect 110708 486372 110709 486436
rect 110643 486371 110709 486372
rect 110830 474741 110890 529075
rect 111750 496093 111810 582523
rect 113514 547174 114134 582618
rect 114507 573204 114573 573205
rect 114507 573140 114508 573204
rect 114572 573140 114573 573204
rect 114507 573139 114573 573140
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111747 496092 111813 496093
rect 111747 496028 111748 496092
rect 111812 496028 111813 496092
rect 111747 496027 111813 496028
rect 111747 492828 111813 492829
rect 111747 492764 111748 492828
rect 111812 492764 111813 492828
rect 111747 492763 111813 492764
rect 110827 474740 110893 474741
rect 110827 474676 110828 474740
rect 110892 474676 110893 474740
rect 110827 474675 110893 474676
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 111750 459645 111810 492763
rect 113035 485076 113101 485077
rect 113035 485012 113036 485076
rect 113100 485012 113101 485076
rect 113035 485011 113101 485012
rect 113038 480861 113098 485011
rect 113035 480860 113101 480861
rect 113035 480796 113036 480860
rect 113100 480796 113101 480860
rect 113035 480795 113101 480796
rect 113514 475174 114134 510618
rect 114510 482357 114570 573139
rect 115982 534717 116042 585107
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 115979 534716 116045 534717
rect 115979 534652 115980 534716
rect 116044 534652 116045 534716
rect 115979 534651 116045 534652
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 115979 497452 116045 497453
rect 115979 497388 115980 497452
rect 116044 497388 116045 497452
rect 115979 497387 116045 497388
rect 114507 482356 114573 482357
rect 114507 482292 114508 482356
rect 114572 482292 114573 482356
rect 114507 482291 114573 482292
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 459644 111813 459645
rect 111747 459580 111748 459644
rect 111812 459580 111813 459644
rect 111747 459579 111813 459580
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 108987 388924 109053 388925
rect 108987 388860 108988 388924
rect 109052 388860 109053 388924
rect 108987 388859 109053 388860
rect 109794 388000 110414 398898
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 114510 402990 114570 482291
rect 115982 437477 116042 497387
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 115979 437476 116045 437477
rect 115979 437412 115980 437476
rect 116044 437412 116045 437476
rect 115979 437411 116045 437412
rect 117234 406894 117854 442338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 124259 582452 124325 582453
rect 124259 582388 124260 582452
rect 124324 582388 124325 582452
rect 124259 582387 124325 582388
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 124262 491877 124322 582387
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 124259 491876 124325 491877
rect 124259 491812 124260 491876
rect 124324 491812 124325 491876
rect 124259 491811 124325 491812
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 122051 486436 122117 486437
rect 122051 486372 122052 486436
rect 122116 486372 122117 486436
rect 122051 486371 122117 486372
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120027 407828 120093 407829
rect 120027 407764 120028 407828
rect 120092 407764 120093 407828
rect 120027 407763 120093 407764
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 114510 402930 115490 402990
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 388000 114134 402618
rect 114691 392596 114757 392597
rect 114691 392532 114692 392596
rect 114756 392532 114757 392596
rect 114691 392531 114757 392532
rect 70044 383150 70410 383210
rect 70044 383148 70045 383150
rect 69979 383147 70045 383148
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 114694 376410 114754 392531
rect 115430 377365 115490 402930
rect 115979 389876 116045 389877
rect 115979 389812 115980 389876
rect 116044 389812 116045 389876
rect 115979 389811 116045 389812
rect 115982 378589 116042 389811
rect 117234 388000 117854 406338
rect 118003 399668 118069 399669
rect 118003 399604 118004 399668
rect 118068 399604 118069 399668
rect 118003 399603 118069 399604
rect 115979 378588 116045 378589
rect 115979 378524 115980 378588
rect 116044 378524 116045 378588
rect 115979 378523 116045 378524
rect 115427 377364 115493 377365
rect 115427 377300 115428 377364
rect 115492 377300 115493 377364
rect 115427 377299 115493 377300
rect 115427 376412 115493 376413
rect 115427 376410 115428 376412
rect 114694 376350 115428 376410
rect 115427 376348 115428 376350
rect 115492 376348 115493 376412
rect 115427 376347 115493 376348
rect 118006 372741 118066 399603
rect 118739 387700 118805 387701
rect 118739 387636 118740 387700
rect 118804 387636 118805 387700
rect 118739 387635 118805 387636
rect 118742 387021 118802 387635
rect 118739 387020 118805 387021
rect 118739 386956 118740 387020
rect 118804 386956 118805 387020
rect 118739 386955 118805 386956
rect 118003 372740 118069 372741
rect 118003 372676 118004 372740
rect 118068 372676 118069 372740
rect 118003 372675 118069 372676
rect 69795 369884 69861 369885
rect 69795 369820 69796 369884
rect 69860 369820 69861 369884
rect 69795 369819 69861 369820
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 70531 341732 70597 341733
rect 70531 341668 70532 341732
rect 70596 341668 70597 341732
rect 70531 341667 70597 341668
rect 69611 340100 69677 340101
rect 69611 340036 69612 340100
rect 69676 340036 69677 340100
rect 69611 340035 69677 340036
rect 70534 335370 70594 341667
rect 70534 335310 71146 335370
rect 70899 332620 70965 332621
rect 70899 332556 70900 332620
rect 70964 332556 70965 332620
rect 70899 332555 70965 332556
rect 69059 325004 69125 325005
rect 69059 324940 69060 325004
rect 69124 324940 69125 325004
rect 69059 324939 69125 324940
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 69062 276317 69122 324939
rect 69243 307868 69309 307869
rect 69243 307804 69244 307868
rect 69308 307804 69309 307868
rect 69243 307803 69309 307804
rect 69059 276316 69125 276317
rect 69059 276252 69060 276316
rect 69124 276252 69125 276316
rect 69059 276251 69125 276252
rect 69246 269517 69306 307803
rect 70902 296730 70962 332555
rect 71086 322149 71146 335310
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 71083 322148 71149 322149
rect 71083 322084 71084 322148
rect 71148 322084 71149 322148
rect 71083 322083 71149 322084
rect 71083 302292 71149 302293
rect 71083 302228 71084 302292
rect 71148 302228 71149 302292
rect 71083 302227 71149 302228
rect 70534 296670 70962 296730
rect 70534 289509 70594 296670
rect 70531 289508 70597 289509
rect 70531 289444 70532 289508
rect 70596 289444 70597 289508
rect 70531 289443 70597 289444
rect 71086 287070 71146 302227
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 331174 114134 338000
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 334894 117854 338000
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 70534 287010 71146 287070
rect 70534 284069 70594 287010
rect 70531 284068 70597 284069
rect 70531 284004 70532 284068
rect 70596 284004 70597 284068
rect 70531 284003 70597 284004
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 69243 269516 69309 269517
rect 69243 269452 69244 269516
rect 69308 269452 69309 269516
rect 69243 269451 69309 269452
rect 118742 267750 118802 386955
rect 120030 358733 120090 407763
rect 120954 374614 121574 410058
rect 121683 385796 121749 385797
rect 121683 385732 121684 385796
rect 121748 385732 121749 385796
rect 121683 385731 121749 385732
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120027 358732 120093 358733
rect 120027 358668 120028 358732
rect 120092 358668 120093 358732
rect 120027 358667 120093 358668
rect 120027 342140 120093 342141
rect 120027 342076 120028 342140
rect 120092 342076 120093 342140
rect 120027 342075 120093 342076
rect 118742 267690 119354 267750
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 119294 247757 119354 267690
rect 119291 247756 119357 247757
rect 119291 247692 119292 247756
rect 119356 247692 119357 247756
rect 119291 247691 119357 247692
rect 70163 246396 70229 246397
rect 70163 246332 70164 246396
rect 70228 246332 70229 246396
rect 70163 246331 70229 246332
rect 69059 240276 69125 240277
rect 69059 240212 69060 240276
rect 69124 240212 69125 240276
rect 69059 240211 69125 240212
rect 69062 228989 69122 240211
rect 70166 239869 70226 246331
rect 120030 245309 120090 342075
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 121686 337925 121746 385731
rect 122054 380221 122114 486371
rect 124075 483172 124141 483173
rect 124075 483108 124076 483172
rect 124140 483108 124141 483172
rect 124075 483107 124141 483108
rect 122603 405108 122669 405109
rect 122603 405044 122604 405108
rect 122668 405044 122669 405108
rect 122603 405043 122669 405044
rect 122051 380220 122117 380221
rect 122051 380156 122052 380220
rect 122116 380156 122117 380220
rect 122051 380155 122117 380156
rect 122051 376820 122117 376821
rect 122051 376756 122052 376820
rect 122116 376756 122117 376820
rect 122051 376755 122117 376756
rect 121683 337924 121749 337925
rect 121683 337860 121684 337924
rect 121748 337860 121749 337924
rect 121683 337859 121749 337860
rect 122054 331805 122114 376755
rect 122606 338061 122666 405043
rect 124078 378725 124138 483107
rect 126835 453932 126901 453933
rect 126835 453868 126836 453932
rect 126900 453868 126901 453932
rect 126835 453867 126901 453868
rect 124259 398036 124325 398037
rect 124259 397972 124260 398036
rect 124324 397972 124325 398036
rect 124259 397971 124325 397972
rect 124075 378724 124141 378725
rect 124075 378660 124076 378724
rect 124140 378660 124141 378724
rect 124075 378659 124141 378660
rect 124262 339421 124322 397971
rect 126838 343637 126898 453867
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 128675 399532 128741 399533
rect 128675 399530 128676 399532
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 126835 343636 126901 343637
rect 126835 343572 126836 343636
rect 126900 343572 126901 343636
rect 126835 343571 126901 343572
rect 124259 339420 124325 339421
rect 124259 339356 124260 339420
rect 124324 339356 124325 339420
rect 124259 339355 124325 339356
rect 122603 338060 122669 338061
rect 122603 337996 122604 338060
rect 122668 337996 122669 338060
rect 122603 337995 122669 337996
rect 122051 331804 122117 331805
rect 122051 331740 122052 331804
rect 122116 331740 122117 331804
rect 122051 331739 122117 331740
rect 124811 331804 124877 331805
rect 124811 331740 124812 331804
rect 124876 331740 124877 331804
rect 124811 331739 124877 331740
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 123339 292636 123405 292637
rect 123339 292572 123340 292636
rect 123404 292572 123405 292636
rect 123339 292571 123405 292572
rect 123342 267069 123402 292571
rect 123339 267068 123405 267069
rect 123339 267004 123340 267068
rect 123404 267004 123405 267068
rect 123339 267003 123405 267004
rect 120027 245308 120093 245309
rect 120027 245244 120028 245308
rect 120092 245244 120093 245308
rect 120027 245243 120093 245244
rect 70531 242452 70597 242453
rect 70531 242388 70532 242452
rect 70596 242450 70597 242452
rect 70596 242390 71146 242450
rect 70596 242388 70597 242390
rect 70531 242387 70597 242388
rect 70531 241636 70597 241637
rect 70531 241572 70532 241636
rect 70596 241572 70597 241636
rect 70531 241571 70597 241572
rect 70347 240956 70413 240957
rect 70347 240892 70348 240956
rect 70412 240892 70413 240956
rect 70347 240891 70413 240892
rect 70163 239868 70229 239869
rect 70163 239804 70164 239868
rect 70228 239804 70229 239868
rect 70163 239803 70229 239804
rect 70350 238645 70410 240891
rect 70534 238770 70594 241571
rect 70534 238710 70962 238770
rect 70347 238644 70413 238645
rect 70347 238580 70348 238644
rect 70412 238580 70413 238644
rect 70347 238579 70413 238580
rect 69059 228988 69125 228989
rect 69059 228924 69060 228988
rect 69124 228924 69125 228988
rect 69059 228923 69125 228924
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 70902 184245 70962 238710
rect 71086 237285 71146 242390
rect 120027 241228 120093 241229
rect 120027 241164 120028 241228
rect 120092 241164 120093 241228
rect 120027 241163 120093 241164
rect 71083 237284 71149 237285
rect 71083 237220 71084 237284
rect 71148 237220 71149 237284
rect 71083 237219 71149 237220
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 70899 184244 70965 184245
rect 70899 184180 70900 184244
rect 70964 184180 70965 184244
rect 70899 184179 70965 184180
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177036 97093 177037
rect 97027 176972 97028 177036
rect 97092 176972 97093 177036
rect 97027 176971 97093 176972
rect 97030 175130 97090 176971
rect 98315 176764 98381 176765
rect 98315 176700 98316 176764
rect 98380 176700 98381 176764
rect 98315 176699 98381 176700
rect 96960 175070 97090 175130
rect 98318 175130 98378 176699
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177716 100773 177717
rect 100707 177652 100708 177716
rect 100772 177652 100773 177716
rect 100707 177651 100773 177652
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177651
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 106963 177716 107029 177717
rect 106963 177652 106964 177716
rect 107028 177652 107029 177716
rect 106963 177651 107029 177652
rect 104571 176764 104637 176765
rect 104571 176700 104572 176764
rect 104636 176700 104637 176764
rect 104571 176699 104637 176700
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 101995 175404 102061 175405
rect 101995 175340 101996 175404
rect 102060 175340 102061 175404
rect 101995 175339 102061 175340
rect 101998 175130 102058 175339
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 176699
rect 105678 175130 105738 177651
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177651
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 177716 110709 177717
rect 110643 177652 110644 177716
rect 110708 177652 110709 177716
rect 110643 177651 110709 177652
rect 112115 177716 112181 177717
rect 112115 177652 112116 177716
rect 112180 177652 112181 177716
rect 112115 177651 112181 177652
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177651
rect 112118 175130 112178 177651
rect 113219 176764 113285 176765
rect 113219 176700 113220 176764
rect 113284 176700 113285 176764
rect 113219 176699 113285 176700
rect 113222 175130 113282 176699
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 120030 217293 120090 241163
rect 124814 239733 124874 331739
rect 127794 309454 128414 344898
rect 128494 399470 128676 399530
rect 128494 331122 128554 399470
rect 128675 399468 128676 399470
rect 128740 399468 128741 399532
rect 128675 399467 128741 399468
rect 129779 391236 129845 391237
rect 129779 391172 129780 391236
rect 129844 391172 129845 391236
rect 129779 391171 129845 391172
rect 128675 378724 128741 378725
rect 128675 378660 128676 378724
rect 128740 378660 128741 378724
rect 128675 378659 128741 378660
rect 128678 338130 128738 378659
rect 128678 338070 129106 338130
rect 128859 331124 128925 331125
rect 128859 331122 128860 331124
rect 128494 331062 128860 331122
rect 128859 331060 128860 331062
rect 128924 331060 128925 331124
rect 128859 331059 128925 331060
rect 129046 328470 129106 338070
rect 128678 328410 129106 328470
rect 128678 318749 128738 328410
rect 128675 318748 128741 318749
rect 128675 318684 128676 318748
rect 128740 318684 128741 318748
rect 128675 318683 128741 318684
rect 125731 309228 125797 309229
rect 125731 309164 125732 309228
rect 125796 309164 125797 309228
rect 125731 309163 125797 309164
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 124811 239732 124877 239733
rect 124811 239668 124812 239732
rect 124876 239668 124877 239732
rect 124811 239667 124877 239668
rect 120954 230614 121574 238000
rect 125734 237149 125794 309163
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 128859 288420 128925 288421
rect 128859 288356 128860 288420
rect 128924 288356 128925 288420
rect 128859 288355 128925 288356
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 128862 255917 128922 288355
rect 128859 255916 128925 255917
rect 128859 255852 128860 255916
rect 128924 255852 128925 255916
rect 128859 255851 128925 255852
rect 129782 238645 129842 391171
rect 131514 385174 132134 420618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 133827 394908 133893 394909
rect 133827 394844 133828 394908
rect 133892 394844 133893 394908
rect 133827 394843 133893 394844
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 133091 342956 133157 342957
rect 133091 342892 133092 342956
rect 133156 342892 133157 342956
rect 133091 342891 133157 342892
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 133094 256733 133154 342891
rect 133830 331805 133890 394843
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 143579 499628 143645 499629
rect 143579 499564 143580 499628
rect 143644 499564 143645 499628
rect 143579 499563 143645 499564
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 141923 449988 141989 449989
rect 141923 449924 141924 449988
rect 141988 449924 141989 449988
rect 141923 449923 141989 449924
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 140819 380220 140885 380221
rect 140819 380156 140820 380220
rect 140884 380156 140885 380220
rect 140819 380155 140885 380156
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 137139 353972 137205 353973
rect 137139 353908 137140 353972
rect 137204 353908 137205 353972
rect 137139 353907 137205 353908
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 133827 331804 133893 331805
rect 133827 331740 133828 331804
rect 133892 331740 133893 331804
rect 133827 331739 133893 331740
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 133091 256732 133157 256733
rect 133091 256668 133092 256732
rect 133156 256668 133157 256732
rect 133091 256667 133157 256668
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 129779 238644 129845 238645
rect 129779 238580 129780 238644
rect 129844 238580 129845 238644
rect 129779 238579 129845 238580
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 125731 237148 125797 237149
rect 125731 237084 125732 237148
rect 125796 237084 125797 237148
rect 125731 237083 125797 237084
rect 127794 237134 128414 237218
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120027 217292 120093 217293
rect 120027 217228 120028 217292
rect 120092 217228 120093 217292
rect 120027 217227 120093 217228
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 115795 177036 115861 177037
rect 115795 176972 115796 177036
rect 115860 176972 115861 177036
rect 115795 176971 115861 176972
rect 114323 176900 114389 176901
rect 114323 176836 114324 176900
rect 114388 176836 114389 176900
rect 114323 176835 114389 176836
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 176835
rect 115798 175130 115858 176971
rect 117234 176600 117854 190338
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 177716 118437 177717
rect 118371 177652 118372 177716
rect 118436 177652 118437 177716
rect 118371 177651 118437 177652
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 116899 175404 116965 175405
rect 116899 175340 116900 175404
rect 116964 175340 116965 175404
rect 116899 175339 116965 175340
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175339
rect 118374 175130 118434 177651
rect 119478 175130 119538 177651
rect 120954 176600 121574 194058
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 129782 233205 129842 238579
rect 129779 233204 129845 233205
rect 129779 233140 129780 233204
rect 129844 233140 129845 233204
rect 129779 233139 129845 233140
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 123155 177716 123221 177717
rect 123155 177652 123156 177716
rect 123220 177652 123221 177716
rect 123155 177651 123221 177652
rect 124443 177716 124509 177717
rect 124443 177652 124444 177716
rect 124508 177652 124509 177716
rect 124443 177651 124509 177652
rect 120763 175404 120829 175405
rect 120763 175340 120764 175404
rect 120828 175340 120829 175404
rect 120763 175339 120829 175340
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 120766 175130 120826 175339
rect 121870 175130 121930 175339
rect 123158 175130 123218 177651
rect 124446 175130 124506 177651
rect 125731 177036 125797 177037
rect 125731 176972 125732 177036
rect 125796 176972 125797 177036
rect 125731 176971 125797 176972
rect 125734 175130 125794 176971
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 131514 176600 132134 204618
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 137142 233069 137202 353907
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 137139 233068 137205 233069
rect 137139 233004 137140 233068
rect 137204 233004 137205 233068
rect 137139 233003 137205 233004
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 130699 175404 130765 175405
rect 130699 175340 130700 175404
rect 130764 175340 130765 175404
rect 130699 175339 130765 175340
rect 130702 175130 130762 175339
rect 132358 175130 132418 177651
rect 134379 177036 134445 177037
rect 134379 176972 134380 177036
rect 134444 176972 134445 177036
rect 134379 176971 134445 176972
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 176699
rect 134382 175130 134442 176971
rect 135234 176600 135854 208338
rect 138954 212614 139574 248058
rect 140822 242861 140882 380155
rect 141926 338330 141986 449923
rect 143582 389061 143642 499563
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 146523 462364 146589 462365
rect 146523 462300 146524 462364
rect 146588 462300 146589 462364
rect 146523 462299 146589 462300
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 143579 389060 143645 389061
rect 143579 388996 143580 389060
rect 143644 388996 143645 389060
rect 143579 388995 143645 388996
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 141926 338270 142354 338330
rect 142294 338061 142354 338270
rect 142291 338060 142357 338061
rect 142291 337996 142292 338060
rect 142356 337996 142357 338060
rect 142291 337995 142357 337996
rect 145794 327454 146414 362898
rect 146526 360365 146586 462299
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 146523 360364 146589 360365
rect 146523 360300 146524 360364
rect 146588 360300 146589 360364
rect 146523 360299 146589 360300
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 140819 242860 140885 242861
rect 140819 242796 140820 242860
rect 140884 242796 140885 242860
rect 140819 242795 140885 242796
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 160691 401708 160757 401709
rect 160691 401644 160692 401708
rect 160756 401644 160757 401708
rect 160691 401643 160757 401644
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 160694 215933 160754 401643
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 160691 215932 160757 215933
rect 160691 215868 160692 215932
rect 160756 215868 160757 215932
rect 160691 215867 160757 215868
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 168971 403068 169037 403069
rect 168971 403004 168972 403068
rect 169036 403004 169037 403068
rect 168971 403003 169037 403004
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 183700 166277 183701
rect 166211 183636 166212 183700
rect 166276 183636 166277 183700
rect 166211 183635 166277 183636
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 156093 166274 183635
rect 166395 180844 166461 180845
rect 166395 180780 166396 180844
rect 166460 180780 166461 180844
rect 166395 180779 166461 180780
rect 166398 158813 166458 180779
rect 167514 169174 168134 204618
rect 168974 181525 169034 403003
rect 170259 389876 170325 389877
rect 170259 389812 170260 389876
rect 170324 389812 170325 389876
rect 170259 389811 170325 389812
rect 168971 181524 169037 181525
rect 168971 181460 168972 181524
rect 169036 181460 169037 181524
rect 168971 181459 169037 181460
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166395 158812 166461 158813
rect 166395 158748 166396 158812
rect 166460 158748 166461 158812
rect 166395 158747 166461 158748
rect 166211 156092 166277 156093
rect 166211 156028 166212 156092
rect 166276 156028 166277 156092
rect 166211 156027 166277 156028
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 167514 133174 168134 168618
rect 168971 144940 169037 144941
rect 168971 144876 168972 144940
rect 169036 144876 169037 144940
rect 168971 144875 169037 144876
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 166395 132836 166461 132837
rect 166395 132772 166396 132836
rect 166460 132772 166461 132836
rect 166395 132771 166461 132772
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 166211 127124 166277 127125
rect 166211 127060 166212 127124
rect 166276 127060 166277 127124
rect 166211 127059 166277 127060
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66115 59940 66181 59941
rect 66115 59876 66116 59940
rect 66180 59876 66181 59940
rect 66115 59875 66181 59876
rect 64459 42260 64525 42261
rect 64459 42196 64460 42260
rect 64524 42196 64525 42260
rect 64459 42195 64525 42196
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 61883 19956 61949 19957
rect 61883 19892 61884 19956
rect 61948 19892 61949 19956
rect 61883 19891 61949 19892
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 85536 94757 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 85533 94756 85599 94757
rect 85533 94692 85534 94756
rect 85598 94692 85599 94756
rect 85533 94691 85599 94692
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 86726 92445 86786 94830
rect 88014 92445 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 86723 92444 86789 92445
rect 86723 92380 86724 92444
rect 86788 92380 86789 92444
rect 86723 92379 86789 92380
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88934 91765 88994 94830
rect 88931 91764 88997 91765
rect 88931 91700 88932 91764
rect 88996 91700 88997 91764
rect 88931 91699 88997 91700
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91221 96722 94830
rect 97214 91493 97274 94830
rect 98134 91493 98194 94830
rect 97211 91492 97277 91493
rect 97211 91428 97212 91492
rect 97276 91428 97277 91492
rect 97211 91427 97277 91428
rect 98131 91492 98197 91493
rect 98131 91428 98132 91492
rect 98196 91428 98197 91492
rect 98131 91427 98197 91428
rect 98502 91357 98562 94830
rect 99054 94830 99196 94890
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99054 91221 99114 94830
rect 99544 94754 99604 95200
rect 100632 94890 100692 95200
rect 100526 94830 100692 94890
rect 99544 94694 100034 94754
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 92445 100034 94694
rect 100526 93261 100586 94830
rect 100768 94754 100828 95200
rect 101856 94754 101916 95200
rect 100710 94694 100828 94754
rect 101814 94694 101916 94754
rect 101992 94754 102052 95200
rect 102944 94890 103004 95200
rect 102550 94830 103004 94890
rect 101992 94694 102058 94754
rect 100523 93260 100589 93261
rect 100523 93196 100524 93260
rect 100588 93196 100589 93260
rect 100523 93195 100589 93196
rect 99971 92444 100037 92445
rect 99971 92380 99972 92444
rect 100036 92380 100037 92444
rect 99971 92379 100037 92380
rect 100710 92309 100770 94694
rect 100707 92308 100773 92309
rect 100707 92244 100708 92308
rect 100772 92244 100773 92308
rect 100707 92243 100773 92244
rect 101814 92173 101874 94694
rect 101998 92445 102058 94694
rect 101995 92444 102061 92445
rect 101995 92380 101996 92444
rect 102060 92380 102061 92444
rect 101995 92379 102061 92380
rect 102550 92309 102610 94830
rect 103216 94754 103276 95200
rect 102734 94694 103276 94754
rect 104304 94754 104364 95200
rect 104440 94890 104500 95200
rect 104440 94830 104634 94890
rect 104304 94694 104450 94754
rect 102734 92445 102794 94694
rect 102731 92444 102797 92445
rect 102731 92380 102732 92444
rect 102796 92380 102797 92444
rect 102731 92379 102797 92380
rect 102547 92308 102613 92309
rect 102547 92244 102548 92308
rect 102612 92244 102613 92308
rect 102547 92243 102613 92244
rect 101811 92172 101877 92173
rect 101811 92108 101812 92172
rect 101876 92108 101877 92172
rect 101811 92107 101877 92108
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104390 92445 104450 94694
rect 104387 92444 104453 92445
rect 104387 92380 104388 92444
rect 104452 92380 104453 92444
rect 104387 92379 104453 92380
rect 104574 92309 104634 94830
rect 105392 94754 105452 95200
rect 105664 94754 105724 95200
rect 106480 94890 106540 95200
rect 106414 94830 106540 94890
rect 105392 94694 105554 94754
rect 105664 94694 105738 94754
rect 105494 92309 105554 94694
rect 105678 92445 105738 94694
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106414 92309 106474 94830
rect 106616 94754 106676 95200
rect 107704 94754 107764 95200
rect 108112 94754 108172 95200
rect 106598 94694 106676 94754
rect 107702 94694 107764 94754
rect 108070 94694 108172 94754
rect 109064 94754 109124 95200
rect 109472 94754 109532 95200
rect 110152 94754 110212 95200
rect 110696 94754 110756 95200
rect 111240 94754 111300 95200
rect 109064 94694 109234 94754
rect 109472 94694 109602 94754
rect 106598 92445 106658 94694
rect 107702 92445 107762 94694
rect 108070 92445 108130 94694
rect 109174 92445 109234 94694
rect 106595 92444 106661 92445
rect 106595 92380 106596 92444
rect 106660 92380 106661 92444
rect 106595 92379 106661 92380
rect 107699 92444 107765 92445
rect 107699 92380 107700 92444
rect 107764 92380 107765 92444
rect 107699 92379 107765 92380
rect 108067 92444 108133 92445
rect 108067 92380 108068 92444
rect 108132 92380 108133 92444
rect 108067 92379 108133 92380
rect 109171 92444 109237 92445
rect 109171 92380 109172 92444
rect 109236 92380 109237 92444
rect 109171 92379 109237 92380
rect 104571 92308 104637 92309
rect 104571 92244 104572 92308
rect 104636 92244 104637 92308
rect 104571 92243 104637 92244
rect 105491 92308 105557 92309
rect 105491 92244 105492 92308
rect 105556 92244 105557 92308
rect 105491 92243 105557 92244
rect 106411 92308 106477 92309
rect 106411 92244 106412 92308
rect 106476 92244 106477 92308
rect 106411 92243 106477 92244
rect 109542 91221 109602 94694
rect 110094 94694 110212 94754
rect 110646 94694 110756 94754
rect 111198 94694 111300 94754
rect 111920 94754 111980 95200
rect 112328 94757 112388 95200
rect 112325 94756 112391 94757
rect 111920 94694 111994 94754
rect 110094 93261 110154 94694
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 92445 110706 94694
rect 110643 92444 110709 92445
rect 110643 92380 110644 92444
rect 110708 92380 110709 92444
rect 110643 92379 110709 92380
rect 111198 91765 111258 94694
rect 111195 91764 111261 91765
rect 111195 91700 111196 91764
rect 111260 91700 111261 91764
rect 111195 91699 111261 91700
rect 111934 91221 111994 94694
rect 112325 94692 112326 94756
rect 112390 94692 112391 94756
rect 113144 94754 113204 95200
rect 113688 94754 113748 95200
rect 114368 94754 114428 95200
rect 114776 94754 114836 95200
rect 115456 94754 115516 95200
rect 115864 94754 115924 95200
rect 113144 94694 113282 94754
rect 113688 94694 114202 94754
rect 114368 94694 114570 94754
rect 114776 94694 114938 94754
rect 112325 94691 112391 94692
rect 113222 92445 113282 94694
rect 114142 93870 114202 94694
rect 114142 93810 114386 93870
rect 113219 92444 113285 92445
rect 113219 92380 113220 92444
rect 113284 92380 113285 92444
rect 113219 92379 113285 92380
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 93810
rect 114510 91765 114570 94694
rect 114507 91764 114573 91765
rect 114507 91700 114508 91764
rect 114572 91700 114573 91764
rect 114507 91699 114573 91700
rect 114878 91221 114938 94694
rect 115430 94694 115516 94754
rect 115798 94694 115924 94754
rect 116680 94754 116740 95200
rect 117088 94754 117148 95200
rect 116680 94694 116778 94754
rect 115430 91221 115490 94694
rect 115798 91357 115858 94694
rect 116718 92309 116778 94694
rect 117086 94694 117148 94754
rect 117904 94754 117964 95200
rect 118176 94754 118236 95200
rect 119400 94754 119460 95200
rect 117904 94694 118066 94754
rect 118176 94694 118250 94754
rect 116715 92308 116781 92309
rect 116715 92244 116716 92308
rect 116780 92244 116781 92308
rect 116715 92243 116781 92244
rect 117086 92173 117146 94694
rect 117083 92172 117149 92173
rect 117083 92108 117084 92172
rect 117148 92108 117149 92172
rect 117083 92107 117149 92108
rect 115795 91356 115861 91357
rect 115795 91292 115796 91356
rect 115860 91292 115861 91356
rect 115795 91291 115861 91292
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 115427 91220 115493 91221
rect 115427 91156 115428 91220
rect 115492 91156 115493 91220
rect 115427 91155 115493 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91629 118066 94694
rect 118003 91628 118069 91629
rect 118003 91564 118004 91628
rect 118068 91564 118069 91628
rect 118003 91563 118069 91564
rect 118190 91221 118250 94694
rect 119294 94694 119460 94754
rect 119536 94754 119596 95200
rect 120216 94754 120276 95200
rect 120624 94754 120684 95200
rect 121712 94754 121772 95200
rect 119536 94694 119722 94754
rect 119294 92445 119354 94694
rect 119662 92445 119722 94694
rect 120214 94694 120276 94754
rect 120582 94694 120684 94754
rect 121686 94694 121772 94754
rect 121984 94754 122044 95200
rect 122800 94757 122860 95200
rect 123208 94890 123268 95200
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124024 94830 124138 94890
rect 122797 94756 122863 94757
rect 121984 94694 122114 94754
rect 119291 92444 119357 92445
rect 119291 92380 119292 92444
rect 119356 92380 119357 92444
rect 119291 92379 119357 92380
rect 119659 92444 119725 92445
rect 119659 92380 119660 92444
rect 119724 92380 119725 92444
rect 119659 92379 119725 92380
rect 120214 91221 120274 94694
rect 120582 91629 120642 94694
rect 120579 91628 120645 91629
rect 120579 91564 120580 91628
rect 120644 91564 120645 91628
rect 120579 91563 120645 91564
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91221 121746 94694
rect 122054 91357 122114 94694
rect 122797 94692 122798 94756
rect 122862 94692 122863 94756
rect 122797 94691 122863 94692
rect 123158 93533 123218 94830
rect 123155 93532 123221 93533
rect 123155 93468 123156 93532
rect 123220 93468 123221 93532
rect 123155 93467 123221 93468
rect 122051 91356 122117 91357
rect 122051 91292 122052 91356
rect 122116 91292 122117 91356
rect 122051 91291 122117 91292
rect 124078 91221 124138 94830
rect 124432 94757 124492 95200
rect 125384 94890 125444 95200
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124429 94756 124495 94757
rect 124429 94692 124430 94756
rect 124494 94692 124495 94756
rect 124429 94691 124495 94692
rect 125366 91221 125426 94830
rect 125734 91221 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 126470 91221 126530 94830
rect 126654 91357 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 126651 91356 126717 91357
rect 126651 91292 126652 91356
rect 126716 91292 126717 91356
rect 126651 91291 126717 91292
rect 127574 91221 127634 94830
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 125731 91220 125797 91221
rect 125731 91156 125732 91220
rect 125796 91156 125797 91220
rect 125731 91155 125797 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 92445 129474 94830
rect 129411 92444 129477 92445
rect 129411 92380 129412 92444
rect 129476 92380 129477 92444
rect 129411 92379 129477 92380
rect 130702 91221 130762 94830
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 90949 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 92445 133154 94830
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 134382 91765 134442 94830
rect 134379 91764 134445 91765
rect 134379 91700 134380 91764
rect 134444 91700 134445 91764
rect 134379 91699 134445 91700
rect 132355 90948 132421 90949
rect 132355 90884 132356 90948
rect 132420 90884 132421 90948
rect 132355 90883 132421 90884
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151310 94830 151556 94890
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91221 151370 94830
rect 151491 94756 151557 94757
rect 151491 94692 151492 94756
rect 151556 94692 151557 94756
rect 151491 94691 151557 94692
rect 151494 92445 151554 94691
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 93669 151738 94150
rect 151675 93668 151741 93669
rect 151675 93604 151676 93668
rect 151740 93604 151741 93668
rect 151675 93603 151741 93604
rect 152046 92445 152106 94830
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151307 91220 151373 91221
rect 151307 91156 151308 91220
rect 151372 91156 151373 91220
rect 151307 91155 151373 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 80069 166274 127059
rect 166398 86869 166458 132771
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 168235 128484 168301 128485
rect 168235 128420 168236 128484
rect 168300 128420 168301 128484
rect 168235 128419 168301 128420
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 86868 166461 86869
rect 166395 86804 166396 86868
rect 166460 86804 166461 86868
rect 166395 86803 166461 86804
rect 166211 80068 166277 80069
rect 166211 80004 166212 80068
rect 166276 80004 166277 80068
rect 166211 80003 166277 80004
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 78573 168298 128419
rect 168974 90949 169034 144875
rect 170262 136101 170322 389811
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 173019 359412 173085 359413
rect 173019 359348 173020 359412
rect 173084 359348 173085 359412
rect 173019 359347 173085 359348
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 170443 136780 170509 136781
rect 170443 136716 170444 136780
rect 170508 136716 170509 136780
rect 170443 136715 170509 136716
rect 170259 136100 170325 136101
rect 170259 136036 170260 136100
rect 170324 136036 170325 136100
rect 170259 136035 170325 136036
rect 169155 135284 169221 135285
rect 169155 135220 169156 135284
rect 169220 135220 169221 135284
rect 169155 135219 169221 135220
rect 168971 90948 169037 90949
rect 168971 90884 168972 90948
rect 169036 90884 169037 90948
rect 168971 90883 169037 90884
rect 169158 84149 169218 135219
rect 170259 132700 170325 132701
rect 170259 132636 170260 132700
rect 170324 132636 170325 132700
rect 170259 132635 170325 132636
rect 169155 84148 169221 84149
rect 169155 84084 169156 84148
rect 169220 84084 169221 84148
rect 169155 84083 169221 84084
rect 168235 78572 168301 78573
rect 168235 78508 168236 78572
rect 168300 78508 168301 78572
rect 168235 78507 168301 78508
rect 170262 78437 170322 132635
rect 170446 82789 170506 136715
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 172099 128620 172165 128621
rect 172099 128556 172100 128620
rect 172164 128556 172165 128620
rect 172099 128555 172165 128556
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 82788 170509 82789
rect 170443 82724 170444 82788
rect 170508 82724 170509 82788
rect 170443 82723 170509 82724
rect 170259 78436 170325 78437
rect 170259 78372 170260 78436
rect 170324 78372 170325 78436
rect 170259 78371 170325 78372
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 172102 81429 172162 128555
rect 173022 83469 173082 359347
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 188291 374644 188357 374645
rect 188291 374580 188292 374644
rect 188356 374580 188357 374644
rect 188291 374579 188357 374580
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 184059 363628 184125 363629
rect 184059 363564 184060 363628
rect 184124 363564 184125 363628
rect 184059 363563 184125 363564
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 178539 320788 178605 320789
rect 178539 320724 178540 320788
rect 178604 320724 178605 320788
rect 178539 320723 178605 320724
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 178542 221509 178602 320723
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 178539 221508 178605 221509
rect 178539 221444 178540 221508
rect 178604 221444 178605 221508
rect 178539 221443 178605 221444
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173939 101420 174005 101421
rect 173939 101356 173940 101420
rect 174004 101356 174005 101420
rect 173939 101355 174005 101356
rect 173019 83468 173085 83469
rect 173019 83404 173020 83468
rect 173084 83404 173085 83468
rect 173019 83403 173085 83404
rect 172099 81428 172165 81429
rect 172099 81364 172100 81428
rect 172164 81364 172165 81428
rect 172099 81363 172165 81364
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 173942 3365 174002 101355
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 173939 3364 174005 3365
rect 173939 3300 173940 3364
rect 174004 3300 174005 3364
rect 173939 3299 174005 3300
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 184062 40629 184122 363563
rect 185514 331174 186134 366618
rect 186819 348396 186885 348397
rect 186819 348332 186820 348396
rect 186884 348332 186885 348396
rect 186819 348331 186885 348332
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 186822 43485 186882 348331
rect 186819 43484 186885 43485
rect 186819 43420 186820 43484
rect 186884 43420 186885 43484
rect 186819 43419 186885 43420
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 184059 40628 184125 40629
rect 184059 40564 184060 40628
rect 184124 40564 184125 40628
rect 184059 40563 184125 40564
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 188294 6901 188354 374579
rect 189234 370894 189854 406338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 191235 387836 191301 387837
rect 191235 387772 191236 387836
rect 191300 387772 191301 387836
rect 191235 387771 191301 387772
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 191051 351116 191117 351117
rect 191051 351052 191052 351116
rect 191116 351052 191117 351116
rect 191051 351051 191117 351052
rect 189947 345676 190013 345677
rect 189947 345612 189948 345676
rect 190012 345612 190013 345676
rect 189947 345611 190013 345612
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189950 46205 190010 345611
rect 189947 46204 190013 46205
rect 189947 46140 189948 46204
rect 190012 46140 190013 46204
rect 189947 46139 190013 46140
rect 191054 28253 191114 351051
rect 191238 87549 191298 387771
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 362000 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 362000 204134 384618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 362000 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 362000 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 362000 218414 362898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 362000 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 362000 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 362000 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 362000 236414 380898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 362000 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 362000 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 362000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 362000 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 362000 258134 366618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 362000 261854 370338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 362000 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 362000 272414 380898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 362000 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 362000 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 362000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 362000 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 362000 294134 366618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 362000 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 362000 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 362000 308414 380898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 362000 312134 384618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 362000 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 362000 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 321507 375460 321573 375461
rect 321507 375396 321508 375460
rect 321572 375396 321573 375460
rect 321507 375395 321573 375396
rect 320219 363220 320285 363221
rect 320219 363156 320220 363220
rect 320284 363156 320285 363220
rect 320219 363155 320285 363156
rect 320035 361860 320101 361861
rect 320035 361796 320036 361860
rect 320100 361796 320101 361860
rect 320035 361795 320101 361796
rect 200619 361724 200685 361725
rect 200619 361660 200620 361724
rect 200684 361660 200685 361724
rect 200619 361659 200685 361660
rect 199331 360228 199397 360229
rect 199331 360164 199332 360228
rect 199396 360164 199397 360228
rect 199331 360163 199397 360164
rect 197859 358324 197925 358325
rect 197859 358260 197860 358324
rect 197924 358260 197925 358324
rect 197859 358259 197925 358260
rect 195099 356692 195165 356693
rect 195099 356628 195100 356692
rect 195164 356628 195165 356692
rect 195099 356627 195165 356628
rect 193811 342956 193877 342957
rect 193811 342892 193812 342956
rect 193876 342892 193877 342956
rect 193811 342891 193877 342892
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192339 251292 192405 251293
rect 192339 251228 192340 251292
rect 192404 251228 192405 251292
rect 192339 251227 192405 251228
rect 192342 228309 192402 251227
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192339 228308 192405 228309
rect 192339 228244 192340 228308
rect 192404 228244 192405 228308
rect 192339 228243 192405 228244
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 191235 87548 191301 87549
rect 191235 87484 191236 87548
rect 191300 87484 191301 87548
rect 191235 87483 191301 87484
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 193814 86189 193874 342891
rect 193811 86188 193877 86189
rect 193811 86124 193812 86188
rect 193876 86124 193877 86188
rect 193811 86123 193877 86124
rect 192954 50614 193574 86058
rect 195102 82109 195162 356627
rect 197862 333301 197922 358259
rect 199334 353973 199394 360163
rect 199331 353972 199397 353973
rect 199331 353908 199332 353972
rect 199396 353908 199397 353972
rect 199331 353907 199397 353908
rect 200622 346357 200682 361659
rect 320038 355333 320098 361795
rect 320035 355332 320101 355333
rect 320035 355268 320036 355332
rect 320100 355268 320101 355332
rect 320035 355267 320101 355268
rect 200619 346356 200685 346357
rect 200619 346292 200620 346356
rect 200684 346292 200685 346356
rect 200619 346291 200685 346292
rect 219568 345454 219888 345486
rect 219568 345218 219610 345454
rect 219846 345218 219888 345454
rect 219568 345134 219888 345218
rect 219568 344898 219610 345134
rect 219846 344898 219888 345134
rect 219568 344866 219888 344898
rect 250288 345454 250608 345486
rect 250288 345218 250330 345454
rect 250566 345218 250608 345454
rect 250288 345134 250608 345218
rect 250288 344898 250330 345134
rect 250566 344898 250608 345134
rect 250288 344866 250608 344898
rect 281008 345454 281328 345486
rect 281008 345218 281050 345454
rect 281286 345218 281328 345454
rect 281008 345134 281328 345218
rect 281008 344898 281050 345134
rect 281286 344898 281328 345134
rect 281008 344866 281328 344898
rect 311728 345454 312048 345486
rect 311728 345218 311770 345454
rect 312006 345218 312048 345454
rect 311728 345134 312048 345218
rect 311728 344898 311770 345134
rect 312006 344898 312048 345134
rect 311728 344866 312048 344898
rect 197859 333300 197925 333301
rect 197859 333236 197860 333300
rect 197924 333236 197925 333300
rect 197859 333235 197925 333236
rect 204208 327454 204528 327486
rect 204208 327218 204250 327454
rect 204486 327218 204528 327454
rect 204208 327134 204528 327218
rect 204208 326898 204250 327134
rect 204486 326898 204528 327134
rect 204208 326866 204528 326898
rect 234928 327454 235248 327486
rect 234928 327218 234970 327454
rect 235206 327218 235248 327454
rect 234928 327134 235248 327218
rect 234928 326898 234970 327134
rect 235206 326898 235248 327134
rect 234928 326866 235248 326898
rect 265648 327454 265968 327486
rect 265648 327218 265690 327454
rect 265926 327218 265968 327454
rect 265648 327134 265968 327218
rect 265648 326898 265690 327134
rect 265926 326898 265968 327134
rect 265648 326866 265968 326898
rect 296368 327454 296688 327486
rect 296368 327218 296410 327454
rect 296646 327218 296688 327454
rect 296368 327134 296688 327218
rect 296368 326898 296410 327134
rect 296646 326898 296688 327134
rect 296368 326866 296688 326898
rect 219568 309454 219888 309486
rect 219568 309218 219610 309454
rect 219846 309218 219888 309454
rect 219568 309134 219888 309218
rect 219568 308898 219610 309134
rect 219846 308898 219888 309134
rect 219568 308866 219888 308898
rect 250288 309454 250608 309486
rect 250288 309218 250330 309454
rect 250566 309218 250608 309454
rect 250288 309134 250608 309218
rect 250288 308898 250330 309134
rect 250566 308898 250608 309134
rect 250288 308866 250608 308898
rect 281008 309454 281328 309486
rect 281008 309218 281050 309454
rect 281286 309218 281328 309454
rect 281008 309134 281328 309218
rect 281008 308898 281050 309134
rect 281286 308898 281328 309134
rect 281008 308866 281328 308898
rect 311728 309454 312048 309486
rect 311728 309218 311770 309454
rect 312006 309218 312048 309454
rect 311728 309134 312048 309218
rect 311728 308898 311770 309134
rect 312006 308898 312048 309134
rect 311728 308866 312048 308898
rect 204208 291454 204528 291486
rect 204208 291218 204250 291454
rect 204486 291218 204528 291454
rect 204208 291134 204528 291218
rect 204208 290898 204250 291134
rect 204486 290898 204528 291134
rect 204208 290866 204528 290898
rect 234928 291454 235248 291486
rect 234928 291218 234970 291454
rect 235206 291218 235248 291454
rect 234928 291134 235248 291218
rect 234928 290898 234970 291134
rect 235206 290898 235248 291134
rect 234928 290866 235248 290898
rect 265648 291454 265968 291486
rect 265648 291218 265690 291454
rect 265926 291218 265968 291454
rect 265648 291134 265968 291218
rect 265648 290898 265690 291134
rect 265926 290898 265968 291134
rect 265648 290866 265968 290898
rect 296368 291454 296688 291486
rect 296368 291218 296410 291454
rect 296646 291218 296688 291454
rect 296368 291134 296688 291218
rect 296368 290898 296410 291134
rect 296646 290898 296688 291134
rect 296368 290866 296688 290898
rect 219568 273454 219888 273486
rect 219568 273218 219610 273454
rect 219846 273218 219888 273454
rect 219568 273134 219888 273218
rect 219568 272898 219610 273134
rect 219846 272898 219888 273134
rect 219568 272866 219888 272898
rect 250288 273454 250608 273486
rect 250288 273218 250330 273454
rect 250566 273218 250608 273454
rect 250288 273134 250608 273218
rect 250288 272898 250330 273134
rect 250566 272898 250608 273134
rect 250288 272866 250608 272898
rect 281008 273454 281328 273486
rect 281008 273218 281050 273454
rect 281286 273218 281328 273454
rect 281008 273134 281328 273218
rect 281008 272898 281050 273134
rect 281286 272898 281328 273134
rect 281008 272866 281328 272898
rect 311728 273454 312048 273486
rect 311728 273218 311770 273454
rect 312006 273218 312048 273454
rect 311728 273134 312048 273218
rect 311728 272898 311770 273134
rect 312006 272898 312048 273134
rect 311728 272866 312048 272898
rect 204208 255454 204528 255486
rect 204208 255218 204250 255454
rect 204486 255218 204528 255454
rect 204208 255134 204528 255218
rect 204208 254898 204250 255134
rect 204486 254898 204528 255134
rect 204208 254866 204528 254898
rect 234928 255454 235248 255486
rect 234928 255218 234970 255454
rect 235206 255218 235248 255454
rect 234928 255134 235248 255218
rect 234928 254898 234970 255134
rect 235206 254898 235248 255134
rect 234928 254866 235248 254898
rect 265648 255454 265968 255486
rect 265648 255218 265690 255454
rect 265926 255218 265968 255454
rect 265648 255134 265968 255218
rect 265648 254898 265690 255134
rect 265926 254898 265968 255134
rect 265648 254866 265968 254898
rect 296368 255454 296688 255486
rect 296368 255218 296410 255454
rect 296646 255218 296688 255454
rect 296368 255134 296688 255218
rect 296368 254898 296410 255134
rect 296646 254898 296688 255134
rect 296368 254866 296688 254898
rect 197123 252516 197189 252517
rect 197123 252452 197124 252516
rect 197188 252452 197189 252516
rect 197123 252451 197189 252452
rect 196571 242180 196637 242181
rect 196571 242116 196572 242180
rect 196636 242116 196637 242180
rect 196571 242115 196637 242116
rect 196574 236061 196634 242115
rect 196571 236060 196637 236061
rect 196571 235996 196572 236060
rect 196636 235996 196637 236060
rect 196571 235995 196637 235996
rect 197126 180029 197186 252451
rect 320035 240412 320101 240413
rect 320035 240348 320036 240412
rect 320100 240348 320101 240412
rect 320035 240347 320101 240348
rect 200619 240276 200685 240277
rect 200619 240212 200620 240276
rect 200684 240212 200685 240276
rect 200619 240211 200685 240212
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 197123 180028 197189 180029
rect 197123 179964 197124 180028
rect 197188 179964 197189 180028
rect 197123 179963 197189 179964
rect 199794 165454 200414 200898
rect 200622 185605 200682 240211
rect 320038 238509 320098 240347
rect 320035 238508 320101 238509
rect 320035 238444 320036 238508
rect 320100 238444 320101 238508
rect 320035 238443 320101 238444
rect 203514 205174 204134 238000
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 200619 185604 200685 185605
rect 200619 185540 200620 185604
rect 200684 185540 200685 185604
rect 200619 185539 200685 185540
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 195099 82108 195165 82109
rect 195099 82044 195100 82108
rect 195164 82044 195165 82108
rect 195099 82043 195165 82044
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 191051 28252 191117 28253
rect 191051 28188 191052 28252
rect 191116 28188 191117 28252
rect 191051 28187 191117 28188
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 188291 6900 188357 6901
rect 188291 6836 188292 6900
rect 188356 6836 188357 6900
rect 188291 6835 188357 6836
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238000
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238000
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238000
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 226894 225854 238000
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 230614 229574 238000
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 239514 205174 240134 238000
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 178000 240134 204618
rect 243234 208894 243854 238000
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 178000 243854 208338
rect 246954 212614 247574 238000
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 178000 247574 212058
rect 253794 219454 254414 238000
rect 255267 231164 255333 231165
rect 255267 231100 255268 231164
rect 255332 231100 255333 231164
rect 255267 231099 255333 231100
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 249195 186964 249261 186965
rect 249195 186900 249196 186964
rect 249260 186900 249261 186964
rect 249195 186899 249261 186900
rect 214419 176900 214485 176901
rect 214419 176836 214420 176900
rect 214484 176836 214485 176900
rect 214419 176835 214485 176836
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 214422 164797 214482 176835
rect 249198 174317 249258 186899
rect 253794 183454 254414 218898
rect 254531 198116 254597 198117
rect 254531 198052 254532 198116
rect 254596 198052 254597 198116
rect 254531 198051 254597 198052
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 181388 252573 181389
rect 252507 181324 252508 181388
rect 252572 181324 252573 181388
rect 252507 181323 252573 181324
rect 249379 178668 249445 178669
rect 249379 178604 249380 178668
rect 249444 178604 249445 178668
rect 249379 178603 249445 178604
rect 249382 174725 249442 178603
rect 249379 174724 249445 174725
rect 249379 174660 249380 174724
rect 249444 174660 249445 174724
rect 249379 174659 249445 174660
rect 249195 174316 249261 174317
rect 249195 174252 249196 174316
rect 249260 174252 249261 174316
rect 249195 174251 249261 174252
rect 227874 165454 228194 165486
rect 227874 165218 227916 165454
rect 228152 165218 228194 165454
rect 227874 165134 228194 165218
rect 227874 164898 227916 165134
rect 228152 164898 228194 165134
rect 227874 164866 228194 164898
rect 237805 165454 238125 165486
rect 237805 165218 237847 165454
rect 238083 165218 238125 165454
rect 237805 165134 238125 165218
rect 237805 164898 237847 165134
rect 238083 164898 238125 165134
rect 237805 164866 238125 164898
rect 214419 164796 214485 164797
rect 214419 164732 214420 164796
rect 214484 164732 214485 164796
rect 214419 164731 214485 164732
rect 251771 149700 251837 149701
rect 251771 149636 251772 149700
rect 251836 149636 251837 149700
rect 251771 149635 251837 149636
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 227874 129454 228194 129486
rect 227874 129218 227916 129454
rect 228152 129218 228194 129454
rect 227874 129134 228194 129218
rect 227874 128898 227916 129134
rect 228152 128898 228194 129134
rect 227874 128866 228194 128898
rect 237805 129454 238125 129486
rect 237805 129218 237847 129454
rect 238083 129218 238125 129454
rect 237805 129134 238125 129218
rect 237805 128898 237847 129134
rect 238083 128898 238125 129134
rect 237805 128866 238125 128898
rect 251774 123045 251834 149635
rect 252510 144669 252570 181323
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 252507 144668 252573 144669
rect 252507 144604 252508 144668
rect 252572 144604 252573 144668
rect 252507 144603 252573 144604
rect 253611 138412 253677 138413
rect 253611 138348 253612 138412
rect 253676 138348 253677 138412
rect 253611 138347 253677 138348
rect 251955 123316 252021 123317
rect 251955 123252 251956 123316
rect 252020 123252 252021 123316
rect 251955 123251 252021 123252
rect 251771 123044 251837 123045
rect 251771 122980 251772 123044
rect 251836 122980 251837 123044
rect 251771 122979 251837 122980
rect 249563 114884 249629 114885
rect 249563 114820 249564 114884
rect 249628 114820 249629 114884
rect 249563 114819 249629 114820
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 214603 105228 214669 105229
rect 214603 105164 214604 105228
rect 214668 105164 214669 105228
rect 214603 105163 214669 105164
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 103596 214485 103597
rect 214419 103532 214420 103596
rect 214484 103532 214485 103596
rect 214419 103531 214485 103532
rect 214422 91085 214482 103531
rect 214606 93805 214666 105163
rect 249566 103530 249626 114819
rect 249198 103470 249626 103530
rect 214603 93804 214669 93805
rect 214603 93740 214604 93804
rect 214668 93740 214669 93804
rect 214603 93739 214669 93740
rect 214419 91084 214485 91085
rect 214419 91020 214420 91084
rect 214484 91020 214485 91084
rect 214419 91019 214485 91020
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 94000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 94000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 94000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 249198 11661 249258 103470
rect 249379 98428 249445 98429
rect 249379 98364 249380 98428
rect 249444 98364 249445 98428
rect 249379 98363 249445 98364
rect 249195 11660 249261 11661
rect 249195 11596 249196 11660
rect 249260 11596 249261 11660
rect 249195 11595 249261 11596
rect 249382 10301 249442 98363
rect 251958 97069 252018 123251
rect 253614 122850 253674 138347
rect 253062 122790 253674 122850
rect 251955 97068 252021 97069
rect 251955 97004 251956 97068
rect 252020 97004 252021 97068
rect 251955 97003 252021 97004
rect 253062 37909 253122 122790
rect 253794 111454 254414 146898
rect 254534 146573 254594 198051
rect 255270 156365 255330 231099
rect 257514 223174 258134 238000
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 261234 226894 261854 238000
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 258579 204916 258645 204917
rect 258579 204852 258580 204916
rect 258644 204852 258645 204916
rect 258579 204851 258645 204852
rect 258395 191180 258461 191181
rect 258395 191116 258396 191180
rect 258460 191116 258461 191180
rect 258395 191115 258461 191116
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 256739 184380 256805 184381
rect 256739 184316 256740 184380
rect 256804 184316 256805 184380
rect 256739 184315 256805 184316
rect 255451 180300 255517 180301
rect 255451 180236 255452 180300
rect 255516 180236 255517 180300
rect 255451 180235 255517 180236
rect 255267 156364 255333 156365
rect 255267 156300 255268 156364
rect 255332 156300 255333 156364
rect 255267 156299 255333 156300
rect 254531 146572 254597 146573
rect 254531 146508 254532 146572
rect 254596 146508 254597 146572
rect 254531 146507 254597 146508
rect 255454 141133 255514 180235
rect 256742 170917 256802 184315
rect 256739 170916 256805 170917
rect 256739 170852 256740 170916
rect 256804 170852 256805 170916
rect 256739 170851 256805 170852
rect 257514 151174 258134 186618
rect 258398 180810 258458 191115
rect 258214 180750 258458 180810
rect 258214 171150 258274 180750
rect 258214 171090 258458 171150
rect 258398 160989 258458 171090
rect 258395 160988 258461 160989
rect 258395 160924 258396 160988
rect 258460 160924 258461 160988
rect 258395 160923 258461 160924
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 255451 141132 255517 141133
rect 255451 141068 255452 141132
rect 255516 141068 255517 141132
rect 255451 141067 255517 141068
rect 257291 134196 257357 134197
rect 257291 134132 257292 134196
rect 257356 134132 257357 134196
rect 257291 134131 257357 134132
rect 255819 128756 255885 128757
rect 255819 128692 255820 128756
rect 255884 128692 255885 128756
rect 255819 128691 255885 128692
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 37908 253125 37909
rect 253059 37844 253060 37908
rect 253124 37844 253125 37908
rect 253059 37843 253125 37844
rect 249379 10300 249445 10301
rect 249379 10236 249380 10300
rect 249444 10236 249445 10300
rect 249379 10235 249445 10236
rect 253794 3454 254414 38898
rect 255822 14517 255882 128691
rect 257294 51781 257354 134131
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257291 51780 257357 51781
rect 257291 51716 257292 51780
rect 257356 51716 257357 51780
rect 257291 51715 257357 51716
rect 257514 43174 258134 78618
rect 258582 67557 258642 204851
rect 259499 200700 259565 200701
rect 259499 200636 259500 200700
rect 259564 200636 259565 200700
rect 259499 200635 259565 200636
rect 259502 145077 259562 200635
rect 259683 191044 259749 191045
rect 259683 190980 259684 191044
rect 259748 190980 259749 191044
rect 259683 190979 259749 190980
rect 259499 145076 259565 145077
rect 259499 145012 259500 145076
rect 259564 145012 259565 145076
rect 259499 145011 259565 145012
rect 259686 140997 259746 190979
rect 261234 190894 261854 226338
rect 264954 230614 265574 238000
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263547 206276 263613 206277
rect 263547 206212 263548 206276
rect 263612 206212 263613 206276
rect 263547 206211 263613 206212
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 262259 189684 262325 189685
rect 262259 189620 262260 189684
rect 262324 189620 262325 189684
rect 262259 189619 262325 189620
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 259683 140996 259749 140997
rect 259683 140932 259684 140996
rect 259748 140932 259749 140996
rect 259683 140931 259749 140932
rect 261234 118894 261854 154338
rect 262262 138277 262322 189619
rect 262443 180164 262509 180165
rect 262443 180100 262444 180164
rect 262508 180100 262509 180164
rect 262443 180099 262509 180100
rect 262446 154597 262506 180099
rect 262443 154596 262509 154597
rect 262443 154532 262444 154596
rect 262508 154532 262509 154596
rect 262443 154531 262509 154532
rect 263550 140861 263610 206211
rect 264954 194614 265574 230058
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 268331 215932 268397 215933
rect 268331 215868 268332 215932
rect 268396 215868 268397 215932
rect 268331 215867 268397 215868
rect 266307 195396 266373 195397
rect 266307 195332 266308 195396
rect 266372 195332 266373 195396
rect 266307 195331 266373 195332
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263731 187100 263797 187101
rect 263731 187036 263732 187100
rect 263796 187036 263797 187100
rect 263731 187035 263797 187036
rect 263734 163165 263794 187035
rect 263731 163164 263797 163165
rect 263731 163100 263732 163164
rect 263796 163100 263797 163164
rect 263731 163099 263797 163100
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 263547 140860 263613 140861
rect 263547 140796 263548 140860
rect 263612 140796 263613 140860
rect 263547 140795 263613 140796
rect 262259 138276 262325 138277
rect 262259 138212 262260 138276
rect 262324 138212 262325 138276
rect 262259 138211 262325 138212
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 258579 67556 258645 67557
rect 258579 67492 258580 67556
rect 258644 67492 258645 67556
rect 258579 67491 258645 67492
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 255819 14516 255885 14517
rect 255819 14452 255820 14516
rect 255884 14452 255885 14516
rect 255819 14451 255885 14452
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 122614 265574 158058
rect 266310 142221 266370 195331
rect 266307 142220 266373 142221
rect 266307 142156 266308 142220
rect 266372 142156 266373 142220
rect 266307 142155 266373 142156
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 268334 35189 268394 215867
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 269067 178804 269133 178805
rect 269067 178740 269068 178804
rect 269132 178740 269133 178804
rect 269067 178739 269133 178740
rect 269070 148069 269130 178739
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 269067 148068 269133 148069
rect 269067 148004 269068 148068
rect 269132 148004 269133 148068
rect 269067 148003 269133 148004
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 268331 35188 268397 35189
rect 268331 35124 268332 35188
rect 268396 35124 268397 35188
rect 268331 35123 268397 35124
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 205174 276134 238000
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 208894 279854 238000
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 212614 283574 238000
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 219454 290414 238000
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 223174 294134 238000
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 226894 297854 238000
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 300954 230614 301574 238000
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 307794 237454 308414 238000
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 311514 205174 312134 238000
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 178000 312134 204618
rect 315234 208894 315854 238000
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 178000 315854 208338
rect 318954 212614 319574 238000
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 178000 319574 212058
rect 320222 175813 320282 363155
rect 321510 352205 321570 375395
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 321507 352204 321573 352205
rect 321507 352140 321508 352204
rect 321572 352140 321573 352204
rect 321507 352139 321573 352140
rect 325794 327454 326414 362898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 332915 369884 332981 369885
rect 332915 369820 332916 369884
rect 332980 369820 332981 369884
rect 332915 369819 332981 369820
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 327027 354244 327093 354245
rect 327027 354180 327028 354244
rect 327092 354180 327093 354244
rect 327027 354179 327093 354180
rect 326659 331124 326725 331125
rect 326659 331060 326660 331124
rect 326724 331060 326725 331124
rect 326659 331059 326725 331060
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 321507 318884 321573 318885
rect 321507 318820 321508 318884
rect 321572 318820 321573 318884
rect 321507 318819 321573 318820
rect 321510 236605 321570 318819
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 321507 236604 321573 236605
rect 321507 236540 321508 236604
rect 321572 236540 321573 236604
rect 321507 236539 321573 236540
rect 321507 224500 321573 224501
rect 321507 224436 321508 224500
rect 321572 224436 321573 224500
rect 321507 224435 321573 224436
rect 321323 181524 321389 181525
rect 321323 181460 321324 181524
rect 321388 181460 321389 181524
rect 321323 181459 321389 181460
rect 320219 175812 320285 175813
rect 320219 175748 320220 175812
rect 320284 175748 320285 175812
rect 320219 175747 320285 175748
rect 321326 170645 321386 181459
rect 321323 170644 321389 170645
rect 321323 170580 321324 170644
rect 321388 170580 321389 170644
rect 321323 170579 321389 170580
rect 314208 165454 314528 165486
rect 314208 165218 314250 165454
rect 314486 165218 314528 165454
rect 314208 165134 314528 165218
rect 314208 164898 314250 165134
rect 314486 164898 314528 165134
rect 314208 164866 314528 164898
rect 317472 165454 317792 165486
rect 317472 165218 317514 165454
rect 317750 165218 317792 165454
rect 317472 165134 317792 165218
rect 317472 164898 317514 165134
rect 317750 164898 317792 165134
rect 317472 164866 317792 164898
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 306971 141268 307037 141269
rect 306971 141204 306972 141268
rect 307036 141204 307037 141268
rect 306971 141203 307037 141204
rect 305499 129844 305565 129845
rect 305499 129780 305500 129844
rect 305564 129780 305565 129844
rect 305499 129779 305565 129780
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 302739 114340 302805 114341
rect 302739 114276 302740 114340
rect 302804 114276 302805 114340
rect 302739 114275 302805 114276
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300715 76532 300781 76533
rect 300715 76468 300716 76532
rect 300780 76468 300781 76532
rect 300715 76467 300781 76468
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 300718 39541 300778 76467
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300715 39540 300781 39541
rect 300715 39476 300716 39540
rect 300780 39476 300781 39540
rect 300715 39475 300781 39476
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 302742 4861 302802 114275
rect 304211 101148 304277 101149
rect 304211 101084 304212 101148
rect 304276 101084 304277 101148
rect 304211 101083 304277 101084
rect 304214 42125 304274 101083
rect 304211 42124 304277 42125
rect 304211 42060 304212 42124
rect 304276 42060 304277 42124
rect 304211 42059 304277 42060
rect 305502 17237 305562 129779
rect 306974 119373 307034 141203
rect 321510 131069 321570 224435
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 321691 176220 321757 176221
rect 321691 176156 321692 176220
rect 321756 176156 321757 176220
rect 321691 176155 321757 176156
rect 321694 155277 321754 176155
rect 321691 155276 321757 155277
rect 321691 155212 321692 155276
rect 321756 155212 321757 155276
rect 321691 155211 321757 155212
rect 325794 147454 326414 182898
rect 326662 149701 326722 331059
rect 326659 149700 326725 149701
rect 326659 149636 326660 149700
rect 326724 149636 326725 149700
rect 326659 149635 326725 149636
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 321507 131068 321573 131069
rect 321507 131004 321508 131068
rect 321572 131004 321573 131068
rect 321507 131003 321573 131004
rect 314208 129454 314528 129486
rect 314208 129218 314250 129454
rect 314486 129218 314528 129454
rect 314208 129134 314528 129218
rect 314208 128898 314250 129134
rect 314486 128898 314528 129134
rect 314208 128866 314528 128898
rect 317472 129454 317792 129486
rect 317472 129218 317514 129454
rect 317750 129218 317792 129454
rect 317472 129134 317792 129218
rect 317472 128898 317514 129134
rect 317750 128898 317792 129134
rect 317472 128866 317792 128898
rect 307155 127668 307221 127669
rect 307155 127604 307156 127668
rect 307220 127604 307221 127668
rect 307155 127603 307221 127604
rect 306971 119372 307037 119373
rect 306971 119308 306972 119372
rect 307036 119308 307037 119372
rect 306971 119307 307037 119308
rect 306971 97068 307037 97069
rect 306971 97004 306972 97068
rect 307036 97004 307037 97068
rect 306971 97003 307037 97004
rect 306974 18597 307034 97003
rect 307158 84829 307218 127603
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 327030 139365 327090 354179
rect 329514 331174 330134 366618
rect 330339 364444 330405 364445
rect 330339 364380 330340 364444
rect 330404 364380 330405 364444
rect 330339 364379 330405 364380
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 328499 232524 328565 232525
rect 328499 232460 328500 232524
rect 328564 232460 328565 232524
rect 328499 232459 328565 232460
rect 327027 139364 327093 139365
rect 327027 139300 327028 139364
rect 327092 139300 327093 139364
rect 327027 139299 327093 139300
rect 328502 125629 328562 232459
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 328499 125628 328565 125629
rect 328499 125564 328500 125628
rect 328564 125564 328565 125628
rect 328499 125563 328565 125564
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 321507 109580 321573 109581
rect 321507 109516 321508 109580
rect 321572 109516 321573 109580
rect 321507 109515 321573 109516
rect 321510 95165 321570 109515
rect 324267 98564 324333 98565
rect 324267 98500 324268 98564
rect 324332 98500 324333 98564
rect 324267 98499 324333 98500
rect 321507 95164 321573 95165
rect 321507 95100 321508 95164
rect 321572 95100 321573 95164
rect 321507 95099 321573 95100
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 84828 307221 84829
rect 307155 84764 307156 84828
rect 307220 84764 307221 84828
rect 307155 84763 307221 84764
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 18596 307037 18597
rect 306971 18532 306972 18596
rect 307036 18532 307037 18596
rect 306971 18531 307037 18532
rect 305499 17236 305565 17237
rect 305499 17172 305500 17236
rect 305564 17172 305565 17236
rect 305499 17171 305565 17172
rect 302739 4860 302805 4861
rect 302739 4796 302740 4860
rect 302804 4796 302805 4860
rect 302739 4795 302805 4796
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 94000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 94000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 94000
rect 324270 93669 324330 98499
rect 324267 93668 324333 93669
rect 324267 93604 324268 93668
rect 324332 93604 324333 93668
rect 324267 93603 324333 93604
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 115174 330134 150618
rect 330342 139501 330402 364379
rect 331259 358052 331325 358053
rect 331259 357988 331260 358052
rect 331324 357988 331325 358052
rect 331259 357987 331325 357988
rect 330339 139500 330405 139501
rect 330339 139436 330340 139500
rect 330404 139436 330405 139500
rect 330339 139435 330405 139436
rect 331262 131205 331322 357987
rect 331443 178668 331509 178669
rect 331443 178604 331444 178668
rect 331508 178604 331509 178668
rect 331443 178603 331509 178604
rect 331446 144125 331506 178603
rect 332918 175269 332978 369819
rect 333234 334894 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 338251 407148 338317 407149
rect 338251 407084 338252 407148
rect 338316 407084 338317 407148
rect 338251 407083 338317 407084
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 334571 360364 334637 360365
rect 334571 360300 334572 360364
rect 334636 360300 334637 360364
rect 334571 360299 334637 360300
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 332915 175268 332981 175269
rect 332915 175204 332916 175268
rect 332980 175204 332981 175268
rect 332915 175203 332981 175204
rect 332915 172548 332981 172549
rect 332915 172484 332916 172548
rect 332980 172484 332981 172548
rect 332915 172483 332981 172484
rect 331443 144124 331509 144125
rect 331443 144060 331444 144124
rect 331508 144060 331509 144124
rect 331443 144059 331509 144060
rect 331259 131204 331325 131205
rect 331259 131140 331260 131204
rect 331324 131140 331325 131204
rect 331259 131139 331325 131140
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 332918 80749 332978 172483
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 334574 117333 334634 360299
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336043 197980 336109 197981
rect 336043 197916 336044 197980
rect 336108 197916 336109 197980
rect 336043 197915 336109 197916
rect 334755 171188 334821 171189
rect 334755 171124 334756 171188
rect 334820 171124 334821 171188
rect 334755 171123 334821 171124
rect 334571 117332 334637 117333
rect 334571 117268 334572 117332
rect 334636 117268 334637 117332
rect 334571 117267 334637 117268
rect 334758 87549 334818 171123
rect 335859 169828 335925 169829
rect 335859 169764 335860 169828
rect 335924 169764 335925 169828
rect 335859 169763 335925 169764
rect 334755 87548 334821 87549
rect 334755 87484 334756 87548
rect 334820 87484 334821 87548
rect 334755 87483 334821 87484
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 332915 80748 332981 80749
rect 332915 80684 332916 80748
rect 332980 80684 332981 80748
rect 332915 80683 332981 80684
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 82338
rect 335862 79389 335922 169763
rect 336046 144805 336106 197915
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336043 144804 336109 144805
rect 336043 144740 336044 144804
rect 336108 144740 336109 144804
rect 336043 144739 336109 144740
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 335859 79388 335925 79389
rect 335859 79324 335860 79388
rect 335924 79324 335925 79388
rect 335859 79323 335925 79324
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 86058
rect 338254 78573 338314 407083
rect 340091 404428 340157 404429
rect 340091 404364 340092 404428
rect 340156 404364 340157 404428
rect 340091 404363 340157 404364
rect 338619 158812 338685 158813
rect 338619 158748 338620 158812
rect 338684 158748 338685 158812
rect 338619 158747 338685 158748
rect 338251 78572 338317 78573
rect 338251 78508 338252 78572
rect 338316 78508 338317 78572
rect 338251 78507 338317 78508
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 338622 45525 338682 158747
rect 340094 148341 340154 404363
rect 340827 385660 340893 385661
rect 340827 385596 340828 385660
rect 340892 385596 340893 385660
rect 340827 385595 340893 385596
rect 340275 162892 340341 162893
rect 340275 162828 340276 162892
rect 340340 162828 340341 162892
rect 340275 162827 340341 162828
rect 340091 148340 340157 148341
rect 340091 148276 340092 148340
rect 340156 148276 340157 148340
rect 340091 148275 340157 148276
rect 340278 83469 340338 162827
rect 340275 83468 340341 83469
rect 340275 83404 340276 83468
rect 340340 83404 340341 83468
rect 340275 83403 340341 83404
rect 340830 46205 340890 385595
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 345611 361996 345677 361997
rect 345611 361932 345612 361996
rect 345676 361932 345677 361996
rect 345611 361931 345677 361932
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342851 178124 342917 178125
rect 342851 178060 342852 178124
rect 342916 178060 342917 178124
rect 342851 178059 342917 178060
rect 342854 84965 342914 178059
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 345614 113253 345674 361931
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 345611 113252 345677 113253
rect 345611 113188 345612 113252
rect 345676 113188 345677 113252
rect 345611 113187 345677 113188
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 342851 84964 342917 84965
rect 342851 84900 342852 84964
rect 342916 84900 342917 84964
rect 342851 84899 342917 84900
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 340827 46204 340893 46205
rect 340827 46140 340828 46204
rect 340892 46140 340893 46204
rect 340827 46139 340893 46140
rect 338619 45524 338685 45525
rect 338619 45460 338620 45524
rect 338684 45460 338685 45524
rect 338619 45459 338685 45460
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 340830 11797 340890 46139
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 340827 11796 340893 11797
rect 340827 11732 340828 11796
rect 340892 11732 340893 11796
rect 340827 11731 340893 11732
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 181600 420134 204618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 181600 423854 208338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 181600 427574 212058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 181600 434414 182898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 181600 438134 186618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 181600 441854 190338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 181600 445574 194058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 181600 452414 200898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 181600 456134 204618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 181600 459854 208338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 181600 463574 212058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 181600 470414 182898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 181600 474134 186618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 181600 477854 190338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 181600 481574 194058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 181600 488414 200898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 181600 492134 204618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 181600 495854 208338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 494099 177308 494165 177309
rect 494099 177244 494100 177308
rect 494164 177244 494165 177308
rect 494099 177243 494165 177244
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 439568 165454 439888 165486
rect 439568 165218 439610 165454
rect 439846 165218 439888 165454
rect 439568 165134 439888 165218
rect 439568 164898 439610 165134
rect 439846 164898 439888 165134
rect 439568 164866 439888 164898
rect 470288 165454 470608 165486
rect 470288 165218 470330 165454
rect 470566 165218 470608 165454
rect 470288 165134 470608 165218
rect 470288 164898 470330 165134
rect 470566 164898 470608 165134
rect 470288 164866 470608 164898
rect 424208 147454 424528 147486
rect 424208 147218 424250 147454
rect 424486 147218 424528 147454
rect 424208 147134 424528 147218
rect 424208 146898 424250 147134
rect 424486 146898 424528 147134
rect 424208 146866 424528 146898
rect 454928 147454 455248 147486
rect 454928 147218 454970 147454
rect 455206 147218 455248 147454
rect 454928 147134 455248 147218
rect 454928 146898 454970 147134
rect 455206 146898 455248 147134
rect 454928 146866 455248 146898
rect 485648 147454 485968 147486
rect 485648 147218 485690 147454
rect 485926 147218 485968 147454
rect 485648 147134 485968 147218
rect 485648 146898 485690 147134
rect 485926 146898 485968 147134
rect 485648 146866 485968 146898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 439568 129454 439888 129486
rect 439568 129218 439610 129454
rect 439846 129218 439888 129454
rect 439568 129134 439888 129218
rect 439568 128898 439610 129134
rect 439846 128898 439888 129134
rect 439568 128866 439888 128898
rect 470288 129454 470608 129486
rect 470288 129218 470330 129454
rect 470566 129218 470608 129454
rect 470288 129134 470608 129218
rect 470288 128898 470330 129134
rect 470566 128898 470608 129134
rect 470288 128866 470608 128898
rect 424208 111454 424528 111486
rect 424208 111218 424250 111454
rect 424486 111218 424528 111454
rect 424208 111134 424528 111218
rect 424208 110898 424250 111134
rect 424486 110898 424528 111134
rect 424208 110866 424528 110898
rect 454928 111454 455248 111486
rect 454928 111218 454970 111454
rect 455206 111218 455248 111454
rect 454928 111134 455248 111218
rect 454928 110898 454970 111134
rect 455206 110898 455248 111134
rect 454928 110866 455248 110898
rect 485648 111454 485968 111486
rect 485648 111218 485690 111454
rect 485926 111218 485968 111454
rect 485648 111134 485968 111218
rect 485648 110898 485690 111134
rect 485926 110898 485968 111134
rect 485648 110866 485968 110898
rect 493915 102236 493981 102237
rect 493915 102172 493916 102236
rect 493980 102172 493981 102236
rect 493915 102171 493981 102172
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 97174 420134 98000
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 98000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 68614 427574 98000
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 75454 434414 98000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 79174 438134 98000
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 82894 441854 98000
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 98000
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 93454 452414 98000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 97174 456134 98000
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 64894 459854 98000
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 68614 463574 98000
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 75454 470414 98000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 79174 474134 98000
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 82894 477854 98000
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 86614 481574 98000
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 93454 488414 98000
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 97174 492134 98000
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 493918 96525 493978 102171
rect 493915 96524 493981 96525
rect 493915 96460 493916 96524
rect 493980 96460 493981 96524
rect 493915 96459 493981 96460
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 494102 15197 494162 177243
rect 498954 176614 499574 212058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 502379 189684 502445 189685
rect 502379 189620 502380 189684
rect 502444 189620 502445 189684
rect 502379 189619 502445 189620
rect 499803 176764 499869 176765
rect 499803 176700 499804 176764
rect 499868 176700 499869 176764
rect 499803 176699 499869 176700
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 496859 174452 496925 174453
rect 496859 174388 496860 174452
rect 496924 174388 496925 174452
rect 496859 174387 496925 174388
rect 494467 171460 494533 171461
rect 494467 171396 494468 171460
rect 494532 171396 494533 171460
rect 494467 171395 494533 171396
rect 494470 98701 494530 171395
rect 494467 98700 494533 98701
rect 494467 98636 494468 98700
rect 494532 98636 494533 98700
rect 494467 98635 494533 98636
rect 495234 64894 495854 98000
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 494099 15196 494165 15197
rect 494099 15132 494100 15196
rect 494164 15132 494165 15196
rect 494099 15131 494165 15132
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28338
rect 496862 4045 496922 174387
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 496859 4044 496925 4045
rect 496859 3980 496860 4044
rect 496924 3980 496925 4044
rect 496859 3979 496925 3980
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 499806 8261 499866 176699
rect 502382 110533 502442 189619
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 502379 110532 502445 110533
rect 502379 110468 502380 110532
rect 502444 110468 502445 110532
rect 502379 110467 502445 110468
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 499803 8260 499869 8261
rect 499803 8196 499804 8260
rect 499868 8196 499869 8260
rect 499803 8195 499869 8196
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 76618 579218 76854 579454
rect 76618 578898 76854 579134
rect 87882 579218 88118 579454
rect 87882 578898 88118 579134
rect 99146 579218 99382 579454
rect 99146 578898 99382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 82250 561218 82486 561454
rect 82250 560898 82486 561134
rect 93514 561218 93750 561454
rect 93514 560898 93750 561134
rect 76618 543218 76854 543454
rect 76618 542898 76854 543134
rect 87882 543218 88118 543454
rect 87882 542898 88118 543134
rect 99146 543218 99382 543454
rect 99146 542898 99382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 75618 471218 75854 471454
rect 75618 470898 75854 471134
rect 84882 471218 85118 471454
rect 84882 470898 85118 471134
rect 94146 471218 94382 471454
rect 94146 470898 94382 471134
rect 80250 453218 80486 453454
rect 80250 452898 80486 453134
rect 89514 453218 89750 453454
rect 89514 452898 89750 453134
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 219610 345218 219846 345454
rect 219610 344898 219846 345134
rect 250330 345218 250566 345454
rect 250330 344898 250566 345134
rect 281050 345218 281286 345454
rect 281050 344898 281286 345134
rect 311770 345218 312006 345454
rect 311770 344898 312006 345134
rect 204250 327218 204486 327454
rect 204250 326898 204486 327134
rect 234970 327218 235206 327454
rect 234970 326898 235206 327134
rect 265690 327218 265926 327454
rect 265690 326898 265926 327134
rect 296410 327218 296646 327454
rect 296410 326898 296646 327134
rect 219610 309218 219846 309454
rect 219610 308898 219846 309134
rect 250330 309218 250566 309454
rect 250330 308898 250566 309134
rect 281050 309218 281286 309454
rect 281050 308898 281286 309134
rect 311770 309218 312006 309454
rect 311770 308898 312006 309134
rect 204250 291218 204486 291454
rect 204250 290898 204486 291134
rect 234970 291218 235206 291454
rect 234970 290898 235206 291134
rect 265690 291218 265926 291454
rect 265690 290898 265926 291134
rect 296410 291218 296646 291454
rect 296410 290898 296646 291134
rect 219610 273218 219846 273454
rect 219610 272898 219846 273134
rect 250330 273218 250566 273454
rect 250330 272898 250566 273134
rect 281050 273218 281286 273454
rect 281050 272898 281286 273134
rect 311770 273218 312006 273454
rect 311770 272898 312006 273134
rect 204250 255218 204486 255454
rect 204250 254898 204486 255134
rect 234970 255218 235206 255454
rect 234970 254898 235206 255134
rect 265690 255218 265926 255454
rect 265690 254898 265926 255134
rect 296410 255218 296646 255454
rect 296410 254898 296646 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 227916 165218 228152 165454
rect 227916 164898 228152 165134
rect 237847 165218 238083 165454
rect 237847 164898 238083 165134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 227916 129218 228152 129454
rect 227916 128898 228152 129134
rect 237847 129218 238083 129454
rect 237847 128898 238083 129134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 314250 165218 314486 165454
rect 314250 164898 314486 165134
rect 317514 165218 317750 165454
rect 317514 164898 317750 165134
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 314250 129218 314486 129454
rect 314250 128898 314486 129134
rect 317514 129218 317750 129454
rect 317514 128898 317750 129134
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 439610 165218 439846 165454
rect 439610 164898 439846 165134
rect 470330 165218 470566 165454
rect 470330 164898 470566 165134
rect 424250 147218 424486 147454
rect 424250 146898 424486 147134
rect 454970 147218 455206 147454
rect 454970 146898 455206 147134
rect 485690 147218 485926 147454
rect 485690 146898 485926 147134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 439610 129218 439846 129454
rect 439610 128898 439846 129134
rect 470330 129218 470566 129454
rect 470330 128898 470566 129134
rect 424250 111218 424486 111454
rect 424250 110898 424486 111134
rect 454970 111218 455206 111454
rect 454970 110898 455206 111134
rect 485690 111218 485926 111454
rect 485690 110898 485926 111134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76618 579454
rect 76854 579218 87882 579454
rect 88118 579218 99146 579454
rect 99382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76618 579134
rect 76854 578898 87882 579134
rect 88118 578898 99146 579134
rect 99382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 82250 561454
rect 82486 561218 93514 561454
rect 93750 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 82250 561134
rect 82486 560898 93514 561134
rect 93750 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76618 543454
rect 76854 543218 87882 543454
rect 88118 543218 99146 543454
rect 99382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76618 543134
rect 76854 542898 87882 543134
rect 88118 542898 99146 543134
rect 99382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 75618 471454
rect 75854 471218 84882 471454
rect 85118 471218 94146 471454
rect 94382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 75618 471134
rect 75854 470898 84882 471134
rect 85118 470898 94146 471134
rect 94382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 80250 453454
rect 80486 453218 89514 453454
rect 89750 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 80250 453134
rect 80486 452898 89514 453134
rect 89750 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 219610 345454
rect 219846 345218 250330 345454
rect 250566 345218 281050 345454
rect 281286 345218 311770 345454
rect 312006 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 219610 345134
rect 219846 344898 250330 345134
rect 250566 344898 281050 345134
rect 281286 344898 311770 345134
rect 312006 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 204250 327454
rect 204486 327218 234970 327454
rect 235206 327218 265690 327454
rect 265926 327218 296410 327454
rect 296646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 204250 327134
rect 204486 326898 234970 327134
rect 235206 326898 265690 327134
rect 265926 326898 296410 327134
rect 296646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 219610 309454
rect 219846 309218 250330 309454
rect 250566 309218 281050 309454
rect 281286 309218 311770 309454
rect 312006 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 219610 309134
rect 219846 308898 250330 309134
rect 250566 308898 281050 309134
rect 281286 308898 311770 309134
rect 312006 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 204250 291454
rect 204486 291218 234970 291454
rect 235206 291218 265690 291454
rect 265926 291218 296410 291454
rect 296646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 204250 291134
rect 204486 290898 234970 291134
rect 235206 290898 265690 291134
rect 265926 290898 296410 291134
rect 296646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219610 273454
rect 219846 273218 250330 273454
rect 250566 273218 281050 273454
rect 281286 273218 311770 273454
rect 312006 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219610 273134
rect 219846 272898 250330 273134
rect 250566 272898 281050 273134
rect 281286 272898 311770 273134
rect 312006 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204250 255454
rect 204486 255218 234970 255454
rect 235206 255218 265690 255454
rect 265926 255218 296410 255454
rect 296646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204250 255134
rect 204486 254898 234970 255134
rect 235206 254898 265690 255134
rect 265926 254898 296410 255134
rect 296646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 227916 165454
rect 228152 165218 237847 165454
rect 238083 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 314250 165454
rect 314486 165218 317514 165454
rect 317750 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 439610 165454
rect 439846 165218 470330 165454
rect 470566 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 227916 165134
rect 228152 164898 237847 165134
rect 238083 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 314250 165134
rect 314486 164898 317514 165134
rect 317750 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 439610 165134
rect 439846 164898 470330 165134
rect 470566 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 424250 147454
rect 424486 147218 454970 147454
rect 455206 147218 485690 147454
rect 485926 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 424250 147134
rect 424486 146898 454970 147134
rect 455206 146898 485690 147134
rect 485926 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 227916 129454
rect 228152 129218 237847 129454
rect 238083 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 314250 129454
rect 314486 129218 317514 129454
rect 317750 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 439610 129454
rect 439846 129218 470330 129454
rect 470566 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 227916 129134
rect 228152 128898 237847 129134
rect 238083 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 314250 129134
rect 314486 128898 317514 129134
rect 317750 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 439610 129134
rect 439846 128898 470330 129134
rect 470566 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 424250 111454
rect 424486 111218 454970 111454
rect 455206 111218 485690 111454
rect 485926 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 424250 111134
rect 424486 110898 454970 111134
rect 455206 110898 485690 111134
rect 485926 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 70000 0 1 440000
box -10 -52 30000 50000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_hack_soc_dffram  wrapped_hack_soc_dffram_11
timestamp 0
transform 1 0 420000 0 1 100000
box 0 0 74470 79600
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 540000
box -10 -52 36000 42000
use wrapped_teras  wrapped_teras_13
timestamp 0
transform 1 0 200000 0 1 240000
box -10 -52 120000 120000
use wrapped_vga_clock  wrapped_vga_clock_1
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 46000 46000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 388000 74414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 492000 74414 538000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 584000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 388000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 362000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 362000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 362000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 181600 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 181600 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 388000 78134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 492000 78134 538000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 584000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 388000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 362000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 362000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 362000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 181600 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 181600 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 388000 81854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 492000 81854 538000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 584000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 388000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 362000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 362000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 362000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 181600 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 181600 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 388000 85574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 492000 85574 538000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 584000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 362000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 362000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 362000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 181600 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 181600 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 178000 243854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 178000 315854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 388000 99854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 492000 99854 538000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 584000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 362000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 362000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 362000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 362000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 181600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 181600 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 181600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 178000 247574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 178000 319574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 388000 103574 538000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 584000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 362000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 362000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 362000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 362000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 181600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 181600 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 178000 236414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 178000 308414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 388000 92414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 492000 92414 538000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 584000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 362000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 362000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 362000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 362000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 181600 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 181600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 178000 240134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 178000 312134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 388000 96134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 492000 96134 538000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 584000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 362000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 362000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 362000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 362000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 181600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 181600 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 181600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
